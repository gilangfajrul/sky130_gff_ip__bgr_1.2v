magic
tech sky130A
magscale 1 2
timestamp 1716599840
<< checkpaint >>
rect 32307 1615 35419 1668
rect 32307 -1472 35958 1615
rect 32846 -1525 35958 -1472
<< error_p >>
rect 12785 13275 12820 13309
rect 12786 13256 12820 13275
rect 12687 13126 12694 13144
rect 12616 12995 12674 13001
rect 12616 12961 12628 12995
rect 12616 12955 12674 12961
rect 12616 12675 12674 12681
rect 12616 12641 12628 12675
rect 12616 12635 12674 12641
rect 12616 12567 12674 12573
rect 12616 12544 12628 12567
rect 12616 12527 12674 12544
rect 12588 12499 12687 12516
rect 12616 12247 12674 12253
rect 12616 12213 12628 12247
rect 12616 12207 12674 12213
rect 12805 11899 12820 13256
rect 12839 13222 12874 13256
rect 12839 11899 12873 13222
rect 12985 13154 13043 13160
rect 12985 13120 12997 13154
rect 12985 13114 13043 13120
rect 13723 13048 13781 13054
rect 13723 13014 13735 13048
rect 13723 13008 13781 13014
rect 12985 12942 13043 12948
rect 12985 12908 12997 12942
rect 17173 12921 17208 12955
rect 12985 12902 13043 12908
rect 17174 12902 17208 12921
rect 14461 12870 14519 12876
rect 12985 12834 13043 12840
rect 13723 12836 13781 12842
rect 14461 12836 14473 12870
rect 12985 12800 12997 12834
rect 13723 12802 13735 12836
rect 14461 12830 14519 12836
rect 12985 12794 13043 12800
rect 13723 12796 13781 12802
rect 13723 12728 13781 12734
rect 13723 12694 13735 12728
rect 13723 12688 13781 12694
rect 14461 12676 14519 12682
rect 14461 12642 14473 12676
rect 16456 12654 16490 12708
rect 14461 12636 14519 12642
rect 12985 12622 13043 12628
rect 12985 12588 12997 12622
rect 12985 12582 13043 12588
rect 13155 12563 13189 12581
rect 13577 12563 13611 12581
rect 13155 12527 13225 12563
rect 12985 12514 13043 12520
rect 12985 12480 12997 12514
rect 13172 12493 13243 12527
rect 12985 12474 13043 12480
rect 12985 12302 13043 12308
rect 12985 12268 12997 12302
rect 12985 12262 13043 12268
rect 12985 12194 13043 12200
rect 12985 12160 12997 12194
rect 12985 12154 13043 12160
rect 12985 11982 13043 11988
rect 12985 11948 12997 11982
rect 12985 11942 13043 11948
rect 12839 11865 12854 11899
rect 13172 11846 13242 12493
rect 13354 12425 13412 12431
rect 13354 12391 13366 12425
rect 13354 12385 13412 12391
rect 13354 12231 13412 12237
rect 13354 12197 13366 12231
rect 13354 12191 13412 12197
rect 13354 12123 13412 12129
rect 13354 12089 13366 12123
rect 13354 12083 13412 12089
rect 13354 11929 13412 11935
rect 13354 11895 13366 11929
rect 13354 11889 13412 11895
rect 13172 11810 13225 11846
rect 13541 11793 13611 12563
rect 14461 12568 14519 12574
rect 14461 12534 14473 12568
rect 14461 12528 14519 12534
rect 13723 12516 13781 12522
rect 13723 12482 13735 12516
rect 13723 12476 13781 12482
rect 13893 12457 13927 12475
rect 13893 12421 13963 12457
rect 13723 12408 13781 12414
rect 13723 12374 13735 12408
rect 13910 12387 13981 12421
rect 13723 12368 13781 12374
rect 13723 12196 13781 12202
rect 13723 12162 13735 12196
rect 13723 12156 13781 12162
rect 13723 12088 13781 12094
rect 13723 12054 13735 12088
rect 13723 12048 13781 12054
rect 13723 11876 13781 11882
rect 13723 11842 13735 11876
rect 13723 11836 13781 11842
rect 13541 11757 13594 11793
rect 13910 11740 13980 12387
rect 14092 12319 14150 12325
rect 14092 12285 14104 12319
rect 14092 12279 14150 12285
rect 14092 12125 14150 12131
rect 14092 12091 14104 12125
rect 14092 12085 14150 12091
rect 14092 12017 14150 12023
rect 14092 11983 14104 12017
rect 14092 11977 14150 11983
rect 14092 11823 14150 11829
rect 14092 11789 14104 11823
rect 14092 11783 14150 11789
rect 13910 11704 13963 11740
rect 14281 11687 14296 12421
rect 14315 11687 14349 12475
rect 14631 12387 14665 12405
rect 14461 12374 14519 12380
rect 14461 12340 14473 12374
rect 14631 12351 14701 12387
rect 14461 12334 14519 12340
rect 14648 12317 14719 12351
rect 14999 12317 15034 12351
rect 14461 12266 14519 12272
rect 14461 12232 14473 12266
rect 14461 12226 14519 12232
rect 14461 12072 14519 12078
rect 14461 12038 14473 12072
rect 14461 12032 14519 12038
rect 14461 11964 14519 11970
rect 14461 11930 14473 11964
rect 14461 11924 14519 11930
rect 14461 11770 14519 11776
rect 14461 11736 14473 11770
rect 14461 11730 14519 11736
rect 14315 11653 14330 11687
rect 14648 11634 14718 12317
rect 15000 12298 15034 12317
rect 14830 12249 14888 12255
rect 14830 12215 14842 12249
rect 14830 12209 14888 12215
rect 14830 12037 14888 12043
rect 14830 12003 14842 12037
rect 14830 11997 14888 12003
rect 14830 11929 14888 11935
rect 14830 11895 14842 11929
rect 14830 11889 14888 11895
rect 14830 11717 14888 11723
rect 14830 11683 14842 11717
rect 14830 11677 14888 11683
rect 14648 11598 14701 11634
rect 15019 11581 15034 12298
rect 15053 12264 15088 12298
rect 15053 11581 15087 12264
rect 15369 12245 15403 12263
rect 15369 12209 15439 12245
rect 15199 12196 15257 12202
rect 15199 12162 15211 12196
rect 15386 12175 15457 12209
rect 15737 12175 15772 12209
rect 15199 12156 15257 12162
rect 15199 11984 15257 11990
rect 15199 11950 15211 11984
rect 15199 11944 15257 11950
rect 15199 11876 15257 11882
rect 15199 11842 15211 11876
rect 15199 11836 15257 11842
rect 15199 11664 15257 11670
rect 15199 11630 15211 11664
rect 15199 11624 15257 11630
rect 15053 11547 15068 11581
rect 15386 11528 15456 12175
rect 15738 12156 15772 12175
rect 15568 12107 15626 12113
rect 15568 12073 15580 12107
rect 15568 12067 15626 12073
rect 15568 11913 15626 11919
rect 15568 11879 15580 11913
rect 15568 11873 15626 11879
rect 15568 11805 15626 11811
rect 15568 11771 15580 11805
rect 15568 11765 15626 11771
rect 15568 11611 15626 11617
rect 15568 11577 15580 11611
rect 15568 11571 15626 11577
rect 15386 11492 15439 11528
rect 15757 11475 15772 12156
rect 15791 12122 15826 12156
rect 15791 11475 15825 12122
rect 15937 12054 15995 12060
rect 15937 12020 15949 12054
rect 15937 12014 15995 12020
rect 15937 11860 15995 11866
rect 15937 11826 15949 11860
rect 15937 11820 15995 11826
rect 15937 11752 15995 11758
rect 15937 11718 15949 11752
rect 15937 11712 15995 11718
rect 15937 11558 15995 11564
rect 15937 11524 15949 11558
rect 15937 11518 15995 11524
rect 15791 11441 15806 11475
rect 16126 11422 16141 12156
rect 16160 11422 16194 12210
rect 16160 11388 16175 11422
rect 16475 11369 16490 12654
rect 16509 12620 16544 12654
rect 16509 11369 16543 12620
rect 16655 12552 16713 12558
rect 16655 12518 16667 12552
rect 16655 12512 16713 12518
rect 16655 12358 16713 12364
rect 16655 12324 16667 12358
rect 16655 12318 16713 12324
rect 16655 12250 16713 12256
rect 16655 12216 16667 12250
rect 16655 12210 16713 12216
rect 16655 12056 16713 12062
rect 16655 12022 16667 12056
rect 16655 12016 16713 12022
rect 16655 11948 16713 11954
rect 16655 11914 16667 11948
rect 16655 11908 16713 11914
rect 16655 11754 16713 11760
rect 16655 11720 16667 11754
rect 16655 11714 16713 11720
rect 16655 11646 16713 11652
rect 16655 11612 16667 11646
rect 16655 11606 16713 11612
rect 16655 11452 16713 11458
rect 16655 11418 16667 11452
rect 16655 11412 16713 11418
rect 16509 11335 16524 11369
rect 16844 11316 16859 12654
rect 16878 11316 16912 12708
rect 16878 11282 16893 11316
rect 17193 11263 17208 12902
rect 17227 12868 17262 12902
rect 17227 11263 17261 12868
rect 17227 11229 17242 11263
rect 28493 968 28528 1002
rect 28494 949 28528 968
rect 28513 436 28528 949
rect 28547 915 28582 949
rect 30832 915 30867 949
rect 28547 436 28581 915
rect 30833 896 30867 915
rect 28547 402 28562 436
rect 30852 383 30867 896
rect 30886 862 30921 896
rect 30886 383 30920 862
rect 30886 349 30901 383
<< error_s >>
rect 25777 1917 25823 1934
rect 25749 1889 25851 1906
rect 25749 1706 25851 1727
rect 25777 1678 25823 1699
rect 1366 26 1368 1314
rect 11643 153 11797 1429
rect 11994 1359 12029 1393
rect 11995 1340 12029 1359
rect 11825 1291 11883 1297
rect 11825 1257 11837 1291
rect 11825 1251 11883 1257
rect 11825 1079 11883 1085
rect 11825 1045 11837 1079
rect 11825 1039 11883 1045
rect 11825 971 11883 977
rect 11825 937 11837 971
rect 11825 931 11883 937
rect 11825 759 11883 765
rect 11825 725 11837 759
rect 11825 719 11883 725
rect 11825 651 11883 657
rect 11825 617 11837 651
rect 11825 611 11883 617
rect 11825 439 11883 445
rect 11825 405 11837 439
rect 11825 399 11883 405
rect 11825 331 11883 337
rect 11825 297 11837 331
rect 11825 291 11883 297
rect 11643 26 11713 153
rect 11825 119 11883 125
rect 11825 85 11837 119
rect 11825 79 11883 85
rect 11643 0 11704 26
rect 11679 -8 11704 0
rect 12014 -17 12029 1340
rect 12048 1306 12083 1340
rect 25749 1306 25851 1309
rect 12048 -17 12082 1306
rect 25777 1278 25823 1281
rect 12194 1238 12252 1244
rect 12194 1204 12206 1238
rect 12194 1198 12252 1204
rect 26155 1038 26189 1056
rect 12194 1026 12252 1032
rect 12194 992 12206 1026
rect 26155 1002 26225 1038
rect 12194 986 12252 992
rect 26172 968 26243 1002
rect 12194 918 12252 924
rect 12194 884 12206 918
rect 12194 878 12252 884
rect 12194 706 12252 712
rect 12194 672 12206 706
rect 12194 666 12252 672
rect 12194 598 12252 604
rect 12194 564 12206 598
rect 12194 558 12252 564
rect 26172 489 26242 968
rect 24455 434 24490 468
rect 26172 453 26225 489
rect 33225 932 33259 950
rect 24456 415 24490 434
rect 12194 386 12252 392
rect 12194 352 12206 386
rect 24286 366 24344 372
rect 12194 346 12252 352
rect 24286 332 24298 366
rect 24286 326 24344 332
rect 12194 278 12252 284
rect 12194 244 12206 278
rect 12194 238 12252 244
rect 24286 172 24344 178
rect 24286 138 24298 172
rect 24286 132 24344 138
rect 12194 66 12252 72
rect 12194 32 12206 66
rect 24475 36 24490 415
rect 24509 381 24544 415
rect 24824 381 24859 415
rect 24509 36 24543 381
rect 24825 362 24859 381
rect 24655 313 24713 319
rect 24655 279 24667 313
rect 24655 273 24713 279
rect 24655 119 24713 125
rect 24655 85 24667 119
rect 24655 79 24713 85
rect 12194 26 12252 32
rect 24509 2 24524 36
rect 24844 -17 24859 362
rect 24878 328 24913 362
rect 25193 328 25228 362
rect 24878 -17 24912 328
rect 25194 309 25228 328
rect 33189 330 33259 932
rect 33549 372 33555 426
rect 25024 260 25082 266
rect 25024 226 25036 260
rect 25024 220 25082 226
rect 25024 66 25082 72
rect 25024 32 25036 66
rect 25024 26 25082 32
rect 12048 -51 12063 -17
rect 24878 -51 24893 -17
rect 25213 -70 25228 309
rect 25247 275 25282 309
rect 33189 294 33242 330
rect 25247 -70 25281 275
rect 25393 207 25451 213
rect 25393 173 25405 207
rect 25393 167 25451 173
rect 25393 13 25451 19
rect 25393 -21 25405 13
rect 25393 -27 25451 -21
rect 25247 -104 25262 -70
rect 33603 -123 33609 372
use op5  x1
timestamp 1716599838
transform 1 0 12487 0 1 13516
box -53 -13622 8878 1258
use Resistor492k_1  x2
timestamp 1716599839
transform 1 0 23704 0 1 1441
box 0 -1600 200 200
use Resistor492k_1  x3
timestamp 1716599839
transform 1 0 23904 0 1 1441
box 0 -1600 200 200
use Resistor50k_1  x4
timestamp 1716599839
transform 1 0 24151 0 1 453
box -47 -612 1482 200
use Startup  x5
timestamp 1716599840
transform 1 0 25686 0 1 2106
box -53 -2265 7934 2299
use sky130_fd_pr__pfet_01v8_M47T9Z  XM1
timestamp 0
transform 1 0 11854 0 1 688
box -211 -741 211 741
use sky130_fd_pr__pfet_01v8_M47T9Z  XM2
timestamp 0
transform 1 0 12223 0 1 635
box -211 -741 211 741
use sky130_fd_pr__nfet_01v8_lvt_69TQ3K  XM3
timestamp 0
transform 1 0 33863 0 1 98
box -296 -310 296 310
use sky130_fd_pr__nfet_01v8_lvt_69TQ3K  XM4
timestamp 0
transform 1 0 34402 0 1 45
box -296 -310 296 310
use sky130_fd_pr__pfet_01v8_6H4VWJ  XM15
timestamp 0
transform 1 0 22508 0 1 814
box -1196 -973 1196 973
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  XQ1 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1716538025
transform 1 0 0 0 1 0
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  XQ2
array 0 7 1288 0 0 1288
timestamp 1716538025
transform 1 0 1340 0 1 0
box 0 0 1340 1340
<< end >>
