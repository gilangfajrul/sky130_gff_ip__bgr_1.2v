magic
tech sky130A
magscale 1 2
timestamp 1716365683
<< metal3 >>
rect -3892 3172 -120 3200
rect -3892 148 -204 3172
rect -140 148 -120 3172
rect -3892 120 -120 148
rect 120 3172 3892 3200
rect 120 148 3808 3172
rect 3872 148 3892 3172
rect 120 120 3892 148
rect -3892 -148 -120 -120
rect -3892 -3172 -204 -148
rect -140 -3172 -120 -148
rect -3892 -3200 -120 -3172
rect 120 -148 3892 -120
rect 120 -3172 3808 -148
rect 3872 -3172 3892 -148
rect 120 -3200 3892 -3172
<< via3 >>
rect -204 148 -140 3172
rect 3808 148 3872 3172
rect -204 -3172 -140 -148
rect 3808 -3172 3872 -148
<< mimcap >>
rect -3852 3120 -452 3160
rect -3852 200 -3812 3120
rect -492 200 -452 3120
rect -3852 160 -452 200
rect 160 3120 3560 3160
rect 160 200 200 3120
rect 3520 200 3560 3120
rect 160 160 3560 200
rect -3852 -200 -452 -160
rect -3852 -3120 -3812 -200
rect -492 -3120 -452 -200
rect -3852 -3160 -452 -3120
rect 160 -200 3560 -160
rect 160 -3120 200 -200
rect 3520 -3120 3560 -200
rect 160 -3160 3560 -3120
<< mimcapcontact >>
rect -3812 200 -492 3120
rect 200 200 3520 3120
rect -3812 -3120 -492 -200
rect 200 -3120 3520 -200
<< metal4 >>
rect -2204 3121 -2100 3320
rect -224 3172 -120 3320
rect -3813 3120 -491 3121
rect -3813 200 -3812 3120
rect -492 200 -491 3120
rect -3813 199 -491 200
rect -2204 -199 -2100 199
rect -224 148 -204 3172
rect -140 148 -120 3172
rect 1808 3121 1912 3320
rect 3788 3172 3892 3320
rect 199 3120 3521 3121
rect 199 200 200 3120
rect 3520 200 3521 3120
rect 199 199 3521 200
rect -224 -148 -120 148
rect -3813 -200 -491 -199
rect -3813 -3120 -3812 -200
rect -492 -3120 -491 -200
rect -3813 -3121 -491 -3120
rect -2204 -3320 -2100 -3121
rect -224 -3172 -204 -148
rect -140 -3172 -120 -148
rect 1808 -199 1912 199
rect 3788 148 3808 3172
rect 3872 148 3892 3172
rect 3788 -148 3892 148
rect 199 -200 3521 -199
rect 199 -3120 200 -200
rect 3520 -3120 3521 -200
rect 199 -3121 3521 -3120
rect -224 -3320 -120 -3172
rect 1808 -3320 1912 -3121
rect 3788 -3172 3808 -148
rect 3872 -3172 3892 -148
rect 3788 -3320 3892 -3172
<< properties >>
string FIXED_BBOX 120 120 3600 3200
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 17 l 15 val 522.159 carea 2.00 cperi 0.19 nx 2 ny 2 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
