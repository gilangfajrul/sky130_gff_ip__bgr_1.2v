magic
tech sky130A
magscale 1 2
timestamp 1717432527
<< error_p >>
rect -29 -87 29 -81
rect -29 -121 -17 -87
rect -29 -127 29 -121
<< nmos >>
rect -15 -49 15 111
<< ndiff >>
rect -73 99 -15 111
rect -73 -37 -61 99
rect -27 -37 -15 99
rect -73 -49 -15 -37
rect 15 99 73 111
rect 15 -37 27 99
rect 61 -37 73 99
rect 15 -49 73 -37
<< ndiffc >>
rect -61 -37 -27 99
rect 27 -37 61 99
<< poly >>
rect -15 111 15 137
rect -15 -71 15 -49
rect -33 -87 33 -71
rect -33 -121 -17 -87
rect 17 -121 33 -87
rect -33 -137 33 -121
<< polycont >>
rect -17 -121 17 -87
<< locali >>
rect -61 99 -27 115
rect -61 -53 -27 -37
rect 27 99 61 115
rect 27 -53 61 -37
rect -33 -121 -17 -87
rect 17 -121 33 -87
<< viali >>
rect -61 -37 -27 99
rect 27 -37 61 99
rect -17 -121 17 -87
<< metal1 >>
rect -67 99 -21 111
rect -67 -37 -61 99
rect -27 -37 -21 99
rect -67 -49 -21 -37
rect 21 99 67 111
rect 21 -37 27 99
rect 61 -37 67 99
rect 21 -49 67 -37
rect -29 -87 29 -81
rect -29 -121 -17 -87
rect 17 -121 29 -87
rect -29 -127 29 -121
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.8 l 0.150 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
