magic
tech sky130A
magscale 1 2
timestamp 1762860936
<< dnwell >>
rect -1012 -8432 27624 10622
<< nwell >>
rect -1092 10416 27704 10702
rect -1092 -8226 -806 10416
rect 27418 -8226 27704 10416
rect -1092 -8512 27704 -8226
<< pwell >>
rect 352 -3415 494 -3301
<< nsubdiff >>
rect -1055 10645 27667 10665
rect -1055 10611 -975 10645
rect 27587 10611 27667 10645
rect -1055 10591 27667 10611
rect -1055 10585 -981 10591
rect -1055 -8395 -1035 10585
rect -1001 -8395 -981 10585
rect -1055 -8401 -981 -8395
rect 27593 10585 27667 10591
rect 27593 -8395 27613 10585
rect 27647 -8395 27667 10585
rect 27593 -8401 27667 -8395
rect -1055 -8421 27667 -8401
rect -1055 -8455 -975 -8421
rect 27587 -8455 27667 -8421
rect -1055 -8475 27667 -8455
<< nsubdiffcont >>
rect -975 10611 27587 10645
rect -1035 -8395 -1001 10585
rect 27613 -8395 27647 10585
rect -975 -8455 27587 -8421
<< locali >>
rect -1035 10611 -975 10645
rect 27587 10611 27647 10645
rect -1035 10585 -1001 10611
rect -1035 -8421 -1001 -8395
rect 27613 10585 27647 10611
rect 27613 -8421 27647 -8395
rect -1035 -8455 -975 -8421
rect 27587 -8455 27647 -8421
<< metal1 >>
rect 17231 5947 17283 5953
rect 17283 5895 19463 5947
rect 19515 5895 19521 5947
rect 17231 5889 17283 5895
rect 19160 2845 19240 2851
rect 16812 2790 16822 2842
rect 18106 2790 18116 2842
rect 19240 2765 19450 2845
rect 19530 2765 19536 2845
rect 19160 2759 19240 2765
rect 18870 -851 18876 -727
rect 19000 -851 29502 -727
rect 29626 -851 29632 -727
rect -4547 -1266 -4537 -1090
rect -4485 -1266 -4475 -1090
rect -3433 -1267 -3423 -1090
rect -3371 -1267 -3361 -1090
rect 9397 -1310 9407 -1238
rect 9479 -1310 19295 -1238
rect 19367 -1310 19377 -1238
rect -3423 -1396 -3371 -1390
rect -494 -1396 -442 -1390
rect -3371 -1448 -494 -1396
rect -3423 -1454 -3371 -1448
rect -494 -1454 -442 -1448
rect -1001 -1494 -949 -1488
rect -4543 -1546 -4537 -1494
rect -4485 -1546 -1001 -1494
rect -1001 -1552 -949 -1546
rect -2786 -1977 -2780 -1925
rect -2728 -1926 -2722 -1925
rect -144 -1926 -138 -1925
rect -2728 -1976 -138 -1926
rect -2728 -1977 -2722 -1976
rect -144 -1977 -138 -1976
rect -86 -1977 -80 -1925
rect 4529 -2291 4581 -2285
rect 4581 -2343 26555 -2291
rect 26607 -2343 26613 -2291
rect 4529 -2349 4581 -2343
rect 26778 -2544 26830 -2538
rect 8635 -2596 8645 -2544
rect 8697 -2596 26778 -2544
rect 26830 -2596 26840 -2544
rect 26778 -2602 26830 -2596
rect 9406 -2719 9416 -2663
rect 9472 -2719 9482 -2663
rect -2790 -2869 -2784 -2817
rect -2732 -2818 -2726 -2817
rect -311 -2818 -305 -2817
rect -2732 -2868 -305 -2818
rect -2732 -2869 -2726 -2868
rect -311 -2869 -305 -2868
rect -253 -2869 -247 -2817
rect 13219 -2821 29848 -2731
rect 29982 -2821 29992 -2731
rect 13219 -3026 13269 -2821
rect 32174 -2987 32184 -2447
rect 32724 -2987 32734 -2447
rect -138 -3084 -86 -3078
rect -86 -3135 272 -3085
rect -138 -3142 -86 -3136
rect -688 -3392 -682 -3326
rect -616 -3392 352 -3326
rect -50 -3709 2 -3703
rect -2794 -3761 -2788 -3709
rect -2736 -3761 -50 -3709
rect -50 -3767 2 -3761
rect -305 -3988 -253 -3982
rect -253 -4039 189 -3989
rect -305 -4046 -253 -4040
rect -2776 -4662 -2770 -4596
rect -2704 -4662 -136 -4596
rect -70 -4662 -64 -4596
rect -500 -4782 -494 -4730
rect -442 -4782 8463 -4730
rect 8515 -4782 8521 -4730
rect 19296 -4813 19368 -4807
rect -3855 -4910 -3845 -4858
rect -3069 -4910 -3059 -4858
rect -2774 -4916 -2768 -4850
rect -2702 -4916 -682 -4850
rect -616 -4916 -610 -4850
rect 8985 -4885 8991 -4813
rect 9063 -4885 19296 -4813
rect 19296 -4891 19368 -4885
rect 26329 -4939 26339 -4938
rect 18892 -5012 18902 -4940
rect 18974 -5012 26339 -4939
rect 26411 -5010 26421 -4938
rect -1007 -5134 -1001 -5082
rect -949 -5134 4126 -5082
rect 4178 -5134 4184 -5082
rect 17287 -5184 17297 -5108
rect 17373 -5184 25868 -5108
rect 25944 -5184 25954 -5108
rect 25626 -5645 25636 -5593
rect 26033 -5645 26043 -5593
rect 25626 -5811 25636 -5759
rect 26033 -5811 26043 -5759
rect 8819 -6309 8829 -6257
rect 9226 -6309 9236 -6257
rect 8282 -6475 8292 -6423
rect 8689 -6475 8699 -6423
rect 25626 -6641 25636 -6589
rect 26033 -6641 26043 -6589
rect 25626 -6807 25636 -6755
rect 26033 -6807 26043 -6755
<< via1 >>
rect 17231 5895 17283 5947
rect 19463 5895 19515 5947
rect 16822 2790 18106 2842
rect 19160 2765 19240 2845
rect 19450 2765 19530 2845
rect 18876 -851 19000 -727
rect 29502 -851 29626 -727
rect -4537 -1266 -4485 -1090
rect -3423 -1267 -3371 -1090
rect 9407 -1310 9479 -1238
rect 19295 -1310 19367 -1238
rect -3423 -1448 -3371 -1396
rect -494 -1448 -442 -1396
rect -4537 -1546 -4485 -1494
rect -1001 -1546 -949 -1494
rect -2780 -1977 -2728 -1925
rect -138 -1977 -86 -1925
rect 4529 -2343 4581 -2291
rect 26555 -2343 26607 -2291
rect 8645 -2596 8697 -2544
rect 26778 -2596 26830 -2544
rect 9416 -2719 9472 -2663
rect -2784 -2869 -2732 -2817
rect -305 -2869 -253 -2817
rect 29848 -2821 29982 -2731
rect 32184 -2987 32724 -2447
rect -138 -3136 -86 -3084
rect -682 -3392 -616 -3326
rect -2788 -3761 -2736 -3709
rect -50 -3761 2 -3709
rect -305 -4040 -253 -3988
rect -2770 -4662 -2704 -4596
rect -136 -4662 -70 -4596
rect -494 -4782 -442 -4730
rect 8463 -4782 8515 -4730
rect -3845 -4910 -3069 -4858
rect -2768 -4916 -2702 -4850
rect -682 -4916 -616 -4850
rect 8991 -4885 9063 -4813
rect 19296 -4885 19368 -4813
rect 18902 -5012 18974 -4940
rect 26339 -5010 26411 -4938
rect -1001 -5134 -949 -5082
rect 4126 -5134 4178 -5082
rect 17297 -5184 17373 -5108
rect 25868 -5184 25944 -5108
rect 25636 -5645 26033 -5593
rect 25636 -5811 26033 -5759
rect 8829 -6309 9226 -6257
rect 8292 -6475 8689 -6423
rect 25636 -6641 26033 -6589
rect 25636 -6807 26033 -6755
<< metal2 >>
rect 17231 5947 17283 7177
rect 19463 5947 19515 5953
rect 17225 5895 17231 5947
rect 17283 5895 17289 5947
rect 18084 2928 19374 2986
rect 16822 2845 18106 2852
rect 16822 2842 19160 2845
rect 18106 2790 19160 2842
rect 16822 2787 19160 2790
rect 16822 2780 18106 2787
rect 18898 2765 19160 2787
rect 19240 2765 19246 2845
rect 9034 1546 9095 1549
rect 9027 1490 9036 1546
rect 9092 1490 9101 1546
rect -4537 -1090 -4485 -1079
rect -4537 -1494 -4485 -1266
rect -3423 -1090 -3371 -1078
rect 9034 -1267 9095 1490
rect 18898 -721 18978 2765
rect 18876 -727 19000 -721
rect 18876 -857 19000 -851
rect -3423 -1396 -3371 -1267
rect 8754 -1328 9095 -1267
rect 9407 -1238 9479 -1228
rect -3429 -1448 -3423 -1396
rect -3371 -1448 -3365 -1396
rect -500 -1448 -494 -1396
rect -442 -1448 -436 -1396
rect -1007 -1546 -1001 -1494
rect -949 -1546 -943 -1494
rect -4537 -1552 -4485 -1546
rect -2780 -1925 -2728 -1919
rect -3845 -1976 -2780 -1926
rect -2780 -1983 -2728 -1977
rect -2784 -2817 -2732 -2811
rect -3846 -2868 -2784 -2818
rect -2784 -2875 -2732 -2869
rect -2788 -3709 -2736 -3703
rect -3844 -3761 -2788 -3709
rect -2788 -3767 -2736 -3761
rect -2770 -4596 -2704 -4590
rect -3845 -4662 -2770 -4596
rect -2770 -4668 -2704 -4662
rect -3845 -4850 -3069 -4848
rect -2768 -4850 -2702 -4844
rect -3845 -4858 -2768 -4850
rect -3069 -4910 -2768 -4858
rect -3845 -4916 -2768 -4910
rect -3845 -4920 -3069 -4916
rect -2768 -4922 -2702 -4916
rect -1001 -5082 -949 -1546
rect -682 -3326 -616 -3320
rect -682 -4850 -616 -3392
rect -494 -4730 -442 -1448
rect -138 -1925 -86 -1919
rect -138 -1983 -86 -1977
rect -305 -2817 -253 -2811
rect -305 -2875 -253 -2869
rect -304 -3988 -254 -2875
rect -137 -3084 -87 -1983
rect 4529 -2291 4581 -1340
rect 4523 -2343 4529 -2291
rect 4581 -2343 4587 -2291
rect 8645 -2544 8697 -1413
rect 8645 -2606 8697 -2596
rect 9407 -2663 9479 -1310
rect 9415 -2719 9416 -2663
rect 9472 -2719 9473 -2663
rect 9415 -2720 9473 -2719
rect 9416 -2729 9472 -2720
rect -144 -3136 -138 -3084
rect -86 -3136 -80 -3084
rect -56 -3761 -50 -3709
rect 2 -3761 190 -3709
rect -311 -4040 -305 -3988
rect -253 -4040 -247 -3988
rect -131 -4239 -75 -4235
rect -136 -4244 -70 -4239
rect -136 -4300 -131 -4244
rect -75 -4300 -70 -4244
rect -136 -4596 -70 -4300
rect -136 -4668 -70 -4662
rect -494 -4788 -442 -4782
rect 8463 -4730 8515 -4724
rect -682 -4922 -616 -4916
rect -1001 -5140 -949 -5134
rect 4126 -5082 4178 -5076
rect 4126 -6423 4178 -5134
rect 8463 -6413 8515 -4782
rect 8991 -4813 9063 -4807
rect 8991 -6247 9063 -4885
rect 18898 -4940 18978 -857
rect 19290 -1238 19374 2928
rect 19463 2851 19515 5895
rect 19450 2845 19530 2851
rect 19450 2759 19530 2765
rect 19290 -1310 19295 -1238
rect 19367 -1310 19374 -1238
rect 19290 -4813 19374 -1310
rect 29502 -727 29626 -721
rect 29502 -1274 29626 -851
rect 29502 -1398 30085 -1274
rect 19290 -4885 19296 -4813
rect 19368 -4885 19374 -4813
rect 26555 -2291 26607 -2285
rect 18898 -5012 18902 -4940
rect 18974 -5012 18978 -4940
rect 18898 -5022 18978 -5012
rect 26339 -4938 26411 -4928
rect 17297 -5108 17373 -5098
rect 25868 -5108 25944 -5098
rect 17293 -5179 17297 -5113
rect 17373 -5179 17377 -5113
rect 17297 -5194 17373 -5184
rect 25868 -5194 25944 -5184
rect 25636 -5591 26033 -5581
rect 25636 -5657 26033 -5647
rect 26339 -5749 26411 -5010
rect 25636 -5759 26411 -5749
rect 26033 -5811 26411 -5759
rect 25636 -5821 26411 -5811
rect 17307 -6099 17363 -6089
rect 17307 -6165 17363 -6155
rect 8829 -6257 9226 -6247
rect 8829 -6319 9226 -6309
rect 8292 -6423 8689 -6413
rect 4126 -6475 4415 -6423
rect 8292 -6485 8689 -6475
rect 25636 -6589 26033 -6579
rect 26555 -6589 26607 -2343
rect 32184 -2447 32724 -2437
rect 26778 -2544 26830 -2534
rect 26772 -2596 26778 -2544
rect 26830 -2596 26836 -2544
rect 26033 -6641 26607 -6589
rect 25636 -6651 26033 -6641
rect 25636 -6755 26033 -6745
rect 26778 -6755 26830 -2596
rect 29848 -2731 29982 -2721
rect 29982 -2821 32184 -2731
rect 29848 -2831 29982 -2821
rect 32184 -2997 32724 -2987
rect 25634 -6807 25636 -6755
rect 26033 -6807 26830 -6755
rect 25636 -6817 26033 -6807
<< via2 >>
rect 9036 1490 9092 1546
rect 9416 -2719 9472 -2663
rect -131 -4300 -75 -4244
rect 17302 -5179 17368 -5113
rect 25868 -5184 25944 -5118
rect 25636 -5593 26033 -5591
rect 25636 -5645 26033 -5593
rect 25636 -5647 26033 -5645
rect 17307 -6155 17363 -6099
<< metal3 >>
rect 9031 1546 9097 1551
rect 9031 1490 9036 1546
rect 9092 1490 9097 1546
rect 9031 1485 9097 1490
rect 9396 -2659 9496 -2641
rect 9396 -2723 9412 -2659
rect 9476 -2723 9496 -2659
rect 9396 -2741 9496 -2723
rect -136 -4244 2600 -4239
rect -136 -4300 -131 -4244
rect -75 -4300 2600 -4244
rect -136 -4305 2600 -4300
rect 17297 -5113 17373 -5108
rect 17297 -5179 17302 -5113
rect 17368 -5179 17373 -5113
rect 17297 -6099 17373 -5179
rect 25858 -5118 25954 -5113
rect 25858 -5184 25868 -5118
rect 25944 -5184 25954 -5118
rect 25858 -5189 25954 -5184
rect 25868 -5586 25944 -5189
rect 25626 -5591 26043 -5586
rect 25626 -5647 25636 -5591
rect 26033 -5647 26043 -5591
rect 25626 -5652 26043 -5647
rect 17297 -6155 17307 -6099
rect 17363 -6155 17373 -6099
rect 17297 -6160 17373 -6155
<< via3 >>
rect 9412 -2663 9476 -2659
rect 9412 -2719 9416 -2663
rect 9416 -2719 9472 -2663
rect 9472 -2719 9476 -2663
rect 9412 -2723 9476 -2719
<< metal4 >>
rect 9411 -2659 9477 -2658
rect 9411 -2723 9412 -2659
rect 9476 -2723 9477 -2659
rect 9411 -2973 9477 -2723
use bjt  bjt_0
timestamp 1762855819
transform -1 0 37289 0 -1 2118
box -387 -387 7328 7279
use digital  digital_0
timestamp 1720189102
transform 1 0 -4922 0 1 -4244
box -397 -1200 2333 5008
use op5  op5_0
timestamp 1762786734
transform 1 0 9786 0 1 -6121
box -9786 6121 9272 13721
use pmos_current_bgr  pmos_current_bgr_0
timestamp 1762753955
transform 1 0 425 0 1 -1186
box -227 -676 8487 506
use res_trim  res_trim_0
timestamp 1720030020
transform 0 1 101 -1 0 -2857
box -31 -51 1533 15873
use resist_const  resist_const_0
timestamp 1720269525
transform -1 0 28465 0 -1 -9225
box 2257 -3964 28483 -2103
use startupcir  startupcir_0
timestamp 1762846550
transform -1 0 21906 0 -1 7909
box -20 -1581 21888 938
<< end >>
