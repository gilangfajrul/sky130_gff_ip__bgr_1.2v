magic
tech sky130A
magscale 1 2
timestamp 1716365683
<< metal3 >>
rect -386 3172 386 3200
rect -386 148 302 3172
rect 366 148 386 3172
rect -386 120 386 148
rect -386 -148 386 -120
rect -386 -3172 302 -148
rect 366 -3172 386 -148
rect -386 -3200 386 -3172
<< via3 >>
rect 302 148 366 3172
rect 302 -3172 366 -148
<< mimcap >>
rect -346 3120 54 3160
rect -346 200 -306 3120
rect 14 200 54 3120
rect -346 160 54 200
rect -346 -200 54 -160
rect -346 -3120 -306 -200
rect 14 -3120 54 -200
rect -346 -3160 54 -3120
<< mimcapcontact >>
rect -306 200 14 3120
rect -306 -3120 14 -200
<< metal4 >>
rect -198 3121 -94 3320
rect 282 3172 386 3320
rect -307 3120 15 3121
rect -307 200 -306 3120
rect 14 200 15 3120
rect -307 199 15 200
rect -198 -199 -94 199
rect 282 148 302 3172
rect 366 148 386 3172
rect 282 -148 386 148
rect -307 -200 15 -199
rect -307 -3120 -306 -200
rect 14 -3120 15 -200
rect -307 -3121 15 -3120
rect -198 -3320 -94 -3121
rect 282 -3172 302 -148
rect 366 -3172 386 -148
rect 282 -3320 386 -3172
<< properties >>
string FIXED_BBOX -386 120 94 3200
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 2.00 l 15 val 66.46 carea 2.00 cperi 0.19 nx 1 ny 2 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
