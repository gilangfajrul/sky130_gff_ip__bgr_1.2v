magic
tech sky130A
magscale 1 2
timestamp 1717771017
<< nwell >>
rect -523 -164 523 198
<< pmos >>
rect -429 -64 -29 136
rect 29 -64 429 136
<< pdiff >>
rect -487 124 -429 136
rect -487 -52 -475 124
rect -441 -52 -429 124
rect -487 -64 -429 -52
rect -29 124 29 136
rect -29 -52 -17 124
rect 17 -52 29 124
rect -29 -64 29 -52
rect 429 124 487 136
rect 429 -52 441 124
rect 475 -52 487 124
rect 429 -64 487 -52
<< pdiffc >>
rect -475 -52 -441 124
rect -17 -52 17 124
rect 441 -52 475 124
<< poly >>
rect -429 136 -29 162
rect 29 136 429 162
rect -429 -111 -29 -64
rect -429 -128 -321 -111
rect -337 -145 -321 -128
rect -137 -128 -29 -111
rect 29 -111 429 -64
rect 29 -128 137 -111
rect -137 -145 -121 -128
rect -337 -161 -121 -145
rect 121 -145 137 -128
rect 321 -128 429 -111
rect 321 -145 337 -128
rect 121 -161 337 -145
<< polycont >>
rect -321 -145 -137 -111
rect 137 -145 321 -111
<< locali >>
rect -475 124 -441 140
rect -475 -68 -441 -52
rect -17 124 17 140
rect -17 -68 17 -52
rect 441 124 475 140
rect 441 -68 475 -52
rect -337 -145 -321 -111
rect -137 -145 -121 -111
rect 121 -145 137 -111
rect 321 -145 337 -111
<< viali >>
rect -475 -52 -441 124
rect -17 -52 17 124
rect 441 -52 475 124
rect -321 -145 -137 -111
rect 137 -145 321 -111
<< metal1 >>
rect -481 124 -435 136
rect -481 -52 -475 124
rect -441 -52 -435 124
rect -481 -64 -435 -52
rect -23 124 23 136
rect -23 -52 -17 124
rect 17 -52 23 124
rect -23 -64 23 -52
rect 435 124 481 136
rect 435 -52 441 124
rect 475 -52 481 124
rect 435 -64 481 -52
rect -333 -111 -125 -105
rect -333 -145 -321 -111
rect -137 -145 -125 -111
rect -333 -151 -125 -145
rect 125 -111 333 -105
rect 125 -145 137 -111
rect 321 -145 333 -111
rect 125 -151 333 -145
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 2 m 1 nf 2 diffcov 100 polycov 50 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
