magic
tech sky130A
magscale 1 2
timestamp 1716599838
<< checkpaint >>
rect 3846 841 10138 2518
rect 2377 752 10138 841
rect 532 -3178 10138 752
rect 2377 -3443 10138 -3178
rect 2726 -3496 10138 -3443
rect 3095 -3549 10138 -3496
rect 3444 -3602 10138 -3549
rect 3846 -14882 10138 -3602
<< error_s >>
rect 298 -241 333 -207
rect 299 -260 333 -241
rect 200 -390 207 -372
rect 129 -521 187 -515
rect 129 -555 141 -521
rect 129 -561 187 -555
rect 129 -841 187 -835
rect 129 -875 141 -841
rect 129 -881 187 -875
rect 129 -949 187 -943
rect 129 -972 141 -949
rect 129 -989 187 -972
rect 101 -1017 200 -1000
rect 129 -1269 187 -1263
rect 129 -1303 141 -1269
rect 129 -1309 187 -1303
rect 318 -1617 333 -260
rect 352 -294 387 -260
rect 352 -1617 386 -294
rect 498 -362 556 -356
rect 498 -396 510 -362
rect 498 -402 556 -396
rect 1236 -468 1294 -462
rect 1236 -502 1248 -468
rect 1236 -508 1294 -502
rect 498 -574 556 -568
rect 498 -608 510 -574
rect 498 -614 556 -608
rect 1974 -646 2032 -640
rect 498 -682 556 -676
rect 1236 -680 1294 -674
rect 1974 -680 1986 -646
rect 498 -716 510 -682
rect 1236 -714 1248 -680
rect 1974 -686 2032 -680
rect 498 -722 556 -716
rect 1236 -720 1294 -714
rect 1236 -788 1294 -782
rect 1236 -822 1248 -788
rect 1236 -828 1294 -822
rect 1974 -840 2032 -834
rect 1974 -874 1986 -840
rect 1974 -880 2032 -874
rect 498 -894 556 -888
rect 498 -928 510 -894
rect 498 -934 556 -928
rect 668 -953 702 -935
rect 1090 -953 1124 -935
rect 668 -989 738 -953
rect 498 -1002 556 -996
rect 498 -1036 510 -1002
rect 685 -1023 756 -989
rect 498 -1042 556 -1036
rect 498 -1214 556 -1208
rect 498 -1248 510 -1214
rect 498 -1254 556 -1248
rect 498 -1322 556 -1316
rect 498 -1356 510 -1322
rect 498 -1362 556 -1356
rect 498 -1534 556 -1528
rect 498 -1568 510 -1534
rect 498 -1574 556 -1568
rect 352 -1651 367 -1617
rect 685 -1670 755 -1023
rect 867 -1091 925 -1085
rect 867 -1125 879 -1091
rect 867 -1131 925 -1125
rect 867 -1285 925 -1279
rect 867 -1319 879 -1285
rect 867 -1325 925 -1319
rect 867 -1393 925 -1387
rect 867 -1427 879 -1393
rect 867 -1433 925 -1427
rect 867 -1587 925 -1581
rect 867 -1621 879 -1587
rect 867 -1627 925 -1621
rect 685 -1706 738 -1670
rect 1054 -1723 1124 -953
rect 1974 -948 2032 -942
rect 1974 -982 1986 -948
rect 1974 -988 2032 -982
rect 1236 -1000 1294 -994
rect 1236 -1034 1248 -1000
rect 1236 -1040 1294 -1034
rect 1406 -1059 1440 -1041
rect 1406 -1095 1476 -1059
rect 1236 -1108 1294 -1102
rect 1236 -1142 1248 -1108
rect 1423 -1129 1494 -1095
rect 1236 -1148 1294 -1142
rect 1236 -1320 1294 -1314
rect 1236 -1354 1248 -1320
rect 1236 -1360 1294 -1354
rect 1236 -1428 1294 -1422
rect 1236 -1462 1248 -1428
rect 1236 -1468 1294 -1462
rect 1236 -1640 1294 -1634
rect 1236 -1674 1248 -1640
rect 1236 -1680 1294 -1674
rect 1054 -1759 1107 -1723
rect 1423 -1776 1493 -1129
rect 1605 -1197 1663 -1191
rect 1605 -1231 1617 -1197
rect 1605 -1237 1663 -1231
rect 1605 -1391 1663 -1385
rect 1605 -1425 1617 -1391
rect 1605 -1431 1663 -1425
rect 1605 -1499 1663 -1493
rect 1605 -1533 1617 -1499
rect 1605 -1539 1663 -1533
rect 1605 -1693 1663 -1687
rect 1605 -1727 1617 -1693
rect 1605 -1733 1663 -1727
rect 1423 -1812 1476 -1776
rect 1794 -1829 1809 -1095
rect 1828 -1829 1862 -1041
rect 2144 -1129 2178 -1111
rect 1974 -1142 2032 -1136
rect 1974 -1176 1986 -1142
rect 2144 -1165 2214 -1129
rect 1974 -1182 2032 -1176
rect 2161 -1199 2232 -1165
rect 2512 -1199 2547 -1165
rect 1974 -1250 2032 -1244
rect 1974 -1284 1986 -1250
rect 1974 -1290 2032 -1284
rect 1974 -1444 2032 -1438
rect 1974 -1478 1986 -1444
rect 1974 -1484 2032 -1478
rect 1974 -1552 2032 -1546
rect 1974 -1586 1986 -1552
rect 1974 -1592 2032 -1586
rect 1974 -1746 2032 -1740
rect 1974 -1780 1986 -1746
rect 1974 -1786 2032 -1780
rect 1828 -1863 1843 -1829
rect 2161 -1882 2231 -1199
rect 2513 -1218 2547 -1199
rect 2343 -1267 2401 -1261
rect 2343 -1301 2355 -1267
rect 2343 -1307 2401 -1301
rect 2343 -1479 2401 -1473
rect 2343 -1513 2355 -1479
rect 2343 -1519 2401 -1513
rect 2343 -1587 2401 -1581
rect 2343 -1621 2355 -1587
rect 2343 -1627 2401 -1621
rect 2343 -1799 2401 -1793
rect 2343 -1833 2355 -1799
rect 2343 -1839 2401 -1833
rect 2161 -1918 2214 -1882
rect 2532 -1935 2547 -1218
rect 2566 -1252 2601 -1218
rect 2566 -1935 2600 -1252
rect 2882 -1271 2916 -1253
rect 2882 -1307 2952 -1271
rect 2712 -1320 2770 -1314
rect 2712 -1354 2724 -1320
rect 2899 -1341 2970 -1307
rect 3250 -1341 3285 -1307
rect 2712 -1360 2770 -1354
rect 2712 -1532 2770 -1526
rect 2712 -1566 2724 -1532
rect 2712 -1572 2770 -1566
rect 2712 -1640 2770 -1634
rect 2712 -1674 2724 -1640
rect 2712 -1680 2770 -1674
rect 2712 -1852 2770 -1846
rect 2712 -1886 2724 -1852
rect 2712 -1892 2770 -1886
rect 2566 -1969 2581 -1935
rect 2899 -1988 2969 -1341
rect 3251 -1360 3285 -1341
rect 3081 -1409 3139 -1403
rect 3081 -1443 3093 -1409
rect 3081 -1449 3139 -1443
rect 3081 -1603 3139 -1597
rect 3081 -1637 3093 -1603
rect 3081 -1643 3139 -1637
rect 3081 -1711 3139 -1705
rect 3081 -1745 3093 -1711
rect 3081 -1751 3139 -1745
rect 3081 -1905 3139 -1899
rect 3081 -1939 3093 -1905
rect 3081 -1945 3139 -1939
rect 2899 -2024 2952 -1988
rect 3270 -2041 3285 -1360
rect 3304 -1394 3339 -1360
rect 3304 -2041 3338 -1394
rect 3450 -1462 3508 -1456
rect 3450 -1496 3462 -1462
rect 3450 -1502 3508 -1496
rect 3450 -1656 3508 -1650
rect 3450 -1690 3462 -1656
rect 3450 -1696 3508 -1690
rect 3450 -1764 3508 -1758
rect 3450 -1798 3462 -1764
rect 3450 -1804 3508 -1798
rect 3450 -1958 3508 -1952
rect 3450 -1992 3462 -1958
rect 3450 -1998 3508 -1992
rect 3304 -2075 3319 -2041
rect 3639 -2094 3654 -1360
rect 3673 -2094 3707 -1306
rect 3673 -2128 3688 -2094
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
use sky130_fd_pr__cap_mim_m3_1_Z4YBWZ  XC1
timestamp 0
transform 1 0 6992 0 1 -6182
box -1886 -7440 1886 7440
use sky130_fd_pr__pfet_01v8_M47XPL  XM1
timestamp 0
transform 1 0 2372 0 1 -1550
box -211 -421 211 421
use sky130_fd_pr__pfet_01v8_M47XPL  XM2
timestamp 0
transform 1 0 2741 0 1 -1603
box -211 -421 211 421
use sky130_fd_pr__nfet_01v8_9XY3GD  XM3
timestamp 0
transform 1 0 2003 0 1 -1213
box -211 -705 211 705
use sky130_fd_pr__nfet_01v8_9XY3GD  XM4
timestamp 0
transform 1 0 4197 0 1 -1531
box -211 -705 211 705
use sky130_fd_pr__nfet_01v8_PTX3GD  XM5
timestamp 0
transform 1 0 896 0 1 -1356
box -211 -403 211 403
use sky130_fd_pr__nfet_01v8_PTX3GD  XM6
timestamp 0
transform 1 0 3110 0 1 -1674
box -211 -403 211 403
use sky130_fd_pr__nfet_01v8_PTX3GD  XM7
timestamp 0
transform 1 0 3479 0 1 -1727
box -211 -403 211 403
use sky130_fd_pr__pfet_01v8_M47T9Z  XM8
timestamp 0
transform 1 0 158 0 1 -912
box -211 -741 211 741
use sky130_fd_pr__pfet_01v8_M47T9Z  XM9
timestamp 0
transform 1 0 527 0 1 -965
box -211 -741 211 741
use sky130_fd_pr__pfet_01v8_M47T9Z  XM10
timestamp 0
transform 1 0 1265 0 1 -1071
box -211 -741 211 741
use sky130_fd_pr__nfet_01v8_PTX3GD  XM11
timestamp 0
transform 1 0 1634 0 1 -1462
box -211 -403 211 403
use sky130_fd_pr__res_high_po_0p35_K5HYSB  XR1
timestamp 0
transform 1 0 4556 0 1 -1407
box -201 -882 201 882
use sky130_fd_pr__res_high_po_0p35_K5HYSB  XR2
timestamp 0
transform 1 0 4905 0 1 -1460
box -201 -882 201 882
use sky130_fd_pr__res_high_po_0p35_K5HYSB  XR4
timestamp 0
transform 1 0 3838 0 1 -1301
box -201 -882 201 882
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 out
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 -
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 +
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 GND
port 4 nsew
<< end >>
