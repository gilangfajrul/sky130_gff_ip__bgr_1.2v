magic
tech sky130A
magscale 1 2
timestamp 1716303658
<< psubdiff >>
rect -239 616 -179 650
rect 8343 616 8403 650
rect -239 590 -205 616
rect 8369 590 8403 616
rect -239 -141 -205 -115
rect 8369 -141 8403 -115
rect -239 -175 -179 -141
rect 8343 -175 8403 -141
<< psubdiffcont >>
rect -179 616 8343 650
rect -239 -115 -205 590
rect 8369 -115 8403 590
rect -179 -175 8343 -141
<< poly >>
rect -93 316 -63 335
rect -170 268 -63 316
rect 1282 309 1995 335
rect 2053 309 2766 335
rect 8227 316 8257 335
rect 1282 265 1908 309
rect 2140 265 2766 309
rect 3314 268 3966 309
rect 4198 268 4824 309
rect 5398 265 6024 309
rect 6256 265 6882 309
rect 8227 268 8334 316
rect -170 160 -63 208
rect 1282 167 1908 211
rect 2140 167 2766 211
rect 3314 167 3966 208
rect 4198 167 4824 208
rect 5398 167 6024 211
rect 6256 167 6882 211
rect 1282 141 1995 167
rect 2053 141 2766 167
rect 8227 160 8334 208
rect 8227 141 8257 160
<< locali >>
rect -239 616 -179 650
rect 8343 616 8403 650
rect -239 590 -205 616
rect 8369 590 8403 616
rect -139 309 -105 335
rect 2007 331 2041 335
rect 8269 309 8303 335
rect -139 133 -105 167
rect 2007 141 2041 145
rect 8269 141 8303 167
rect -239 -141 -205 -115
rect 8369 -141 8403 -115
rect -239 -175 -179 -141
rect 8343 -175 8403 -141
<< viali >>
rect 1998 616 2050 650
rect 6114 616 6166 650
rect -239 275 -205 309
rect -157 275 -93 309
rect 1295 275 1895 309
rect 2153 275 2753 309
rect 3327 275 3953 309
rect 4211 275 4811 309
rect 5411 275 6011 309
rect 6269 275 6869 309
rect 8257 275 8321 309
rect 8369 275 8403 309
rect -239 167 -205 201
rect -157 167 -93 201
rect 1295 167 1895 201
rect 2153 167 2753 201
rect 3327 167 3953 201
rect 4211 167 4811 201
rect 5411 167 6011 201
rect 6269 167 6869 201
rect 8257 167 8321 201
rect 8369 167 8403 201
rect 1998 -175 2050 -141
rect 6114 -175 6166 -141
<< metal1 >>
rect 1988 656 1998 659
rect 1986 610 1998 656
rect 2050 656 2060 659
rect 6104 656 6114 659
rect 1988 607 1998 610
rect 2050 610 2062 656
rect 6102 610 6114 656
rect 6166 656 6176 659
rect 2050 607 2060 610
rect 6104 607 6114 610
rect 6166 610 6178 656
rect 6166 607 6176 610
rect -57 531 8221 579
rect -57 457 -11 531
rect 1988 347 1998 483
rect 2050 347 2060 483
rect 4059 442 4105 531
rect 6104 347 6114 483
rect 6166 347 6176 483
rect 8175 446 8221 531
rect -145 315 -99 335
rect -251 309 -81 315
rect -251 275 -239 309
rect -205 275 -157 309
rect -93 275 -81 309
rect -251 269 -81 275
rect 1283 266 1295 318
rect 1895 266 1907 318
rect -251 201 -81 207
rect -251 167 -239 201
rect -205 167 -157 201
rect -93 167 -81 201
rect -251 161 -81 167
rect -145 135 -99 161
rect 1283 158 1295 210
rect 1895 158 1907 210
rect 2001 141 2047 335
rect 2141 266 2153 318
rect 2753 266 2765 318
rect 3315 309 3965 315
rect 3315 275 3327 309
rect 3953 307 3965 309
rect 4199 309 4823 315
rect 4199 307 4211 309
rect 3953 275 4211 307
rect 4811 275 4823 309
rect 3315 267 4823 275
rect 5399 266 5411 318
rect 6011 266 6023 318
rect 2141 158 2153 210
rect 2753 158 2765 210
rect 3315 201 4823 209
rect 3315 167 3327 201
rect 3953 169 4211 201
rect 3953 167 3965 169
rect 3315 161 3965 167
rect 4199 167 4211 169
rect 4811 167 4823 201
rect 4199 161 4823 167
rect 5399 158 5411 210
rect 6011 158 6023 210
rect 6117 132 6163 347
rect 6257 266 6269 318
rect 6869 266 6881 318
rect 8263 315 8309 335
rect 8245 309 8415 315
rect 8245 275 8257 309
rect 8321 275 8369 309
rect 8403 275 8415 309
rect 8245 269 8415 275
rect 6257 158 6269 210
rect 6869 158 6881 210
rect 8245 201 8415 207
rect 8245 167 8257 201
rect 8321 167 8369 201
rect 8403 167 8415 201
rect 8245 161 8415 167
rect 8263 141 8309 161
rect 6117 130 6163 131
rect -57 -56 -11 29
rect 1988 -7 1998 129
rect 2050 -7 2060 129
rect 4059 -56 4105 66
rect 6104 -7 6114 129
rect 6166 -7 6176 129
rect 8175 -56 8221 18
rect -57 -104 8221 -56
rect 1988 -135 1998 -132
rect 1986 -181 1998 -135
rect 2050 -135 2060 -132
rect 6104 -135 6114 -132
rect 1988 -184 1998 -181
rect 2050 -181 2062 -135
rect 6102 -181 6114 -135
rect 6166 -135 6176 -132
rect 2050 -184 2060 -181
rect 6104 -184 6114 -181
rect 6166 -181 6178 -135
rect 6166 -184 6176 -181
<< via1 >>
rect 1998 650 2050 659
rect 1998 616 2050 650
rect 1998 607 2050 616
rect 6114 650 6166 659
rect 6114 616 6166 650
rect 6114 607 6166 616
rect 1998 347 2050 483
rect 6114 347 6166 483
rect 1295 309 1895 318
rect 1295 275 1895 309
rect 1295 266 1895 275
rect 1295 201 1895 210
rect 1295 167 1895 201
rect 1295 158 1895 167
rect 2153 309 2753 318
rect 2153 275 2753 309
rect 2153 266 2753 275
rect 5411 309 6011 318
rect 5411 275 6011 309
rect 5411 266 6011 275
rect 2153 201 2753 210
rect 2153 167 2753 201
rect 2153 158 2753 167
rect 5411 201 6011 210
rect 5411 167 6011 201
rect 5411 158 6011 167
rect 6269 309 6869 318
rect 6269 275 6869 309
rect 6269 266 6869 275
rect 6269 201 6869 210
rect 6269 167 6869 201
rect 6269 158 6869 167
rect 1998 -7 2050 129
rect 6114 -7 6166 129
rect 1998 -141 2050 -132
rect 1998 -175 2050 -141
rect 1998 -184 2050 -175
rect 6114 -141 6166 -132
rect 6114 -175 6166 -141
rect 6114 -184 6166 -175
<< metal2 >>
rect 1998 659 2050 669
rect 1998 483 2050 607
rect 1998 337 2050 347
rect 6114 659 6166 669
rect 6114 483 6166 607
rect 6114 337 6166 347
rect 1295 320 1895 330
rect 2153 318 2753 328
rect 1295 254 1895 264
rect 2007 275 2153 309
rect 1295 210 1895 220
rect 2007 201 2041 275
rect 2153 256 2753 266
rect 5411 318 6011 328
rect 6269 320 6869 330
rect 6011 275 6157 309
rect 5411 256 6011 266
rect 1895 167 2041 201
rect 2153 212 2753 222
rect 1295 148 1895 158
rect 2153 146 2753 156
rect 5411 212 6011 222
rect 6123 201 6157 275
rect 6269 254 6869 264
rect 6269 210 6869 220
rect 6123 167 6269 201
rect 5411 146 6011 156
rect 6269 148 6869 158
rect 1998 129 2050 139
rect 1998 -132 2050 -7
rect 1998 -194 2050 -184
rect 6114 129 6166 139
rect 6114 -132 6166 -7
rect 6114 -194 6166 -184
<< via2 >>
rect 1295 318 1895 320
rect 1295 266 1895 318
rect 1295 264 1895 266
rect 6269 318 6869 320
rect 2153 210 2753 212
rect 2153 158 2753 210
rect 2153 156 2753 158
rect 5411 210 6011 212
rect 5411 158 6011 210
rect 6269 266 6869 318
rect 6269 264 6869 266
rect 5411 156 6011 158
<< metal3 >>
rect 1285 323 1905 325
rect 6259 323 6879 325
rect 1285 320 2055 323
rect 1285 264 1295 320
rect 1895 264 2055 320
rect 1285 261 2055 264
rect 1285 259 1905 261
rect 1993 215 2055 261
rect 6109 320 6879 323
rect 6109 264 6269 320
rect 6869 264 6879 320
rect 6109 261 6879 264
rect 2143 215 2763 217
rect 1993 212 2763 215
rect 1993 156 2153 212
rect 2753 156 2763 212
rect 1993 153 2763 156
rect 2143 151 2763 153
rect 5401 215 6021 217
rect 6109 215 6171 261
rect 6259 259 6879 261
rect 5401 212 6171 215
rect 5401 156 5411 212
rect 6011 156 6171 212
rect 5401 153 6171 156
rect 5401 151 6021 153
use sky130_fd_pr__nfet_01v8_4VSDG9  sky130_fd_pr__nfet_01v8_4VSDG9_0
timestamp 1716303658
transform 1 0 -78 0 1 415
box -73 -106 73 106
use sky130_fd_pr__nfet_01v8_4VSDG9  sky130_fd_pr__nfet_01v8_4VSDG9_1
timestamp 1716303658
transform 1 0 8242 0 1 415
box -73 -106 73 106
use sky130_fd_pr__nfet_01v8_4VSDG9  sky130_fd_pr__nfet_01v8_4VSDG9_2
timestamp 1716303658
transform 1 0 8242 0 1 61
box -73 -106 73 106
use sky130_fd_pr__nfet_01v8_4VSDG9  sky130_fd_pr__nfet_01v8_4VSDG9_3
timestamp 1716303658
transform 1 0 -78 0 1 61
box -73 -106 73 106
use sky130_fd_pr__nfet_01v8_EDB9KC  sky130_fd_pr__nfet_01v8_EDB9KC_0
timestamp 1716303658
transform 1 0 148 0 1 207
box 0 0 1 1
use sky130_fd_pr__nfet_01v8_X627NV  sky130_fd_pr__nfet_01v8_X627NV_0
timestamp 1716303658
transform -1 0 4082 0 1 415
box -4145 -106 4145 106
use sky130_fd_pr__nfet_01v8_X627NV  sky130_fd_pr__nfet_01v8_X627NV_1
timestamp 1716303658
transform -1 0 4082 0 1 61
box -4145 -106 4145 106
<< end >>
