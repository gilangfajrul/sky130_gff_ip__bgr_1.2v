magic
tech sky130A
magscale 1 2
timestamp 1720118050
<< psubdiff >>
rect -309 1533 -249 1567
rect 8527 1533 8587 1567
rect -309 1485 -275 1533
rect 8553 1485 8587 1533
rect -309 -95 -275 -69
rect 8553 -95 8587 -69
rect -309 -129 -249 -95
rect 8527 -129 8587 -95
<< psubdiffcont >>
rect -249 1533 8527 1567
rect -309 -69 -275 1485
rect 8553 -69 8587 1485
rect -249 -129 8527 -95
<< poly >>
rect -208 1482 -116 1498
rect -208 1448 -192 1482
rect -158 1448 -116 1482
rect -208 1432 -116 1448
rect 8394 1482 8486 1498
rect 8394 1448 8436 1482
rect 8470 1448 8486 1482
rect 8394 1432 8486 1448
rect -208 1088 -116 1104
rect -208 1054 -192 1088
rect -158 1054 -116 1088
rect -208 1038 -116 1054
rect 54 1042 8224 1185
rect 8394 1088 8486 1104
rect 8394 1054 8436 1088
rect 8470 1054 8486 1088
rect 8394 1038 8486 1054
rect 54 648 8224 791
rect -208 384 -116 400
rect -208 350 -192 384
rect -158 350 -116 384
rect -208 334 -116 350
rect 54 254 8224 397
rect 8394 384 8486 400
rect 8394 350 8436 384
rect 8470 350 8486 384
rect 8394 334 8486 350
rect -146 6 -116 7
rect -208 -10 -116 6
rect -208 -44 -192 -10
rect -158 -44 -116 -10
rect -208 -60 -116 -44
rect 8394 -10 8486 6
rect 8394 -44 8436 -10
rect 8470 -44 8486 -10
rect 8394 -60 8486 -44
<< polycont >>
rect -192 1448 -158 1482
rect 8436 1448 8470 1482
rect -192 1054 -158 1088
rect 8436 1054 8470 1088
rect -192 350 -158 384
rect 8436 350 8470 384
rect -192 -44 -158 -10
rect 8436 -44 8470 -10
<< locali >>
rect -192 1482 -158 1498
rect -192 1411 -158 1448
rect 8436 1482 8470 1498
rect -104 1398 -70 1411
rect 8436 1408 8470 1448
rect -192 1088 -158 1104
rect -192 1013 -158 1054
rect 8436 1088 8470 1104
rect 8436 1007 8470 1054
rect -192 384 -158 425
rect -192 334 -158 350
rect 8436 384 8470 444
rect 8436 334 8470 350
rect -192 -10 -158 34
rect -192 -60 -158 -44
rect 8436 -10 8470 46
rect 8436 -60 8470 -44
<< viali >>
rect -309 1533 -249 1567
rect -249 1533 8527 1567
rect 8527 1533 8587 1567
rect -309 1485 -275 1533
rect -309 -69 -275 1485
rect -192 1448 -158 1482
rect 8436 1448 8470 1482
rect 8553 1485 8587 1533
rect -192 1054 -158 1088
rect 8436 1054 8470 1088
rect -192 350 -158 384
rect 8436 350 8470 384
rect -192 -44 -158 -10
rect 8436 -44 8470 -10
rect -309 -95 -275 -69
rect 8553 -69 8587 1485
rect 8553 -95 8587 -69
rect -309 -129 -249 -95
rect -249 -129 8527 -95
rect 8527 -129 8587 -95
<< metal1 >>
rect -315 1573 -269 1579
rect 4060 1573 4106 1579
rect 8547 1573 8593 1579
rect -321 1567 8599 1573
rect -321 1527 -309 1567
rect -315 -89 -309 1527
rect -321 -129 -309 -89
rect -275 1527 8553 1533
rect -275 -89 -269 1527
rect -198 1482 -152 1494
rect -198 1448 -192 1482
rect -158 1448 -152 1482
rect -198 1410 -152 1448
rect 8 1443 1089 1489
rect 8 1410 42 1443
rect -198 1406 48 1410
rect -164 1210 48 1406
rect 4060 1405 4106 1527
rect 8430 1482 8476 1494
rect 8430 1448 8436 1482
rect 8470 1448 8476 1482
rect 8430 1410 8476 1448
rect 8230 1406 8476 1410
rect 8230 1398 8461 1406
rect -198 1088 -152 1100
rect -198 1054 -192 1088
rect -158 1054 -152 1088
rect -198 1016 -152 1054
rect 4060 1016 4106 1227
rect 4153 1222 4163 1398
rect 4227 1222 4237 1398
rect 8230 1222 8283 1398
rect 8335 1222 8461 1398
rect 8230 1210 8461 1222
rect 8430 1088 8476 1100
rect 8430 1054 8436 1088
rect 8470 1054 8476 1088
rect 8430 1016 8476 1054
rect -198 1012 48 1016
rect -161 1004 48 1012
rect -161 828 -57 1004
rect -5 828 48 1004
rect -161 816 48 828
rect -165 610 48 622
rect -165 434 -57 610
rect -5 434 48 610
rect -165 428 48 434
rect -198 422 48 428
rect 4060 450 4217 1016
rect 8230 1011 8476 1016
rect 8230 1004 8474 1011
rect 8230 828 8283 1004
rect 8335 828 8474 1004
rect 8230 816 8474 828
rect 8230 610 8464 622
rect 4060 422 4218 450
rect 8230 434 8283 610
rect 8335 436 8464 610
rect 8335 434 8476 436
rect 8230 422 8476 434
rect -198 384 -152 422
rect -198 350 -192 384
rect -158 350 -152 384
rect -198 338 -152 350
rect -177 216 48 228
rect 4172 216 4218 422
rect 8430 384 8476 422
rect 8430 350 8436 384
rect 8470 350 8476 384
rect 8430 338 8476 350
rect -177 40 -57 216
rect -5 40 48 216
rect 4041 40 4051 216
rect 4115 40 4125 216
rect 8230 41 8441 228
rect -177 38 48 40
rect -198 28 48 38
rect -198 -10 -152 28
rect -198 -44 -192 -10
rect -158 -44 -152 -10
rect -198 -56 -152 -44
rect 4172 -89 4218 40
rect 8230 28 8476 41
rect 8236 -3 8270 28
rect 7161 -49 8270 -3
rect 8430 -10 8476 28
rect 8430 -44 8436 -10
rect 8470 -44 8476 -10
rect 8430 -56 8476 -44
rect 8547 -89 8553 1527
rect -275 -95 8553 -89
rect 8587 1527 8599 1567
rect 8587 -89 8593 1527
rect 8587 -129 8599 -89
rect -321 -135 8599 -129
rect -315 -141 -269 -135
rect 4172 -141 4218 -135
rect 8547 -141 8593 -135
<< via1 >>
rect 4163 1222 4227 1398
rect 8283 1222 8335 1398
rect -57 828 -5 1004
rect -57 434 -5 610
rect 8283 828 8335 1004
rect 8283 434 8335 610
rect -57 40 -5 216
rect 4051 40 4115 216
<< metal2 >>
rect 4163 1398 4227 1408
rect 4163 1212 4227 1222
rect 8283 1398 8335 1408
rect 8283 1139 8335 1222
rect -270 1087 8548 1139
rect -270 351 -218 1087
rect -57 1004 -5 1014
rect -57 745 -5 828
rect 8281 1004 8337 1014
rect 8281 818 8337 828
rect -57 693 8335 745
rect -59 610 -3 620
rect -59 424 -3 434
rect 8283 610 8335 693
rect 8283 424 8335 434
rect 8496 351 8548 1087
rect -270 299 8548 351
rect -57 216 -5 299
rect -57 30 -5 40
rect 4051 216 4115 226
rect 4051 30 4115 40
<< via2 >>
rect 4163 1222 4227 1398
rect 8281 828 8283 1004
rect 8283 828 8335 1004
rect 8335 828 8337 1004
rect -59 434 -57 610
rect -57 434 -5 610
rect -5 434 -3 610
rect 4051 40 4115 216
<< metal3 >>
rect 4153 1398 4237 1403
rect 4153 1222 4163 1398
rect 4227 1222 4237 1398
rect 4153 1217 4237 1222
rect 8271 1004 8347 1009
rect 8271 828 8281 1004
rect 8337 828 8347 1004
rect 8271 823 8347 828
rect 8279 749 8339 823
rect -61 689 8339 749
rect -61 615 -1 689
rect -69 610 7 615
rect -69 434 -59 610
rect -3 434 7 610
rect -69 429 7 434
rect 4041 216 4125 221
rect 4041 40 4051 216
rect 4115 40 4125 216
rect 4041 35 4125 40
<< via3 >>
rect 4163 1222 4227 1398
rect 4051 40 4115 216
<< metal4 >>
rect 4106 1398 4228 1399
rect 4106 1222 4163 1398
rect 4227 1222 4228 1398
rect 4106 1221 4228 1222
rect 4106 217 4172 1221
rect 4050 216 4172 217
rect 4050 40 4051 216
rect 4115 40 4172 216
rect 4050 39 4172 40
use sky130_fd_pr__nfet_01v8_3KF9AC  sky130_fd_pr__nfet_01v8_3KF9AC_0
timestamp 1717076529
transform 1 0 2054 0 1 1341
box -2058 -157 2058 157
use sky130_fd_pr__nfet_01v8_3YKU97  sky130_fd_pr__nfet_01v8_3YKU97_0
timestamp 1717076529
transform 1 0 6224 0 1 97
box -2058 -157 2058 157
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_0
timestamp 1717432527
transform 1 0 -131 0 1 916
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_1
timestamp 1717432527
transform 1 0 -131 0 1 1310
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_2
timestamp 1717432527
transform 1 0 -131 0 1 522
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_3
timestamp 1717432527
transform 1 0 -131 0 1 128
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_4
timestamp 1717432527
transform 1 0 8409 0 1 128
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_5
timestamp 1717432527
transform 1 0 8409 0 1 522
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_6
timestamp 1717432527
transform 1 0 8409 0 1 916
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_7
timestamp 1717432527
transform 1 0 8409 0 1 1310
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_BSRS8Q  sky130_fd_pr__nfet_01v8_BSRS8Q_0
timestamp 1717249617
transform 1 0 6224 0 1 1310
box -2058 -126 2058 126
use sky130_fd_pr__nfet_01v8_P5G96Q  sky130_fd_pr__nfet_01v8_P5G96Q_1
timestamp 1716212328
transform 1 0 2054 0 1 128
box -2058 -126 2058 126
use sky130_fd_pr__nfet_01v8_P5G96Q  sky130_fd_pr__nfet_01v8_P5G96Q_4
timestamp 1716212328
transform 1 0 6224 0 1 522
box -2058 -126 2058 126
use sky130_fd_pr__nfet_01v8_P5G96Q  sky130_fd_pr__nfet_01v8_P5G96Q_5
timestamp 1716212328
transform 1 0 2054 0 1 522
box -2058 -126 2058 126
use sky130_fd_pr__nfet_01v8_P5G96Q  sky130_fd_pr__nfet_01v8_P5G96Q_6
timestamp 1716212328
transform 1 0 6224 0 1 916
box -2058 -126 2058 126
use sky130_fd_pr__nfet_01v8_P5G96Q  sky130_fd_pr__nfet_01v8_P5G96Q_7
timestamp 1716212328
transform 1 0 2054 0 1 916
box -2058 -126 2058 126
<< labels >>
flabel metal2 8302 652 8302 652 0 FreeSans 160 0 0 0 D3
port 2 nsew
flabel metal3 8310 784 8310 784 0 FreeSans 160 0 0 0 D4
port 1 nsew
flabel metal2 8306 1160 8306 1160 0 FreeSans 160 0 0 0 D1
port 0 nsew
flabel metal4 4136 80 4136 80 0 FreeSans 160 0 0 0 S2
port 5 nsew
flabel metal1 8562 -136 8562 -136 0 FreeSans 160 0 0 0 AVSS
port 6 nsew
flabel metal1 8310 134 8310 134 0 FreeSans 160 0 0 0 D2
port 3 nsew
<< end >>
