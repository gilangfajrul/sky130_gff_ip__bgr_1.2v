magic
tech sky130A
magscale 1 2
timestamp 1716351939
<< xpolycontact >>
rect -654 590 -516 1022
rect -654 52 -516 484
rect -420 590 -282 1022
rect -420 52 -282 484
rect -186 590 -48 1022
rect -186 52 -48 484
rect 48 590 186 1022
rect 48 52 186 484
rect 282 590 420 1022
rect 282 52 420 484
rect 516 590 654 1022
rect 516 52 654 484
rect -654 -484 -516 -52
rect -654 -1022 -516 -590
rect -420 -484 -282 -52
rect -420 -1022 -282 -590
rect -186 -484 -48 -52
rect -186 -1022 -48 -590
rect 48 -484 186 -52
rect 48 -1022 186 -590
rect 282 -484 420 -52
rect 282 -1022 420 -590
rect 516 -484 654 -52
rect 516 -1022 654 -590
<< ppolyres >>
rect -654 484 -516 590
rect -420 484 -282 590
rect -186 484 -48 590
rect 48 484 186 590
rect 282 484 420 590
rect 516 484 654 590
rect -654 -590 -516 -484
rect -420 -590 -282 -484
rect -186 -590 -48 -484
rect 48 -590 186 -484
rect 282 -590 420 -484
rect 516 -590 654 -484
<< viali >>
rect -638 607 -532 1004
rect -404 607 -298 1004
rect -170 607 -64 1004
rect 64 607 170 1004
rect 298 607 404 1004
rect 532 607 638 1004
rect -638 70 -532 467
rect -404 70 -298 467
rect -170 70 -64 467
rect 64 70 170 467
rect 298 70 404 467
rect 532 70 638 467
rect -638 -467 -532 -70
rect -404 -467 -298 -70
rect -170 -467 -64 -70
rect 64 -467 170 -70
rect 298 -467 404 -70
rect 532 -467 638 -70
rect -638 -1004 -532 -607
rect -404 -1004 -298 -607
rect -170 -1004 -64 -607
rect 64 -1004 170 -607
rect 298 -1004 404 -607
rect 532 -1004 638 -607
<< metal1 >>
rect -644 1004 -526 1016
rect -644 607 -638 1004
rect -532 607 -526 1004
rect -644 595 -526 607
rect -410 1004 -292 1016
rect -410 607 -404 1004
rect -298 607 -292 1004
rect -410 595 -292 607
rect -176 1004 -58 1016
rect -176 607 -170 1004
rect -64 607 -58 1004
rect -176 595 -58 607
rect 58 1004 176 1016
rect 58 607 64 1004
rect 170 607 176 1004
rect 58 595 176 607
rect 292 1004 410 1016
rect 292 607 298 1004
rect 404 607 410 1004
rect 292 595 410 607
rect 526 1004 644 1016
rect 526 607 532 1004
rect 638 607 644 1004
rect 526 595 644 607
rect -644 467 -526 479
rect -644 70 -638 467
rect -532 70 -526 467
rect -644 58 -526 70
rect -410 467 -292 479
rect -410 70 -404 467
rect -298 70 -292 467
rect -410 58 -292 70
rect -176 467 -58 479
rect -176 70 -170 467
rect -64 70 -58 467
rect -176 58 -58 70
rect 58 467 176 479
rect 58 70 64 467
rect 170 70 176 467
rect 58 58 176 70
rect 292 467 410 479
rect 292 70 298 467
rect 404 70 410 467
rect 292 58 410 70
rect 526 467 644 479
rect 526 70 532 467
rect 638 70 644 467
rect 526 58 644 70
rect -644 -70 -526 -58
rect -644 -467 -638 -70
rect -532 -467 -526 -70
rect -644 -479 -526 -467
rect -410 -70 -292 -58
rect -410 -467 -404 -70
rect -298 -467 -292 -70
rect -410 -479 -292 -467
rect -176 -70 -58 -58
rect -176 -467 -170 -70
rect -64 -467 -58 -70
rect -176 -479 -58 -467
rect 58 -70 176 -58
rect 58 -467 64 -70
rect 170 -467 176 -70
rect 58 -479 176 -467
rect 292 -70 410 -58
rect 292 -467 298 -70
rect 404 -467 410 -70
rect 292 -479 410 -467
rect 526 -70 644 -58
rect 526 -467 532 -70
rect 638 -467 644 -70
rect 526 -479 644 -467
rect -644 -607 -526 -595
rect -644 -1004 -638 -607
rect -532 -1004 -526 -607
rect -644 -1016 -526 -1004
rect -410 -607 -292 -595
rect -410 -1004 -404 -607
rect -298 -1004 -292 -607
rect -410 -1016 -292 -1004
rect -176 -607 -58 -595
rect -176 -1004 -170 -607
rect -64 -1004 -58 -607
rect -176 -1016 -58 -1004
rect 58 -607 176 -595
rect 58 -1004 64 -607
rect 170 -1004 176 -607
rect 58 -1016 176 -1004
rect 292 -607 410 -595
rect 292 -1004 298 -607
rect 404 -1004 410 -607
rect 292 -1016 410 -1004
rect 526 -607 644 -595
rect 526 -1004 532 -607
rect 638 -1004 644 -607
rect 526 -1016 644 -1004
<< properties >>
string gencell sky130_fd_pr__res_high_po_0p69
string library sky130
string parameters w 0.690 l 0.69 m 2 nx 6 wmin 0.690 lmin 0.50 rho 319.8 val 884.495 dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.690 n_guard 1 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
