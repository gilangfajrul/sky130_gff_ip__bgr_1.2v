magic
tech sky130A
magscale 1 2
timestamp 1716998311
<< nwell >>
rect -177 -62 4422 780
<< nsubdiff >>
rect -141 710 -81 744
rect 4326 710 4386 744
rect -141 684 -107 710
rect 4352 684 4386 710
rect -141 8 -107 34
rect 4352 8 4386 34
rect -141 -26 -81 8
rect 4326 -26 4386 8
<< nsubdiffcont >>
rect -81 710 4326 744
rect -141 34 -107 684
rect 4352 34 4386 684
rect -81 -26 4326 8
<< poly >>
rect -41 395 36 431
rect 593 395 1595 430
rect 2651 395 3653 430
rect 4210 395 4287 431
rect -41 287 36 323
rect 2651 288 3653 323
rect 4210 287 4287 323
<< locali >>
rect -141 710 -81 744
rect 4326 710 4386 744
rect -141 684 -107 710
rect 4352 684 4386 710
rect -40 430 -6 471
rect 4252 430 4286 470
rect -40 254 -6 288
rect 4252 249 4286 288
rect -141 8 -107 34
rect 4352 8 4386 34
rect -141 -26 -81 8
rect 4326 -26 4386 8
<< viali >>
rect 2106 710 2140 744
rect -141 396 -107 430
rect -40 396 -6 430
rect 594 396 1594 430
rect 2652 396 3652 430
rect 4252 396 4286 430
rect 4352 396 4386 430
rect -141 288 -107 322
rect -40 288 -6 322
rect 594 288 1594 322
rect 2652 288 3652 322
rect 4252 288 4286 322
rect 4352 288 4386 322
rect 2106 -26 2140 8
<< metal1 >>
rect 2094 744 2152 750
rect 2094 710 2106 744
rect 2140 710 2152 744
rect 2094 704 2152 710
rect 2100 655 2146 704
rect 2087 468 2097 644
rect 2149 468 2159 644
rect -46 436 0 463
rect -153 430 6 436
rect -153 396 -141 430
rect -107 396 -40 430
rect -6 396 6 430
rect -153 390 6 396
rect 42 428 88 464
rect 582 430 1606 436
rect 582 428 594 430
rect 42 396 594 428
rect 1594 428 1606 430
rect 2640 430 3664 436
rect 2640 428 2652 430
rect 1594 396 2652 428
rect 3652 396 3664 430
rect 4158 428 4204 456
rect 4246 436 4292 463
rect 42 382 3664 396
rect 3908 382 4204 428
rect 4240 430 4398 436
rect 4240 396 4252 430
rect 4286 396 4352 430
rect 4386 396 4398 430
rect 4240 390 4398 396
rect 3908 336 3954 382
rect -153 322 1606 328
rect -153 288 -141 322
rect -107 288 -40 322
rect -6 288 594 322
rect 1594 288 1606 322
rect -153 282 1606 288
rect 2640 322 3954 336
rect 2640 288 2652 322
rect 3652 290 3954 322
rect 4240 322 4398 328
rect 3652 288 3664 290
rect 2640 282 3664 288
rect 4240 288 4252 322
rect 4286 288 4352 322
rect 4386 288 4398 322
rect 4240 282 4398 288
rect -46 254 0 282
rect 42 246 88 282
rect 4246 250 4292 282
rect 2087 74 2097 250
rect 2149 74 2159 250
rect 2100 14 2146 72
rect 2094 8 2152 14
rect 2094 -26 2106 8
rect 2140 -26 2152 8
rect 2094 -32 2152 -26
<< via1 >>
rect 2097 468 2149 644
rect 2097 74 2149 250
<< metal2 >>
rect 2097 644 2149 654
rect 2097 250 2149 468
rect 2097 64 2149 74
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_0
timestamp 1716916329
transform 1 0 4225 0 1 162
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_1
timestamp 1716916329
transform 1 0 21 0 1 162
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_2
timestamp 1716916329
transform 1 0 21 0 1 556
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_3
timestamp 1716916329
transform 1 0 4225 0 1 556
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_UK88DC  sky130_fd_pr__pfet_01v8_UK88DC_0
timestamp 1716916205
transform 1 0 2123 0 1 556
box -2123 -162 2123 162
use sky130_fd_pr__pfet_01v8_UK88DC  sky130_fd_pr__pfet_01v8_UK88DC_1
timestamp 1716916205
transform 1 0 2123 0 1 162
box -2123 -162 2123 162
<< end >>
