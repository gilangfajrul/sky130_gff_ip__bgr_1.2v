magic
tech sky130A
magscale 1 2
timestamp 1762753955
<< nwell >>
rect -227 -676 8487 506
<< nsubdiff >>
rect -191 436 -131 470
rect 8391 436 8451 470
rect -191 410 -157 436
rect 8417 410 8451 436
rect -191 -606 -157 -580
rect 8417 -606 8451 -580
rect -191 -640 -131 -606
rect 8391 -640 8451 -606
<< nsubdiffcont >>
rect -131 436 8391 470
rect -191 -580 -157 410
rect 8417 -580 8451 410
rect -131 -640 8391 -606
<< poly >>
rect -86 393 -15 409
rect -86 359 -70 393
rect -36 359 -15 393
rect -86 343 -15 359
rect -45 312 -15 343
rect 8275 393 8346 409
rect 8275 359 8296 393
rect 8330 359 8346 393
rect 8275 343 8346 359
rect 8275 312 8305 343
rect -45 -513 -15 -489
rect -86 -529 -15 -513
rect -86 -563 -70 -529
rect -36 -563 -15 -529
rect -86 -579 -15 -563
rect 8275 -513 8305 -491
rect 8275 -529 8346 -513
rect 8275 -563 8296 -529
rect 8330 -563 8346 -529
rect 8275 -579 8346 -563
<< polycont >>
rect -70 359 -36 393
rect 8296 359 8330 393
rect -70 -563 -36 -529
rect 8296 -563 8330 -529
<< locali >>
rect -86 359 -70 393
rect -36 359 -20 393
rect 8280 359 8296 393
rect 8330 359 8346 393
rect -86 -563 -70 -529
rect -36 -563 -20 -529
rect 8280 -563 8296 -529
rect 8330 -563 8346 -529
<< viali >>
rect -191 436 -131 470
rect -131 436 8391 470
rect 8391 436 8451 470
rect -191 410 -157 436
rect -191 -580 -157 410
rect 8417 410 8451 436
rect -70 359 -36 393
rect 8296 359 8330 393
rect -70 -563 -36 -529
rect 8296 -563 8330 -529
rect -191 -606 -157 -580
rect 8417 -580 8451 410
rect 8417 -606 8451 -580
rect -191 -640 -131 -606
rect -131 -640 8391 -606
rect 8391 -640 8451 -606
<< metal1 >>
rect -197 476 -151 482
rect 2040 476 2046 479
rect -203 470 2046 476
rect 2098 476 2104 479
rect 6156 476 6162 479
rect 2098 470 6162 476
rect 6214 476 6220 479
rect 8411 476 8457 482
rect 6214 470 8463 476
rect -203 430 -191 470
rect -197 -600 -191 430
rect -203 -640 -191 -600
rect -157 430 2046 436
rect -157 -600 -151 430
rect 2040 427 2046 430
rect 2098 430 6162 436
rect 2098 427 2104 430
rect 6156 427 6162 430
rect 6214 430 8417 436
rect 6214 427 6220 430
rect -97 393 -24 399
rect -97 359 -70 393
rect -36 359 -24 393
rect -97 353 -24 359
rect 8284 393 8357 399
rect 8284 359 8296 393
rect 8330 359 8357 393
rect 8284 353 8357 359
rect -97 300 -51 353
rect 8311 300 8357 353
rect -97 295 -12 300
rect -83 124 -12 295
rect 40 124 50 300
rect 2036 124 2046 300
rect 2098 124 2108 300
rect 4094 124 4104 300
rect 4156 124 4166 300
rect 6152 124 6162 300
rect 6214 124 6224 300
rect 8210 124 8220 300
rect 8272 286 8357 300
rect 8272 124 8347 286
rect -101 22 -95 74
rect -43 71 -37 74
rect 8294 71 8300 74
rect -43 25 76 71
rect 8185 25 8300 71
rect -43 22 -37 25
rect 8294 22 8300 25
rect 8352 22 8358 74
rect -22 -61 -12 -9
rect 40 -61 4208 -9
rect 4260 -61 8220 -9
rect 8272 -61 8282 -9
rect -12 -109 40 -103
rect -22 -161 -12 -109
rect 40 -161 4000 -109
rect 4052 -161 8220 -109
rect 8272 -161 8282 -109
rect -12 -167 40 -161
rect -101 -244 -95 -192
rect -43 -195 -37 -192
rect 8294 -195 8300 -192
rect -43 -241 92 -195
rect 8204 -241 8300 -195
rect -43 -244 -37 -241
rect 8294 -244 8300 -241
rect 8352 -244 8358 -192
rect -89 -448 -12 -294
rect -97 -470 -12 -448
rect 40 -470 50 -294
rect 2036 -470 2046 -294
rect 2098 -470 2108 -294
rect 4094 -470 4104 -294
rect 4156 -470 4166 -294
rect 6152 -470 6162 -294
rect 6214 -470 6224 -294
rect 8210 -470 8220 -294
rect 8272 -470 8357 -294
rect -97 -523 -51 -470
rect 8311 -523 8357 -470
rect -97 -529 -24 -523
rect -97 -563 -70 -529
rect -36 -563 -24 -529
rect -97 -569 -24 -563
rect 8284 -529 8357 -523
rect 8284 -563 8296 -529
rect 8330 -563 8357 -529
rect 8284 -569 8357 -563
rect 2040 -600 2046 -597
rect -157 -606 2046 -600
rect 2098 -600 2104 -597
rect 6156 -600 6162 -597
rect 2098 -606 6162 -600
rect 6214 -600 6220 -597
rect 8411 -600 8417 430
rect 6214 -606 8417 -600
rect 8451 430 8463 470
rect 8451 -600 8457 430
rect 8451 -640 8463 -600
rect -203 -646 2046 -640
rect -197 -652 -151 -646
rect 2040 -649 2046 -646
rect 2098 -646 6162 -640
rect 2098 -649 2104 -646
rect 6156 -649 6162 -646
rect 6214 -646 8463 -640
rect 6214 -649 6220 -646
rect 8411 -652 8457 -646
<< via1 >>
rect 2046 470 2098 479
rect 6162 470 6214 479
rect 2046 436 2098 470
rect 6162 436 6214 470
rect 2046 427 2098 436
rect 6162 427 6214 436
rect -12 124 40 300
rect 2046 124 2098 300
rect 4104 124 4156 300
rect 6162 124 6214 300
rect 8220 124 8272 300
rect -95 22 -43 74
rect 8300 22 8352 74
rect -12 -61 40 -9
rect 4208 -61 4260 -9
rect 8220 -61 8272 -9
rect -12 -161 40 -109
rect 4000 -161 4052 -109
rect 8220 -161 8272 -109
rect -95 -244 -43 -192
rect 8300 -244 8352 -192
rect -12 -470 40 -294
rect 2046 -470 2098 -294
rect 4104 -470 4156 -294
rect 6162 -470 6214 -294
rect 8220 -470 8272 -294
rect 2046 -606 2098 -597
rect 6162 -606 6214 -597
rect 2046 -640 2098 -606
rect 6162 -640 6214 -606
rect 2046 -649 2098 -640
rect 6162 -649 6214 -640
<< metal2 >>
rect 2046 479 2098 485
rect -12 300 40 310
rect -95 74 -43 80
rect -95 16 -43 22
rect -92 -186 -46 16
rect -12 -9 40 124
rect -12 -71 40 -61
rect 2046 300 2098 427
rect 6162 479 6214 485
rect -12 -109 40 -99
rect -18 -161 -12 -109
rect 40 -161 46 -109
rect -95 -192 -43 -186
rect -95 -250 -43 -244
rect -12 -294 40 -161
rect -12 -480 40 -470
rect 2046 -294 2098 124
rect 4104 300 4156 310
rect 4104 -9 4156 124
rect 6162 300 6214 427
rect 4000 -61 4156 -9
rect 4208 -9 4260 3
rect 4000 -109 4052 -61
rect 4208 -109 4260 -61
rect 4000 -167 4052 -161
rect 4104 -161 4260 -109
rect 2046 -597 2098 -470
rect 4104 -294 4156 -161
rect 4104 -480 4156 -470
rect 6162 -294 6214 124
rect 8220 300 8272 310
rect 8220 -9 8272 124
rect 8300 74 8352 80
rect 8300 16 8352 22
rect 8220 -71 8272 -61
rect 2046 -655 2098 -649
rect 6162 -597 6214 -470
rect 8220 -109 8272 -99
rect 8220 -294 8272 -161
rect 8303 -186 8349 16
rect 8300 -192 8352 -186
rect 8300 -250 8352 -244
rect 8220 -480 8272 -470
rect 6162 -655 6214 -649
use sky130_fd_pr__pfet_01v8_P4G5X4  sky130_fd_pr__pfet_01v8_P4G5X4_0
timestamp 1762752159
transform -1 0 -30 0 -1 212
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_P4G5X4  sky130_fd_pr__pfet_01v8_P4G5X4_1
timestamp 1762752159
transform -1 0 -30 0 -1 -382
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_P4G5X4  sky130_fd_pr__pfet_01v8_P4G5X4_2
timestamp 1762752159
transform -1 0 8290 0 -1 -382
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_P4G5X4  sky130_fd_pr__pfet_01v8_P4G5X4_3
timestamp 1762752159
transform -1 0 8290 0 -1 212
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_PDVD34  sky130_fd_pr__pfet_01v8_PDVD34_0
timestamp 1762752159
transform 1 0 4130 0 1 212
box -4181 -200 4181 200
use sky130_fd_pr__pfet_01v8_PDVD34  sky130_fd_pr__pfet_01v8_PDVD34_1
timestamp 1762752159
transform 1 0 4130 0 1 -382
box -4181 -200 4181 200
<< labels >>
rlabel polycont 8313 -546 8313 -546 0 G
port 2 nsew
rlabel polycont -53 -546 -53 -546 0 G
port 2 nsew
flabel metal2 6185 -580 6185 -580 0 FreeSans 160 0 0 0 vdde
port 3 nsew
flabel metal2 8329 -97 8329 -97 0 FreeSans 160 0 0 0 d10
port 1 nsew
flabel metal2 8254 9 8254 9 0 FreeSans 160 0 0 0 d1
port 0 nsew
flabel metal2 8244 -180 8244 -180 0 FreeSans 160 0 0 0 d2
port 4 nsew
<< end >>
