* PEX produced on Min 07 Jul 2024 12:20:57  WIB using ./iic-pex.sh with m=3 and s=1
* NGSPICE file created from bgr_op5_block_rev1.ext - technology: sky130A

.subckt bgr_op5_block_rev1 ENA AVDD DVDD VREF VBGSC TRIM3 TRIM2 IPTAT VENA DVSS TRIM0
+ TRIM1 AVSS VBGTC
X0 VREF.t12 VREF.t10 VREF.t11 digital_0.VDDE.t35 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
X1 pmos_current_bgr_2_0.D3.t15 pmos_current_bgr_2_0.D3.t13 pmos_current_bgr_2_0.D3.t14 AVSS.t117 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
X2 digital_0.S1.t41 TRIM0.t0 bjt_0.B.t29 DVSS.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X3 digital_0.D3.t13 TRIM3.t0 digital_0.S3.t3 DVSS.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X4 digital_0.S3.t21 digital_0.S3.t20 digital_0.S3.t21 DVSS.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.29 as=0 ps=0 w=4 l=0.15
X5 pmos_iptat_0.G.t21 resistor_op_tt_0.C.t16 digital_0.VDDE.t20 digital_0.VDDE.t19 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=10
X6 AVSS.t80 AVSS.t81 bjt_0.B.t27 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720 d=11121552,65696
X7 AVSS.t110 AVSS.t109 AVSS.t84 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720 d=11121552,65696
X8 pmos_startup_0.D3.t17 pmos_startup_0.D4.t3 AVSS.t19 AVSS.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X9 digital_0.VDDE.t3 pmos_current_bgr_2_0.D4.t4 pmos_current_bgr_2_0.D4.t5 digital_0.VDDE.t2 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=10
X10 a_n4883_22159.t1 a_n547_22325.t0 AVSS.t9 sky130_fd_pr__res_high_po_0p35 l=17
X11 a_n17355_21661.t0 a_n13555_21661.t1 AVSS.t17 sky130_fd_pr__res_high_po_0p35 l=17
X12 pmos_current_bgr_2_0.D4.t16 pmos_current_bgr_2_0.D4.t14 pmos_current_bgr_2_0.D4.t15 digital_0.VDDE.t13 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
X13 bjt_0.B.t28 TRIM0.t1 digital_0.S1.t40 DVSS.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X14 pmos_startup_0.D3.t11 pmos_startup_0.D3.t9 pmos_startup_0.D3.t10 AVSS.t2 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
X15 a_n13555_21329.t1 a_n9219_21163.t1 AVSS.t16 sky130_fd_pr__res_high_po_0p35 l=17
X16 a_n13555_20997.t1 a_n9219_20997.t1 AVSS.t16 sky130_fd_pr__res_high_po_0p35 l=17
X17 pmos_startup_0.D3.t8 pmos_startup_0.D3.t7 pmos_startup_0.D3.t8 AVSS.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.15
X18 a_n9219_19433.t1 a_n4883_19433.t1 AVSS.t6 sky130_fd_pr__res_high_po_0p35 l=17
X19 pmos_current_bgr_2_0.D4.t0 pmos_current_bgr_2_0.D3.t17 resistor_op_tt_0.A.t2 AVSS.t117 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=20
X20 digital_0.S3.t8 digital_0.D3.t16 AVSS.t10 sky130_fd_pr__res_high_po_0p35 l=8.4
X21 pmos_startup_0.D3.t6 pmos_startup_0.D3.t5 pmos_startup_0.D3.t6 digital_0.VDDE.t5 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.15
X22 a_n4883_22325.t0 a_n547_22159.t0 AVSS.t9 sky130_fd_pr__res_high_po_0p35 l=17
X23 a_n17355_21495.t1 a_n13555_21495.t0 AVSS.t17 sky130_fd_pr__res_high_po_0p35 l=17
X24 a_n9219_20595.t0 a_n4883_20595.t1 AVSS.t6 sky130_fd_pr__res_high_po_0p35 l=17
X25 a_n4883_19931.t1 a_n547_19931.t1 AVSS.t9 sky130_fd_pr__res_high_po_0p35 l=17
X26 digital_0.S3.t10 digital_0.S2.t26 AVSS.t13 sky130_fd_pr__res_high_po_0p35 l=8.4
X27 pmos_iptat_0.G.t22 resistor_op_tt_0.D.t7 sky130_fd_pr__cap_mim_m3_1 l=17 w=17
X28 IPTAT.t9 IPTAT.t7 IPTAT.t8 digital_0.VDDE.t8 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
X29 digital_0.VDDE.t61 digital_0.VDDE.t59 digital_0.VDDE.t60 DVDD.t0 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0 ps=0 w=2 l=0.15
X30 digital_0.VDDE.t58 digital_0.VDDE.t57 digital_0.VDDE.t58 digital_0.VDDE.t21 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=10
X31 AVSS.t121 pmos_current_bgr_2_0.D3.t18 pmos_iptat_0.G.t1 AVSS.t15 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=20
X32 a_n547_22159.t1 a_3789_22325.t0 AVSS.t23 sky130_fd_pr__res_high_po_0p35 l=17
X33 VREF.t9 VREF.t8 VREF.t9 digital_0.VDDE.t4 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.15
X34 bjt_0.B.t35 bjt_0.B.t36 AVSS.t10 sky130_fd_pr__res_high_po_0p35 l=8.4
X35 pmos_current_bgr_0.D1.t4 pmos_iptat_0.G.t23 digital_0.VDDE.t67 digital_0.VDDE.t45 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=10
X36 a_n9219_21827.t1 digital_0.SVBGSC.t1 AVSS.t6 sky130_fd_pr__res_high_po_0p35 l=17
X37 a_n4883_19765.t1 a_n547_19765.t1 AVSS.t9 sky130_fd_pr__res_high_po_0p35 l=17
X38 digital_0.S1.t57 bjt_0.B.t40 AVSS.t13 sky130_fd_pr__res_high_po_0p35 l=8.4
X39 bjt_0.B.t38 bjt_0.B.t39 AVSS.t10 sky130_fd_pr__res_high_po_0p35 l=8.4
X40 differential_pair_0.S.t11 differential_pair_0.S.t9 differential_pair_0.S.t10 AVSS.t47 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
X41 AVSS.t73 AVSS.t74 sky130_fd_pr__cap_mim_m3_1 l=17 w=17
X42 a_n4883_20429.t1 a_n547_20429.t1 AVSS.t9 sky130_fd_pr__res_high_po_0p35 l=17
X43 AVSS.t71 AVSS.t72 sky130_fd_pr__cap_mim_m3_1 l=17 w=17
X44 digital_0.VDDE.t56 digital_0.VDDE.t55 digital_0.VDDE.t56 digital_0.VDDE.t16 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=10
X45 a_3789_22159.t0 a_8125_21993.t0 AVSS.t23 sky130_fd_pr__res_high_po_0p35 l=17
X46 a_n9219_21163.t0 a_n4883_21329.t1 AVSS.t6 sky130_fd_pr__res_high_po_0p35 l=17
X47 AVSS.t80 AVSS.t79 bjt_0.B.t26 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720 d=11121552,65696
X48 a_n547_22325.t1 a_3789_22159.t1 AVSS.t34 sky130_fd_pr__res_high_po_0p35 l=17
X49 a_n547_19931.t0 a_3789_19931.t1 AVSS.t33 sky130_fd_pr__res_high_po_0p35 l=17
X50 resistor_op_tt_0.C.t15 differential_pair_0.D4.t16 digital_0.VDDE.t70 digital_0.VDDE.t0 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=10
X51 digital_0.S1.t53 digital_0.S1.t52 digital_0.S1.t53 DVSS.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.29 as=0 ps=0 w=4 l=0.15
X52 AVSS.t108 AVSS.t107 AVSS.t84 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720 d=11121552,65696
X53 pmos_current_bgr_2_0.D4.t13 pmos_current_bgr_2_0.D4.t11 pmos_current_bgr_2_0.D4.t12 AVSS.t117 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
X54 a_n4883_19599.t1 a_n547_19599.t0 AVSS.t9 sky130_fd_pr__res_high_po_0p35 l=17
X55 digital_0.S1.t14 digital_0.S1.t15 AVSS.t10 sky130_fd_pr__res_high_po_0p35 l=8.4
X56 pmos_startup_0.D3.t16 pmos_startup_0.D4.t4 AVSS.t1 AVSS.t0 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X57 AVSS.t90 AVSS.t105 AVSS.t106 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720 d=11121552,65696
X58 a_n4883_21661.t1 digital_0.D3.t15 AVSS.t9 sky130_fd_pr__res_high_po_0p35 l=17
X59 digital_0.S1.t12 digital_0.S1.t13 AVSS.t10 sky130_fd_pr__res_high_po_0p35 l=8.4
X60 pmos_iptat_0.G.t17 pmos_iptat_0.G.t15 pmos_iptat_0.G.t16 digital_0.VDDE.t35 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
X61 digital_0.S2.t22 digital_0.S2.t20 digital_0.S2.t21 DVSS.t0 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=0 ps=0 w=4 l=0.15
X62 a_n4883_22491.t0 a_n547_22491.t0 AVSS.t9 sky130_fd_pr__res_high_po_0p35 l=17
X63 a_3789_22325.t1 a_8125_21827.t0 AVSS.t34 sky130_fd_pr__res_high_po_0p35 l=17
X64 a_3789_19931.t0 a_8125_19931.t0 AVSS.t33 sky130_fd_pr__res_high_po_0p35 l=17
X65 pmos_startup_0.D3.t4 pmos_startup_0.D3.t2 pmos_startup_0.D3.t3 AVSS.t0 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
X66 AVSS.t69 AVSS.t70 sky130_fd_pr__cap_mim_m3_1 l=17 w=17
X67 digital_0.S3.t2 TRIM3.t1 digital_0.D3.t12 DVSS.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X68 digital_0.D3.t9 digital_0.D3.t7 digital_0.D3.t8 DVSS.t3 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=0 ps=0 w=4 l=0.15
X69 differential_pair_0.D4.t15 differential_pair_0.D4.t13 differential_pair_0.D4.t14 AVSS.t28 sky130_fd_pr__nfet_01v8 ad=0.261 pd=2.38 as=0 ps=0 w=0.9 l=0.15
X70 VREF.t13 pmos_iptat_0.G.t24 digital_0.VDDE.t65 digital_0.VDDE.t19 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=10
X71 pmos_iptat_0.G.t0 pmos_current_bgr_2_0.D3.t19 AVSS.t120 AVSS.t47 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=20
X72 digital_0.SVBGSC.t0 VENA.t0 VBGSC.t7 DVSS.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X73 VBGTC.t5 VBGTC.t3 VBGTC.t4 DVSS.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
X74 a_n547_19765.t0 a_3789_19765.t0 AVSS.t32 sky130_fd_pr__res_high_po_0p35 l=17
X75 digital_0.VDDE.t34 pmos_iptat_0.G.t25 VREF.t1 digital_0.VDDE.t32 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=10
X76 digital_0.S2.t5 TRIM2.t0 digital_0.S3.t5 DVSS.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X77 pmos_startup_0.D3.t1 pmos_startup_0.D3.t0 pmos_startup_0.D3.t1 AVSS.t0 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.15
X78 AVSS.t90 AVSS.t103 AVSS.t104 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720 d=11121552,65696
X79 differential_pair_0.PLUS.t1 a_n13555_21163.t1 AVSS.t17 sky130_fd_pr__res_high_po_0p35 l=17
X80 a_n547_20429.t0 a_3789_20429.t0 AVSS.t14 sky130_fd_pr__res_high_po_0p35 l=17
X81 digital_0.S2.t0 digital_0.S1.t0 AVSS.t13 sky130_fd_pr__res_high_po_0p35 l=8.4
X82 AVSS.t67 AVSS.t68 sky130_fd_pr__cap_mim_m3_1 l=17 w=17
X83 AVSS.t129 a_n13555_20997.t0 AVSS.t17 sky130_fd_pr__res_high_po_0p35 l=17
X84 a_n9219_20263.t0 a_n4883_20263.t1 AVSS.t6 sky130_fd_pr__res_high_po_0p35 l=17
X85 digital_0.S1.t37 bjt_0.B.t19 AVSS.t10 sky130_fd_pr__res_high_po_0p35 l=8.4
X86 AVSS.t80 AVSS.t114 bjt_0.B.t25 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720 d=11121552,65696
X87 a_3789_19765.t1 a_8125_19599.t1 AVSS.t32 sky130_fd_pr__res_high_po_0p35 l=17
X88 digital_0.VDDE.t9 differential_pair_0.D4.t4 differential_pair_0.D4.t5 digital_0.VDDE.t2 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=10
X89 digital_0.VDDE.t72 ENA.t0 AVDD.t3 DVDD.t1 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X90 a_3789_20429.t1 a_8125_20263.t1 AVSS.t14 sky130_fd_pr__res_high_po_0p35 l=17
X91 differential_pair_0.D4.t12 differential_pair_0.D4.t10 differential_pair_0.D4.t11 digital_0.VDDE.t13 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
X92 AVDD.t2 ENA.t1 digital_0.VDDE.t11 DVDD.t1 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X93 digital_0.VDDE.t54 digital_0.VDDE.t52 digital_0.VDDE.t53 DVDD.t1 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.15
X94 digital_0.S1.t51 digital_0.S1.t49 digital_0.S1.t50 DVSS.t3 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=0 ps=0 w=4 l=0.15
X95 digital_0.S2.t12 TRIM1.t0 digital_0.S1.t31 DVSS.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X96 differential_pair_0.D4.t1 bjt_0.A.t2 differential_pair_0.S.t3 AVSS.t27 sky130_fd_pr__nfet_01v8 ad=0.1305 pd=1.19 as=0.1305 ps=1.19 w=0.9 l=13
X97 a_n547_19599.t1 a_3789_19599.t1 AVSS.t39 sky130_fd_pr__res_high_po_0p35 l=17
X98 AVSS.t3 pmos_startup_0.D4.t5 pmos_startup_0.D3.t15 AVSS.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X99 digital_0.D3.t6 digital_0.D3.t5 digital_0.D3.t6 DVSS.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.29 as=0 ps=0 w=4 l=0.15
X100 a_n547_21993.t1 a_3789_21827.t0 AVSS.t42 sky130_fd_pr__res_high_po_0p35 l=17
X101 resistor_op_tt_0.C.t14 resistor_op_tt_0.C.t13 resistor_op_tt_0.C.t14 AVSS.t28 sky130_fd_pr__nfet_01v8 ad=0.1305 pd=1.19 as=0 ps=0 w=0.9 l=0.15
X102 a_n13555_22159.t1 a_n9219_22325.t1 AVSS.t16 sky130_fd_pr__res_high_po_0p35 l=17
X103 differential_pair_0.PLUS.t0 a_n4883_21661.t0 AVSS.t6 sky130_fd_pr__res_high_po_0p35 l=17
X104 digital_0.S1.t32 bjt_0.B.t17 AVSS.t13 sky130_fd_pr__res_high_po_0p35 l=8.4
X105 a_n547_22491.t1 a_3789_22491.t0 AVSS.t35 sky130_fd_pr__res_high_po_0p35 l=17
X106 a_n9219_20097.t1 a_n4883_20097.t0 AVSS.t6 sky130_fd_pr__res_high_po_0p35 l=17
X107 a_n4883_19433.t0 a_n547_19433.t0 AVSS.t9 sky130_fd_pr__res_high_po_0p35 l=17
X108 digital_0.S2.t24 digital_0.S2.t25 AVSS.t13 sky130_fd_pr__res_high_po_0p35 l=8.4
X109 digital_0.VDDE.t23 pmos_iptat_0.G.t26 pmos_current_bgr_0.D1.t3 digital_0.VDDE.t21 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=10
X110 pmos_current_bgr_2_0.D4.t10 pmos_current_bgr_2_0.D4.t9 pmos_current_bgr_2_0.D4.t10 digital_0.VDDE.t25 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.15
X111 pmos_iptat_0.G.t27 resistor_op_tt_0.D.t6 sky130_fd_pr__cap_mim_m3_1 l=17 w=17
X112 digital_0.S1.t6 TRIM1.t1 digital_0.S2.t2 DVSS.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X113 a_3789_19599.t0 a_8125_19599.t0 AVSS.t39 sky130_fd_pr__res_high_po_0p35 l=17
X114 resistor_op_tt_0.A.t1 pmos_current_bgr_2_0.D3.t20 pmos_current_bgr_2_0.D4.t1 AVSS.t5 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=20
X115 digital_0.SVBGTC.t3 a_8125_21827.t1 AVSS.t42 sky130_fd_pr__res_high_po_0p35 l=17
X116 a_n4883_20595.t0 a_n547_20595.t0 AVSS.t9 sky130_fd_pr__res_high_po_0p35 l=17
X117 pmos_iptat_0.G.t14 pmos_iptat_0.G.t12 pmos_iptat_0.G.t13 AVSS.t47 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
X118 digital_0.VDDE.t31 pmos_iptat_0.G.t28 IPTAT.t13 digital_0.VDDE.t29 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=10
X119 digital_0.S2.t19 digital_0.S2.t18 digital_0.S2.t19 DVSS.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.29 as=0 ps=0 w=4 l=0.15
X120 AVSS.t102 AVSS.t101 AVSS.t84 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720 d=11121552,65696
X121 a_3789_22491.t1 AVSS.t125 AVSS.t35 sky130_fd_pr__res_high_po_0p35 l=17
X122 digital_0.VDDE.t51 digital_0.VDDE.t50 digital_0.VDDE.t51 digital_0.VDDE.t45 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=10
X123 a_n13555_22325.t1 a_n9219_22159.t1 AVSS.t16 sky130_fd_pr__res_high_po_0p35 l=17
X124 a_n9219_21661.t0 a_n4883_21495.t0 AVSS.t6 sky130_fd_pr__res_high_po_0p35 l=17
X125 a_n13019_19765.t1 a_n9219_19931.t1 AVSS.t16 sky130_fd_pr__res_high_po_0p35 l=17
X126 digital_0.S1.t27 digital_0.S1.t28 AVSS.t10 sky130_fd_pr__res_high_po_0p35 l=8.4
X127 bjt_0.B.t37 digital_0.S1.t56 AVSS.t10 sky130_fd_pr__res_high_po_0p35 l=8.4
X128 digital_0.S2.t7 digital_0.S1.t9 AVSS.t10 sky130_fd_pr__res_high_po_0p35 l=8.4
X129 differential_pair_0.D4.t9 differential_pair_0.D4.t8 differential_pair_0.D4.t9 digital_0.VDDE.t25 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.15
X130 AVSS.t76 AVSS.t100 AVSS.t76 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720 d=11121552,65696
X131 pmos_startup_0.D4.t1 pmos_startup_0.D4.t0 pmos_startup_0.D4.t1 digital_0.VDDE.t5 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.15
X132 pmos_iptat_0.G.t11 pmos_iptat_0.G.t9 pmos_iptat_0.G.t10 digital_0.VDDE.t35 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
X133 a_n9219_21993.t1 a_n547_21993.t0 AVSS.t9 sky130_fd_pr__res_high_po_0p35 l=17
X134 differential_pair_0.S.t0 differential_pair_0.PLUS.t2 resistor_op_tt_0.C.t1 AVSS.t27 sky130_fd_pr__nfet_01v8 ad=0.1305 pd=1.19 as=0.1305 ps=1.19 w=0.9 l=13
X135 a_n547_19433.t1 a_3789_19433.t0 AVSS.t46 sky130_fd_pr__res_high_po_0p35 l=17
X136 IPTAT.t6 IPTAT.t5 IPTAT.t6 digital_0.VDDE.t18 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.15
X137 AVSS.t65 AVSS.t66 sky130_fd_pr__cap_mim_m3_1 l=17 w=17
X138 a_n13019_19765.t0 a_n9219_19765.t1 AVSS.t16 sky130_fd_pr__res_high_po_0p35 l=17
X139 AVDD.t1 ENA.t2 digital_0.VDDE.t62 DVDD.t0 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X140 digital_0.VDDE.t6 ENA.t3 AVDD.t0 DVDD.t0 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X141 AVSS.t90 AVSS.t98 AVSS.t99 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720 d=11121552,65696
X142 AVSS.t76 AVSS.t97 AVSS.t76 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720 d=11121552,65696
X143 AVSS.t41 a_n9219_20429.t1 AVSS.t16 sky130_fd_pr__res_high_po_0p35 l=17
X144 digital_0.S1.t26 digital_0.S2.t9 AVSS.t10 sky130_fd_pr__res_high_po_0p35 l=8.4
X145 digital_0.S1.t11 bjt_0.B.t6 AVSS.t10 sky130_fd_pr__res_high_po_0p35 l=8.4
X146 pmos_iptat_0.G.t8 pmos_iptat_0.G.t6 pmos_iptat_0.G.t7 AVSS.t15 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
X147 digital_0.VDDE.t49 digital_0.VDDE.t47 digital_0.VDDE.t48 DVDD.t0 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.15
X148 pmos_startup_0.D3.t13 pmos_startup_0.D3.t12 digital_0.VDDE.t68 digital_0.VDDE.t14 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=10
X149 a_n4883_21163.t0 a_n547_21329.t0 AVSS.t9 sky130_fd_pr__res_high_po_0p35 l=17
X150 a_n547_20595.t1 a_3789_20595.t1 AVSS.t44 sky130_fd_pr__res_high_po_0p35 l=17
X151 IPTAT.t12 pmos_iptat_0.G.t29 digital_0.VDDE.t28 digital_0.VDDE.t26 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=10
X152 AVSS.t78 AVSS.t96 AVSS.t78 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720 d=11121552,65696
X153 AVSS.t95 AVSS.t94 AVSS.t84 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720 d=11121552,65696
X154 a_3789_19433.t1 AVSS.t122 AVSS.t46 sky130_fd_pr__res_high_po_0p35 l=17
X155 digital_0.S3.t6 TRIM2.t1 digital_0.S2.t6 DVSS.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X156 digital_0.VDDE.t63 resistor_op_tt_0.C.t17 pmos_iptat_0.G.t20 digital_0.VDDE.t32 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=10
X157 resistor_op_tt_0.D.t1 resistor_op_tt_0.D.t2 sky130_fd_pr__cap_mim_m3_1 l=17 w=17
X158 a_3789_20595.t0 AVSS.t45 AVSS.t44 sky130_fd_pr__res_high_po_0p35 l=17
X159 pmos_startup_0.D2.t1 a_n9219_19599.t1 AVSS.t16 sky130_fd_pr__res_high_po_0p35 l=17
X160 AVSS.t4 pmos_startup_0.D4.t6 pmos_startup_0.D3.t14 AVSS.t0 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X161 a_n13555_21993.t0 a_n9219_21827.t0 AVSS.t16 sky130_fd_pr__res_high_po_0p35 l=17
X162 AVSS.t78 AVSS.t93 AVSS.t78 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720 d=11121552,65696
X163 digital_0.SVBGSC.t2 digital_0.SVBGTC.t2 AVSS.t38 sky130_fd_pr__res_high_po_0p35 l=17
X164 digital_0.S1.t42 digital_0.S1.t43 AVSS.t10 sky130_fd_pr__res_high_po_0p35 l=8.4
X165 digital_0.S1.t23 digital_0.S1.t24 AVSS.t10 sky130_fd_pr__res_high_po_0p35 l=8.4
X166 digital_0.S3.t19 digital_0.S3.t17 digital_0.S3.t18 DVSS.t0 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=0 ps=0 w=4 l=0.15
X167 a_n13555_22491.t1 a_n9219_22491.t1 AVSS.t16 sky130_fd_pr__res_high_po_0p35 l=17
X168 pmos_current_bgr_2_0.D3.t12 pmos_current_bgr_2_0.D3.t11 pmos_current_bgr_2_0.D3.t12 digital_0.VDDE.t25 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.15
X169 differential_pair_0.S.t5 pmos_current_bgr_2_0.D3.t21 AVSS.t119 AVSS.t15 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=20
X170 VREF.t0 a_n13555_22325.t0 AVSS.t17 sky130_fd_pr__res_high_po_0p35 l=17
X171 a_n4883_20263.t0 a_n547_20263.t0 AVSS.t9 sky130_fd_pr__res_high_po_0p35 l=17
X172 VREF.t7 VREF.t6 VREF.t7 digital_0.VDDE.t4 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.15
X173 AVSS.t63 AVSS.t64 sky130_fd_pr__cap_mim_m3_1 l=17 w=17
X174 a_3789_21827.t1 a_8125_21993.t1 AVSS.t38 sky130_fd_pr__res_high_po_0p35 l=17
X175 a_n547_21163.t1 a_3789_21329.t0 AVSS.t50 sky130_fd_pr__res_high_po_0p35 l=17
X176 pmos_iptat_0.G.t27 resistor_op_tt_0.D.t5 sky130_fd_pr__cap_mim_m3_1 l=17 w=17
X177 VBGSC.t5 VBGSC.t3 VBGSC.t4 DVSS.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
X178 a_n9219_21329.t1 a_n4883_21163.t1 AVSS.t6 sky130_fd_pr__res_high_po_0p35 l=17
X179 a_n9219_20997.t0 a_n4883_20997.t0 AVSS.t6 sky130_fd_pr__res_high_po_0p35 l=17
X180 bjt_0.B.t15 digital_0.S1.t25 AVSS.t10 sky130_fd_pr__res_high_po_0p35 l=8.4
X181 digital_0.S2.t28 digital_0.S1.t55 AVSS.t10 sky130_fd_pr__res_high_po_0p35 l=8.4
X182 digital_0.VDDE.t46 digital_0.VDDE.t44 digital_0.VDDE.t46 digital_0.VDDE.t45 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=10
X183 digital_0.S1.t17 bjt_0.B.t8 AVSS.t10 sky130_fd_pr__res_high_po_0p35 l=8.4
X184 AVSS.t124 a_220_15663.t1 AVSS.t123 sky130_fd_pr__res_high_po_0p35 l=4.5
X185 a_n4883_21495.t2 a_n4883_21495.t3 AVSS.t9 sky130_fd_pr__res_high_po_0p35 l=17
X186 a_3789_21163.t0 a_8125_21329.t1 AVSS.t50 sky130_fd_pr__res_high_po_0p35 l=17
X187 VBGTC.t7 VENA.t1 digital_0.SVBGTC.t1 DVSS.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X188 pmos_current_bgr_0.D1.t0 a_n13555_22159.t0 AVSS.t17 sky130_fd_pr__res_high_po_0p35 l=17
X189 a_n4883_20097.t1 a_n547_20097.t1 AVSS.t9 sky130_fd_pr__res_high_po_0p35 l=17
X190 digital_0.S1.t4 digital_0.S1.t5 AVSS.t10 sky130_fd_pr__res_high_po_0p35 l=8.4
X191 bjt_0.B.t16 digital_0.S1.t29 AVSS.t10 sky130_fd_pr__res_high_po_0p35 l=8.4
X192 digital_0.S2.t17 digital_0.S2.t15 digital_0.S2.t16 DVSS.t3 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=0 ps=0 w=4 l=0.15
X193 AVSS.t90 AVSS.t91 AVSS.t92 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720 d=11121552,65696
X194 AVSS.t29 a_n9219_19433.t0 AVSS.t16 sky130_fd_pr__res_high_po_0p35 l=17
X195 digital_0.S1.t59 digital_0.S2.t31 AVSS.t10 sky130_fd_pr__res_high_po_0p35 l=8.4
X196 digital_0.S1.t10 bjt_0.B.t5 AVSS.t10 sky130_fd_pr__res_high_po_0p35 l=8.4
X197 AVSS.t61 AVSS.t62 sky130_fd_pr__cap_mim_m3_1 l=17 w=17
X198 AVSS.t76 AVSS.t113 bjt_0.B.t24 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720 d=11121552,65696
X199 bjt_0.B.t32 bjt_0.B.t33 AVSS.t10 sky130_fd_pr__res_high_po_0p35 l=8.4
X200 resistor_op_tt_0.D.t0 a_220_14999.t1 AVSS.t37 sky130_fd_pr__res_high_po_0p35 l=4.5
X201 a_n547_20263.t1 a_3789_20263.t1 AVSS.t12 sky130_fd_pr__res_high_po_0p35 l=17
X202 VREF.t5 VREF.t3 VREF.t4 digital_0.VDDE.t35 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
X203 VREF.t14 pmos_iptat_0.G.t24 digital_0.VDDE.t64 digital_0.VDDE.t19 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=10
X204 a_n9219_21495.t1 a_n547_21495.t0 AVSS.t9 sky130_fd_pr__res_high_po_0p35 l=17
X205 AVSS.t43 a_n9219_20595.t1 AVSS.t16 sky130_fd_pr__res_high_po_0p35 l=17
X206 digital_0.S2.t27 TRIM2.t2 digital_0.S3.t11 DVSS.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X207 pmos_startup_0.D2.t4 pmos_startup_0.D2.t2 pmos_startup_0.D2.t3 digital_0.VDDE.t12 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
X208 differential_pair_0.S.t8 differential_pair_0.S.t6 differential_pair_0.S.t7 AVSS.t15 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
X209 digital_0.D3.t11 TRIM3.t2 digital_0.S3.t0 DVSS.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X210 IPTAT.t4 IPTAT.t2 IPTAT.t3 digital_0.VDDE.t8 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
X211 digital_0.S2.t30 digital_0.S3.t23 AVSS.t10 sky130_fd_pr__res_high_po_0p35 l=8.4
X212 digital_0.S1.t39 TRIM0.t2 bjt_0.B.t31 DVSS.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X213 digital_0.VDDE.t69 resistor_op_tt_0.C.t18 pmos_iptat_0.G.t19 digital_0.VDDE.t32 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=10
X214 pmos_current_bgr_2_0.D4.t8 pmos_current_bgr_2_0.D4.t6 pmos_current_bgr_2_0.D4.t7 AVSS.t5 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
X215 digital_0.S3.t16 digital_0.S3.t15 digital_0.S3.t16 DVSS.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.29 as=0 ps=0 w=4 l=0.15
X216 a_220_15663.t0 AVSS.t31 AVSS.t30 sky130_fd_pr__res_high_po_0p35 l=4.5
X217 a_3789_20263.t0 a_8125_20263.t0 AVSS.t12 sky130_fd_pr__res_high_po_0p35 l=17
X218 resistor_op_tt_0.C.t12 resistor_op_tt_0.C.t10 resistor_op_tt_0.C.t11 AVSS.t27 sky130_fd_pr__nfet_01v8 ad=0.261 pd=2.38 as=0 ps=0 w=0.9 l=0.15
X219 a_n547_21495.t1 a_3789_21661.t0 AVSS.t11 sky130_fd_pr__res_high_po_0p35 l=17
X220 AVSS.t59 AVSS.t60 sky130_fd_pr__cap_mim_m3_1 l=17 w=17
X221 AVSS.t57 AVSS.t58 sky130_fd_pr__cap_mim_m3_1 l=17 w=17
X222 AVSS.t78 AVSS.t77 bjt_0.B.t23 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720 d=11121552,65696
X223 a_n547_20097.t0 a_3789_20097.t0 AVSS.t36 sky130_fd_pr__res_high_po_0p35 l=17
X224 digital_0.S2.t23 digital_0.S1.t36 AVSS.t10 sky130_fd_pr__res_high_po_0p35 l=8.4
X225 a_n13555_21827.t0 a_n9219_21993.t0 AVSS.t16 sky130_fd_pr__res_high_po_0p35 l=17
X226 bjt_0.B.t30 TRIM0.t3 digital_0.S1.t38 DVSS.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X227 AVSS.t90 AVSS.t88 AVSS.t89 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720 d=11121552,65696
X228 VBGSC.t2 VBGSC.t0 VBGSC.t1 DVSS.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.15
X229 VBGTC.t2 VBGTC.t0 VBGTC.t1 DVSS.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.15
X230 a_n17355_21661.t1 a_n13555_21827.t1 AVSS.t17 sky130_fd_pr__res_high_po_0p35 l=17
X231 AVSS.t18 a_n13555_22491.t0 AVSS.t17 sky130_fd_pr__res_high_po_0p35 l=17
X232 a_3789_21495.t0 a_8125_21329.t0 AVSS.t11 sky130_fd_pr__res_high_po_0p35 l=17
X233 AVSS.t118 pmos_current_bgr_2_0.D3.t3 pmos_current_bgr_2_0.D3.t4 AVSS.t117 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=20
X234 a_220_15165.t3 resistor_op_tt_0.A.t3 AVSS.t130 sky130_fd_pr__res_high_po_0p35 l=4.5
X235 a_n13555_21163.t0 a_n9219_21329.t0 AVSS.t16 sky130_fd_pr__res_high_po_0p35 l=17
X236 a_3789_20097.t1 a_8125_19931.t1 AVSS.t36 sky130_fd_pr__res_high_po_0p35 l=17
X237 digital_0.SVBGTC.t0 VENA.t2 VBGTC.t6 DVSS.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X238 a_n4883_21495.t1 a_3789_21495.t1 AVSS.t40 sky130_fd_pr__res_high_po_0p35 l=17
X239 bjt_0.B.t34 digital_0.S1.t54 AVSS.t10 sky130_fd_pr__res_high_po_0p35 l=8.4
X240 digital_0.VDDE.t22 pmos_iptat_0.G.t26 pmos_current_bgr_0.D1.t2 digital_0.VDDE.t21 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=10
X241 pmos_current_bgr_2_0.D3.t2 pmos_current_bgr_2_0.D3.t1 AVSS.t116 AVSS.t5 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=20
X242 AVSS.t52 a_220_15165.t2 AVSS.t51 sky130_fd_pr__res_high_po_0p35 l=4.5
X243 digital_0.S1.t16 bjt_0.B.t7 AVSS.t10 sky130_fd_pr__res_high_po_0p35 l=8.4
X244 digital_0.S2.t14 digital_0.S2.t13 digital_0.S2.t14 DVSS.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.29 as=0 ps=0 w=4 l=0.15
X245 differential_pair_0.D4.t7 differential_pair_0.D4.t6 differential_pair_0.D4.t7 AVSS.t27 sky130_fd_pr__nfet_01v8 ad=0.1305 pd=1.19 as=0 ps=0 w=0.9 l=0.15
X246 pmos_startup_0.D4.t2 pmos_startup_0.D2.t5 digital_0.VDDE.t15 digital_0.VDDE.t14 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=10
X247 pmos_iptat_0.G.t5 pmos_iptat_0.G.t4 pmos_iptat_0.G.t5 digital_0.VDDE.t4 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.15
X248 bjt_0.B.t4 digital_0.S1.t8 AVSS.t10 sky130_fd_pr__res_high_po_0p35 l=8.4
X249 a_3789_21661.t1 a_8125_21163.t1 AVSS.t40 sky130_fd_pr__res_high_po_0p35 l=17
X250 digital_0.S1.t34 digital_0.S1.t35 AVSS.t10 sky130_fd_pr__res_high_po_0p35 l=8.4
X251 bjt_0.B.t3 digital_0.S1.t3 AVSS.t10 sky130_fd_pr__res_high_po_0p35 l=8.4
X252 pmos_current_bgr_0.D1.t1 pmos_iptat_0.G.t23 digital_0.VDDE.t66 digital_0.VDDE.t45 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=10
X253 resistor_op_tt_0.C.t9 resistor_op_tt_0.C.t8 resistor_op_tt_0.C.t9 digital_0.VDDE.t25 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.15
X254 AVSS.t76 AVSS.t75 bjt_0.B.t22 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720 d=11121552,65696
X255 bjt_0.B.t0 bjt_0.B.t1 AVSS.t10 sky130_fd_pr__res_high_po_0p35 l=8.4
X256 bjt_0.B.t13 bjt_0.B.t14 AVSS.t10 sky130_fd_pr__res_high_po_0p35 l=8.4
X257 pmos_current_bgr_2_0.D4.t3 pmos_current_bgr_2_0.D4.t2 digital_0.VDDE.t1 digital_0.VDDE.t0 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=10
X258 AVSS.t26 a_220_15165.t1 AVSS.t25 sky130_fd_pr__res_high_po_0p35 l=4.5
X259 resistor_op_tt_0.D.t3 a_220_14999.t3 AVSS.t128 sky130_fd_pr__res_high_po_0p35 l=4.5
X260 a_n9219_22159.t0 a_n4883_22325.t1 AVSS.t6 sky130_fd_pr__res_high_po_0p35 l=17
X261 a_n4883_21329.t0 a_n547_21163.t0 AVSS.t9 sky130_fd_pr__res_high_po_0p35 l=17
X262 a_n4883_20997.t1 a_n547_20997.t1 AVSS.t9 sky130_fd_pr__res_high_po_0p35 l=17
X263 a_n13019_20097.t1 a_n9219_20263.t1 AVSS.t16 sky130_fd_pr__res_high_po_0p35 l=17
X264 digital_0.S1.t7 digital_0.S2.t4 AVSS.t10 sky130_fd_pr__res_high_po_0p35 l=8.4
X265 AVSS.t80 AVSS.t87 AVSS.t80 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720 d=11121552,65696
X266 digital_0.S1.t20 digital_0.S2.t8 AVSS.t10 sky130_fd_pr__res_high_po_0p35 l=8.4
X267 a_220_14999.t0 resistor_op_tt_0.C.t0 AVSS.t24 sky130_fd_pr__res_high_po_0p35 l=4.5
X268 differential_pair_0.D4.t3 differential_pair_0.D4.t2 digital_0.VDDE.t7 digital_0.VDDE.t0 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=10
X269 digital_0.S1.t48 digital_0.S1.t47 digital_0.S1.t48 DVSS.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.29 as=0 ps=0 w=4 l=0.15
X270 AVSS.t78 AVSS.t112 bjt_0.B.t21 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720 d=11121552,65696
X271 digital_0.S3.t4 digital_0.S2.t3 AVSS.t10 sky130_fd_pr__res_high_po_0p35 l=8.4
X272 pmos_iptat_0.G.t18 resistor_op_tt_0.C.t19 digital_0.VDDE.t71 digital_0.VDDE.t19 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=10
X273 digital_0.S3.t9 TRIM2.t3 digital_0.S2.t11 DVSS.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X274 a_n13555_21495.t1 a_n9219_21661.t1 AVSS.t16 sky130_fd_pr__res_high_po_0p35 l=17
X275 pmos_current_bgr_2_0.D3.t10 pmos_current_bgr_2_0.D3.t8 pmos_current_bgr_2_0.D3.t9 AVSS.t5 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
X276 a_n9219_22325.t0 a_n4883_22159.t0 AVSS.t6 sky130_fd_pr__res_high_po_0p35 l=17
X277 a_n13019_20097.t0 a_n9219_20097.t0 AVSS.t16 sky130_fd_pr__res_high_po_0p35 l=17
X278 a_n9219_19931.t0 a_n4883_19931.t0 AVSS.t6 sky130_fd_pr__res_high_po_0p35 l=17
X279 AVSS.t80 AVSS.t86 AVSS.t80 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720 d=11121552,65696
X280 AVSS.t76 AVSS.t111 bjt_0.B.t20 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720 d=11121552,65696
X281 AVSS.t115 pmos_current_bgr_2_0.D3.t22 differential_pair_0.S.t4 AVSS.t47 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=20
X282 digital_0.VDDE.t33 pmos_iptat_0.G.t25 VREF.t2 digital_0.VDDE.t32 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=10
X283 pmos_current_bgr_2_0.D3.t7 pmos_current_bgr_2_0.D3.t5 pmos_current_bgr_2_0.D3.t6 digital_0.VDDE.t13 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
X284 digital_0.VDDE.t24 pmos_current_bgr_2_0.D4.t17 pmos_current_bgr_2_0.D3.t0 digital_0.VDDE.t2 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=10
X285 VBGSC.t6 VENA.t3 digital_0.SVBGSC.t3 DVSS.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X286 digital_0.S3.t1 TRIM3.t3 digital_0.D3.t10 DVSS.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X287 digital_0.D3.t4 digital_0.D3.t2 digital_0.D3.t3 DVSS.t0 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=0 ps=0 w=4 l=0.15
X288 a_220_14999.t2 resistor_op_tt_0.C.t4 AVSS.t127 sky130_fd_pr__res_high_po_0p35 l=4.5
X289 a_n17355_21495.t0 a_n13555_21993.t1 AVSS.t17 sky130_fd_pr__res_high_po_0p35 l=17
X290 digital_0.S3.t14 digital_0.S3.t12 digital_0.S3.t13 DVSS.t3 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=0 ps=0 w=4 l=0.15
X291 resistor_op_tt_0.C.t2 differential_pair_0.PLUS.t3 differential_pair_0.S.t1 AVSS.t28 sky130_fd_pr__nfet_01v8 ad=0.1305 pd=1.19 as=0.1305 ps=1.19 w=0.9 l=13
X292 a_220_15165.t0 resistor_op_tt_0.A.t0 AVSS.t22 sky130_fd_pr__res_high_po_0p35 l=4.5
X293 digital_0.VDDE.t17 pmos_startup_0.D3.t18 pmos_startup_0.D2.t0 digital_0.VDDE.t16 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=10
X294 digital_0.VDDE.t30 pmos_iptat_0.G.t28 IPTAT.t11 digital_0.VDDE.t29 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=10
X295 a_n547_21329.t1 a_3789_21163.t1 AVSS.t126 sky130_fd_pr__res_high_po_0p35 l=17
X296 a_n547_20997.t0 a_3789_20997.t1 AVSS.t7 sky130_fd_pr__res_high_po_0p35 l=17
X297 digital_0.S1.t2 bjt_0.B.t2 AVSS.t10 sky130_fd_pr__res_high_po_0p35 l=8.4
X298 AVSS.t21 a_220_14833.t0 AVSS.t20 sky130_fd_pr__res_high_po_0p35 l=4.5
X299 a_n13555_21661.t0 a_n9219_21495.t0 AVSS.t16 sky130_fd_pr__res_high_po_0p35 l=17
X300 bjt_0.B.t42 bjt_0.B.t43 AVSS.t10 sky130_fd_pr__res_high_po_0p35 l=8.4
X301 pmos_iptat_0.G.t22 resistor_op_tt_0.D.t4 sky130_fd_pr__cap_mim_m3_1 l=17 w=17
X302 a_n9219_19765.t0 a_n4883_19765.t0 AVSS.t6 sky130_fd_pr__res_high_po_0p35 l=17
X303 AVSS.t55 AVSS.t56 sky130_fd_pr__cap_mim_m3_1 l=17 w=17
X304 bjt_0.A.t0 a_n13555_21329.t0 AVSS.t17 sky130_fd_pr__res_high_po_0p35 l=17
X305 a_n9219_20429.t0 a_n4883_20429.t0 AVSS.t6 sky130_fd_pr__res_high_po_0p35 l=17
X306 resistor_op_tt_0.C.t7 resistor_op_tt_0.C.t5 resistor_op_tt_0.C.t6 digital_0.VDDE.t13 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
X307 digital_0.VDDE.t10 differential_pair_0.D4.t17 resistor_op_tt_0.C.t3 digital_0.VDDE.t2 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=10
X308 AVSS.t78 AVSS.t82 bjt_0.A.t1 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720 d=11121552,65696
X309 bjt_0.B.t18 digital_0.S1.t33 AVSS.t10 sky130_fd_pr__res_high_po_0p35 l=8.4
X310 pmos_iptat_0.G.t3 pmos_iptat_0.G.t2 pmos_iptat_0.G.t3 digital_0.VDDE.t4 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.15
X311 digital_0.S2.t10 TRIM1.t2 digital_0.S1.t30 DVSS.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X312 digital_0.VDDE.t43 digital_0.VDDE.t41 digital_0.VDDE.t42 digital_0.VDDE.t12 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.15
X313 a_3789_21329.t1 a_8125_21163.t0 AVSS.t126 sky130_fd_pr__res_high_po_0p35 l=17
X314 a_3789_20997.t0 AVSS.t8 AVSS.t7 sky130_fd_pr__res_high_po_0p35 l=17
X315 digital_0.S1.t21 digital_0.S1.t22 AVSS.t13 sky130_fd_pr__res_high_po_0p35 l=8.4
X316 digital_0.S1.t18 digital_0.S1.t19 AVSS.t13 sky130_fd_pr__res_high_po_0p35 l=8.4
X317 bjt_0.B.t41 digital_0.S1.t58 AVSS.t10 sky130_fd_pr__res_high_po_0p35 l=8.4
X318 IPTAT.t10 pmos_iptat_0.G.t29 digital_0.VDDE.t27 digital_0.VDDE.t26 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=10
X319 digital_0.S1.t46 digital_0.S1.t44 digital_0.S1.t45 DVSS.t0 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=0 ps=0 w=4 l=0.15
X320 digital_0.D3.t1 digital_0.D3.t0 digital_0.D3.t1 DVSS.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.29 as=0 ps=0 w=4 l=0.15
X321 digital_0.VDDE.t40 digital_0.VDDE.t39 digital_0.VDDE.t40 digital_0.VDDE.t21 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=10
X322 IPTAT.t1 IPTAT.t0 IPTAT.t1 digital_0.VDDE.t18 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.15
X323 pmos_current_bgr_2_0.D3.t16 pmos_current_bgr_2_0.D4.t18 digital_0.VDDE.t73 digital_0.VDDE.t0 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=10
X324 a_n9219_19599.t0 a_n4883_19599.t0 AVSS.t6 sky130_fd_pr__res_high_po_0p35 l=17
X325 a_n9219_21993.t2 a_n9219_21993.t3 AVSS.t6 sky130_fd_pr__res_high_po_0p35 l=17
X326 AVSS.t53 AVSS.t54 sky130_fd_pr__cap_mim_m3_1 l=17 w=17
X327 digital_0.S1.t1 TRIM1.t3 digital_0.S2.t1 DVSS.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X328 bjt_0.B.t11 bjt_0.B.t12 AVSS.t10 sky130_fd_pr__res_high_po_0p35 l=8.4
X329 bjt_0.B.t9 bjt_0.B.t10 AVSS.t10 sky130_fd_pr__res_high_po_0p35 l=8.4
X330 digital_0.VDDE.t38 digital_0.VDDE.t36 digital_0.VDDE.t37 DVDD.t1 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0 ps=0 w=2 l=0.15
X331 AVSS.t85 AVSS.t83 AVSS.t84 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720 d=11121552,65696
X332 a_n9219_22491.t0 a_n4883_22491.t1 AVSS.t6 sky130_fd_pr__res_high_po_0p35 l=17
X333 digital_0.D3.t14 digital_0.S3.t7 AVSS.t13 sky130_fd_pr__res_high_po_0p35 l=8.4
X334 digital_0.S2.t29 digital_0.S3.t22 AVSS.t10 sky130_fd_pr__res_high_po_0p35 l=8.4
X335 differential_pair_0.S.t2 bjt_0.A.t3 differential_pair_0.D4.t0 AVSS.t28 sky130_fd_pr__nfet_01v8 ad=0.1305 pd=1.19 as=0.1305 ps=1.19 w=0.9 l=13
X336 a_220_14833.t1 AVSS.t49 AVSS.t48 sky130_fd_pr__res_high_po_0p35 l=4.5
R0 VREF.n8 VREF.t3 341.837
R1 VREF.n8 VREF.t10 341.837
R2 VREF.n2 VREF.t8 341.837
R3 VREF.n2 VREF.t6 341.837
R4 VREF.n9 VREF.t12 228.784
R5 VREF.n3 VREF.t9 228.784
R6 VREF.n3 VREF.t7 228.784
R7 VREF.n7 VREF.t5 228.215
R8 VREF.n11 VREF.n4 200.219
R9 VREF.n12 VREF.n1 200.219
R10 VREF VREF.n0 200.071
R11 VREF.n7 VREF.n5 199.65
R12 VREF.n9 VREF.n8 161.3
R13 VREF.n3 VREF.n2 161.3
R14 VREF.n6 VREF.t0 42.5516
R15 VREF.n5 VREF.t2 28.5655
R16 VREF.n5 VREF.t4 28.5655
R17 VREF.n4 VREF.t1 28.5655
R18 VREF.n4 VREF.t11 28.5655
R19 VREF.t9 VREF.n0 28.5655
R20 VREF.n0 VREF.t13 28.5655
R21 VREF.t7 VREF.n1 28.5655
R22 VREF.n1 VREF.t14 28.5655
R23 VREF.n12 VREF.n11 22.2635
R24 VREF VREF.n6 4.99763
R25 VREF.n7 VREF 3.72328
R26 VREF.n6 VREF 0.320143
R27 VREF.n12 VREF.n3 0.212038
R28 VREF.n10 VREF.n7 0.202854
R29 VREF VREF.n12 0.147239
R30 VREF.n10 VREF.n9 0.0810264
R31 VREF.n11 VREF.n10 0.0810264
R32 digital_0.VDDE.n80 digital_0.VDDE.n43 18850.6
R33 digital_0.VDDE.n80 digital_0.VDDE.n44 18847.1
R34 digital_0.VDDE.n101 digital_0.VDDE.n43 18822.4
R35 digital_0.VDDE.n101 digital_0.VDDE.n44 18818.8
R36 digital_0.VDDE.n107 digital_0.VDDE.n106 11410.6
R37 digital_0.VDDE.n107 digital_0.VDDE.n14 11410.6
R38 digital_0.VDDE.n16 digital_0.VDDE.n14 11410.6
R39 digital_0.VDDE.n106 digital_0.VDDE.n16 11410.6
R40 digital_0.VDDE.n76 digital_0.VDDE.n72 9504.71
R41 digital_0.VDDE.n77 digital_0.VDDE.n76 9504.71
R42 digital_0.VDDE.n82 digital_0.VDDE.n72 9501.18
R43 digital_0.VDDE.n82 digital_0.VDDE.n77 9501.18
R44 digital_0.VDDE.n110 digital_0.VDDE.n29 9310.59
R45 digital_0.VDDE.n41 digital_0.VDDE.n29 9310.59
R46 digital_0.VDDE.n41 digital_0.VDDE.n28 9310.59
R47 digital_0.VDDE.n110 digital_0.VDDE.n28 9310.59
R48 digital_0.VDDE.n94 digital_0.VDDE.n47 2009.22
R49 digital_0.VDDE.n98 digital_0.VDDE.n47 2008.85
R50 digital_0.VDDE.n100 digital_0.VDDE.n45 2007.72
R51 digital_0.VDDE.n100 digital_0.VDDE.n99 2007.34
R52 digital_0.VDDE.n15 digital_0.VDDE.n13 1217.13
R53 digital_0.VDDE.n116 digital_0.VDDE.n13 1217.13
R54 digital_0.VDDE.n116 digital_0.VDDE.n115 1217.13
R55 digital_0.VDDE.n115 digital_0.VDDE.n15 1217.13
R56 digital_0.VDDE.n75 digital_0.VDDE.n70 1013.84
R57 digital_0.VDDE.n75 digital_0.VDDE.n71 1013.84
R58 digital_0.VDDE.n83 digital_0.VDDE.n70 1013.46
R59 digital_0.VDDE.n83 digital_0.VDDE.n71 1013.46
R60 digital_0.VDDE.n111 digital_0.VDDE.n26 993.13
R61 digital_0.VDDE.n111 digital_0.VDDE.n27 993.13
R62 digital_0.VDDE.n40 digital_0.VDDE.n26 993.13
R63 digital_0.VDDE.n40 digital_0.VDDE.n27 993.13
R64 digital_0.VDDE.t45 digital_0.VDDE.t32 640.596
R65 digital_0.VDDE.n121 digital_0.VDDE.t36 442.656
R66 digital_0.VDDE.n121 digital_0.VDDE.t59 442.656
R67 digital_0.VDDE.n120 digital_0.VDDE.t52 442.656
R68 digital_0.VDDE.n120 digital_0.VDDE.t47 442.656
R69 digital_0.VDDE.n36 digital_0.VDDE.t41 394.608
R70 digital_0.VDDE.t32 digital_0.VDDE.t35 333.995
R71 digital_0.VDDE.t26 digital_0.VDDE.t4 323.723
R72 digital_0.VDDE.t2 digital_0.VDDE.t12 323.411
R73 digital_0.VDDE.t29 digital_0.VDDE.n78 320.298
R74 digital_0.VDDE.n79 digital_0.VDDE.t21 320.298
R75 digital_0.VDDE.n78 digital_0.VDDE.t19 310.026
R76 digital_0.VDDE.n109 digital_0.VDDE.t0 309.716
R77 digital_0.VDDE.n108 digital_0.VDDE.t16 309.716
R78 digital_0.VDDE.n81 digital_0.VDDE.t45 267.382
R79 digital_0.VDDE.t25 digital_0.VDDE.t14 250.129
R80 digital_0.VDDE.n37 digital_0.VDDE.t43 223.565
R81 digital_0.VDDE.n33 digital_0.VDDE.n32 205.286
R82 digital_0.VDDE.n23 digital_0.VDDE.n22 201.9
R83 digital_0.VDDE.n21 digital_0.VDDE.n20 201.9
R84 digital_0.VDDE.n52 digital_0.VDDE.n51 201.9
R85 digital_0.VDDE.n50 digital_0.VDDE.n49 201.9
R86 digital_0.VDDE.n91 digital_0.VDDE.n90 201.9
R87 digital_0.VDDE.n89 digital_0.VDDE.n88 201.9
R88 digital_0.VDDE.n19 digital_0.VDDE.n18 199.65
R89 digital_0.VDDE.n24 digital_0.VDDE.n17 199.65
R90 digital_0.VDDE.n68 digital_0.VDDE.n67 199.65
R91 digital_0.VDDE.n69 digital_0.VDDE.n66 199.65
R92 digital_0.VDDE.n92 digital_0.VDDE.n58 199.65
R93 digital_0.VDDE.n57 digital_0.VDDE.n55 199.65
R94 digital_0.VDDE.n62 digital_0.VDDE.n61 199.65
R95 digital_0.VDDE.n56 digital_0.VDDE.n53 199.65
R96 digital_0.VDDE.n59 digital_0.VDDE.n48 199.65
R97 digital_0.VDDE.n87 digital_0.VDDE.n63 199.65
R98 digital_0.VDDE.n38 digital_0.VDDE.n35 199.65
R99 digital_0.VDDE.n34 digital_0.VDDE.n33 199.65
R100 digital_0.VDDE.n122 digital_0.VDDE.n121 161.3
R101 digital_0.VDDE.n5 digital_0.VDDE.n120 161.3
R102 digital_0.VDDE.n122 digital_0.VDDE.t38 114.451
R103 digital_0.VDDE.n122 digital_0.VDDE.t61 114.451
R104 digital_0.VDDE.n9 digital_0.VDDE.t53 113.644
R105 digital_0.VDDE.n11 digital_0.VDDE.t48 113.644
R106 digital_0.pmos_ena_0.VDDE digital_0.VDDE.n123 100.168
R107 digital_0.pmos_ena_0.VDDE digital_0.VDDE.n124 100.144
R108 digital_0.VDDE.n9 digital_0.VDDE.n8 99.3605
R109 digital_0.VDDE.n11 digital_0.VDDE.n10 99.3605
R110 digital_0.VDDE.n103 digital_0.VDDE.n102 82.4874
R111 digital_0.VDDE.t35 digital_0.VDDE.n80 77.1997
R112 digital_0.VDDE.n37 digital_0.VDDE.n36 61.7417
R113 digital_0.VDDE.t18 digital_0.VDDE.n42 49.8039
R114 digital_0.VDDE.n81 digital_0.VDDE.t8 49.4926
R115 digital_0.VDDE.n105 digital_0.VDDE.t5 45.6005
R116 digital_0.VDDE.t13 digital_0.VDDE.n104 34.2403
R117 digital_0.VDDE.n104 digital_0.VDDE.n103 33.6178
R118 digital_0.VDDE.n22 digital_0.VDDE.t7 28.5655
R119 digital_0.VDDE.n22 digital_0.VDDE.t10 28.5655
R120 digital_0.VDDE.n20 digital_0.VDDE.t70 28.5655
R121 digital_0.VDDE.n20 digital_0.VDDE.t9 28.5655
R122 digital_0.VDDE.n18 digital_0.VDDE.t1 28.5655
R123 digital_0.VDDE.n18 digital_0.VDDE.t24 28.5655
R124 digital_0.VDDE.n17 digital_0.VDDE.t73 28.5655
R125 digital_0.VDDE.n17 digital_0.VDDE.t3 28.5655
R126 digital_0.VDDE.n67 digital_0.VDDE.t27 28.5655
R127 digital_0.VDDE.n67 digital_0.VDDE.t31 28.5655
R128 digital_0.VDDE.n66 digital_0.VDDE.t28 28.5655
R129 digital_0.VDDE.n66 digital_0.VDDE.t30 28.5655
R130 digital_0.VDDE.n58 digital_0.VDDE.t20 28.5655
R131 digital_0.VDDE.n58 digital_0.VDDE.t58 28.5655
R132 digital_0.VDDE.t58 digital_0.VDDE.n57 28.5655
R133 digital_0.VDDE.n57 digital_0.VDDE.t46 28.5655
R134 digital_0.VDDE.t40 digital_0.VDDE.n62 28.5655
R135 digital_0.VDDE.n62 digital_0.VDDE.t51 28.5655
R136 digital_0.VDDE.t46 digital_0.VDDE.n56 28.5655
R137 digital_0.VDDE.n56 digital_0.VDDE.t69 28.5655
R138 digital_0.VDDE.n51 digital_0.VDDE.t66 28.5655
R139 digital_0.VDDE.n51 digital_0.VDDE.t33 28.5655
R140 digital_0.VDDE.n49 digital_0.VDDE.t67 28.5655
R141 digital_0.VDDE.n49 digital_0.VDDE.t34 28.5655
R142 digital_0.VDDE.t51 digital_0.VDDE.n59 28.5655
R143 digital_0.VDDE.n59 digital_0.VDDE.t63 28.5655
R144 digital_0.VDDE.n90 digital_0.VDDE.t65 28.5655
R145 digital_0.VDDE.n90 digital_0.VDDE.t23 28.5655
R146 digital_0.VDDE.n88 digital_0.VDDE.t64 28.5655
R147 digital_0.VDDE.n88 digital_0.VDDE.t22 28.5655
R148 digital_0.VDDE.n63 digital_0.VDDE.t71 28.5655
R149 digital_0.VDDE.n63 digital_0.VDDE.t40 28.5655
R150 digital_0.VDDE.n35 digital_0.VDDE.t56 28.5655
R151 digital_0.VDDE.n35 digital_0.VDDE.t42 28.5655
R152 digital_0.VDDE.n34 digital_0.VDDE.t15 28.5655
R153 digital_0.VDDE.t56 digital_0.VDDE.n34 28.5655
R154 digital_0.VDDE.n32 digital_0.VDDE.t68 28.5655
R155 digital_0.VDDE.n32 digital_0.VDDE.t17 28.5655
R156 digital_0.VDDE.n106 digital_0.VDDE.n105 19.7826
R157 digital_0.VDDE.n28 digital_0.VDDE.n26 16.8187
R158 digital_0.VDDE.n105 digital_0.VDDE.n28 16.8187
R159 digital_0.VDDE.n29 digital_0.VDDE.n27 16.8187
R160 digital_0.VDDE.n104 digital_0.VDDE.n29 16.8187
R161 digital_0.VDDE.n83 digital_0.VDDE.n82 15.4172
R162 digital_0.VDDE.n82 digital_0.VDDE.n81 15.4172
R163 digital_0.VDDE.n76 digital_0.VDDE.n75 15.4172
R164 digital_0.VDDE.n76 digital_0.VDDE.n42 15.4172
R165 digital_0.VDDE.n119 digital_0.VDDE.n11 15.3143
R166 digital_0.VDDE.n54 digital_0.VDDE.t44 14.3181
R167 digital_0.VDDE.n54 digital_0.VDDE.t57 14.3181
R168 digital_0.VDDE.n60 digital_0.VDDE.t50 14.3181
R169 digital_0.VDDE.n60 digital_0.VDDE.t39 14.3181
R170 digital_0.VDDE.n124 digital_0.VDDE.t11 14.283
R171 digital_0.VDDE.n124 digital_0.VDDE.t37 14.283
R172 digital_0.VDDE.n8 digital_0.VDDE.t54 14.283
R173 digital_0.VDDE.n8 digital_0.VDDE.t72 14.283
R174 digital_0.VDDE.n10 digital_0.VDDE.t49 14.283
R175 digital_0.VDDE.n10 digital_0.VDDE.t6 14.283
R176 digital_0.VDDE.n123 digital_0.VDDE.t62 14.283
R177 digital_0.VDDE.n123 digital_0.VDDE.t60 14.283
R178 digital_0.VDDE.n31 digital_0.VDDE.t55 11.5219
R179 digital_0.VDDE.t5 digital_0.VDDE.t25 10.7672
R180 digital_0.VDDE.n109 digital_0.VDDE.n108 10.5837
R181 digital_0.VDDE.t16 digital_0.VDDE.t2 10.5837
R182 digital_0.VDDE.t12 digital_0.VDDE.t13 10.5837
R183 digital_0.VDDE.t4 digital_0.VDDE.t18 10.2725
R184 digital_0.VDDE.t19 digital_0.VDDE.t26 10.2725
R185 digital_0.VDDE.t21 digital_0.VDDE.t29 10.2725
R186 digital_0.VDDE.n36 digital_0.VDDE.n30 9.47441
R187 digital_0.VDDE.n96 digital_0.VDDE.n95 8.90539
R188 digital_0.VDDE.n97 digital_0.VDDE.n96 8.90267
R189 digital_0.VDDE.n93 digital_0.VDDE.n46 8.88365
R190 digital_0.VDDE.n25 pmos_current_bgr_2_0.vdde 8.76952
R191 digital_0.VDDE.n117 pmos_current_bgr_2_0.vdde 8.76952
R192 digital_0.VDDE.n119 digital_0.VDDE.n1 8.95156
R193 digital_0.VDDE.n102 digital_0.VDDE.n42 7.78228
R194 digital_0.VDDE.n74 pmos_iptat_0.VDDE 7.30213
R195 digital_0.VDDE.n84 pmos_iptat_0.VDDE 7.29941
R196 digital_0.VDDE.n23 digital_0.VDDE.n21 7.1617
R197 pmos_startup_0.VDDE digital_0.VDDE.n4 7.15267
R198 digital_0.VDDE.n112 digital_0.VDDE.n4 7.15267
R199 digital_0.VDDE.n106 digital_0.VDDE.n15 7.11588
R200 digital_0.VDDE.n116 digital_0.VDDE.n14 7.11588
R201 digital_0.VDDE.n103 digital_0.VDDE.n14 7.11588
R202 digital_0.VDDE.n80 digital_0.VDDE.n47 6.85235
R203 digital_0.VDDE.n101 digital_0.VDDE.n100 6.85235
R204 digital_0.VDDE.n102 digital_0.VDDE.n101 6.85235
R205 digital_0.VDDE.n114 pmos_current_bgr_2_0.VDDE 6.30485
R206 pmos_current_bgr_0.vdde digital_0.VDDE.n64 6.22061
R207 digital_0.VDDE.n73 digital_0.VDDE.n65 6.03782
R208 digital_0.VDDE.n7 digital_0.VDDE.n93 5.59289
R209 pmos_startup_0.VDDE digital_0.VDDE.n39 5.59289
R210 digital_0.VDDE.n6 digital_0.VDDE.n97 5.58202
R211 digital_0.VDDE.n95 digital_0.VDDE.n7 5.58202
R212 digital_0.VDDE.n69 digital_0.VDDE.n68 5.44762
R213 digital_0.VDDE.t14 digital_0.VDDE.t0 5.33758
R214 digital_0.VDDE.n38 digital_0.VDDE.n37 4.6505
R215 digital_0.VDDE.t8 digital_0.VDDE.n79 3.42448
R216 digital_0.VDDE.n53 digital_0.VDDE.n52 3.40194
R217 digital_0.VDDE.n50 digital_0.VDDE.n48 3.40194
R218 digital_0.VDDE.n92 digital_0.VDDE.n91 3.40194
R219 digital_0.VDDE.n89 digital_0.VDDE.n87 3.40194
R220 digital_0.VDDE.n24 digital_0.VDDE.n23 3.24863
R221 digital_0.VDDE.n21 digital_0.VDDE.n19 3.24667
R222 digital_0.VDDE.n33 digital_0.VDDE.n31 3.0935
R223 digital_0.VDDE.n86 digital_0.VDDE.n65 3.0005
R224 pmos_current_bgr_0.vdde digital_0.VDDE.n86 2.98963
R225 digital_0.VDDE.n31 digital_0.VDDE.n30 2.90811
R226 digital_0.VDDE.n3 digital_0.VDDE.n39 1.55683
R227 digital_0.VDDE.n77 digital_0.VDDE.n71 2.84665
R228 digital_0.VDDE.n78 digital_0.VDDE.n77 2.84665
R229 digital_0.VDDE.n72 digital_0.VDDE.n70 2.84665
R230 digital_0.VDDE.n78 digital_0.VDDE.n72 2.84665
R231 digital_0.VDDE.n111 digital_0.VDDE.n110 2.84665
R232 digital_0.VDDE.n110 digital_0.VDDE.n109 2.84665
R233 digital_0.VDDE.n41 digital_0.VDDE.n40 2.84665
R234 digital_0.VDDE.n109 digital_0.VDDE.n41 2.84665
R235 digital_0.VDDE.n115 digital_0.VDDE.n16 2.80353
R236 digital_0.VDDE.n108 digital_0.VDDE.n16 2.80353
R237 digital_0.VDDE.n107 digital_0.VDDE.n13 2.80353
R238 digital_0.VDDE.n108 digital_0.VDDE.n107 2.80353
R239 digital_0.VDDE.n2 digital_0.VDDE.n12 2.65147
R240 digital_0.VDDE.n64 digital_0.VDDE.n46 2.6245
R241 digital_0.VDDE.n118 digital_0.VDDE.n12 2.56843
R242 digital_0.VDDE.n118 digital_0.VDDE.n117 2.48542
R243 pmos_current_bgr_2_0.VDDE digital_0.VDDE.n25 2.46517
R244 digital_0.pmos_ena_0.VDDE digital_0.VDDE.n5 2.40529
R245 digital_0.VDDE.n85 digital_0.VDDE.n84 2.03039
R246 digital_0.VDDE.n2 digital_0.VDDE.n3 0.976616
R247 digital_0.VDDE.n94 digital_0.VDDE.n45 1.50638
R248 digital_0.VDDE.n99 digital_0.VDDE.n98 1.50638
R249 digital_0.VDDE.n99 digital_0.VDDE.n44 1.45719
R250 digital_0.VDDE.n79 digital_0.VDDE.n44 1.45719
R251 digital_0.VDDE.n45 digital_0.VDDE.n43 1.45719
R252 digital_0.VDDE.n79 digital_0.VDDE.n43 1.45719
R253 digital_0.VDDE.n113 digital_0.VDDE.n112 1.33202
R254 digital_0.VDDE.n114 digital_0.VDDE.n113 1.23963
R255 digital_0.VDDE.n52 digital_0.VDDE.n50 1.13031
R256 digital_0.VDDE.n91 digital_0.VDDE.n89 1.13031
R257 digital_0.VDDE.n74 digital_0.VDDE.n73 1.08707
R258 digital_0.VDDE.n26 digital_0.VDDE.n4 0.845955
R259 digital_0.VDDE.n75 digital_0.VDDE.n74 0.7755
R260 digital_0.VDDE.n84 digital_0.VDDE.n83 0.7755
R261 digital_0.VDDE.n5 digital_0.VDDE.n119 0.708631
R262 digital_0.VDDE.n86 digital_0.VDDE.n85 0.663329
R263 digital_0.VDDE.n7 digital_0.VDDE.n55 0.639087
R264 digital_0.VDDE.n61 digital_0.VDDE.n6 0.63637
R265 digital_0.VDDE.n113 digital_0.VDDE.n12 0.626276
R266 digital_0.VDDE.n114 digital_0.VDDE.n24 0.566321
R267 digital_0.VDDE.n95 digital_0.VDDE.n53 0.552734
R268 digital_0.VDDE.n93 digital_0.VDDE.n92 0.552734
R269 digital_0.VDDE.n97 digital_0.VDDE.n48 0.550017
R270 digital_0.VDDE.n87 pmos_current_bgr_0.vdde 0.550017
R271 digital_0.VDDE.n19 pmos_current_bgr_2_0.vdde 0.520126
R272 digital_0.VDDE.n68 digital_0.VDDE.n65 0.504571
R273 digital_0.VDDE.n85 digital_0.VDDE.n6 0.413543
R274 pmos_iptat_0.VDDE digital_0.VDDE.n69 0.396812
R275 digital_0.VDDE.n1 digital_0.VDDE.n0 0.019801
R276 digital_0.VDDE.n55 digital_0.VDDE.n54 0.383652
R277 digital_0.VDDE.n61 digital_0.VDDE.n60 0.383652
R278 digital_0.VDDE.n25 digital_0.VDDE.n15 0.3725
R279 digital_0.VDDE.n117 digital_0.VDDE.n116 0.3725
R280 digital_0.VDDE.n100 digital_0.VDDE.n46 0.344944
R281 digital_0.VDDE.n96 digital_0.VDDE.n47 0.344944
R282 digital_0.VDDE.n33 pmos_startup_0.VDDE 0.289147
R283 digital_0.VDDE.n39 digital_0.VDDE.n38 0.224218
R284 digital_0.VDDE.n5 digital_0.VDDE.n9 0.203505
R285 digital_0.VDDE.n40 pmos_startup_0.VDDE 0.175293
R286 digital_0.VDDE.n70 digital_0.VDDE.n65 0.148119
R287 digital_0.VDDE.n112 digital_0.VDDE.n111 0.148119
R288 digital_0.VDDE.n115 digital_0.VDDE.n114 0.143577
R289 digital_0.pmos_ena_0.VDDE digital_0.VDDE.n122 0.139087
R290 digital_0.VDDE.n3 digital_0.VDDE.n27 0.879945
R291 digital_0.VDDE.n71 pmos_iptat_0.VDDE 0.206309
R292 digital_0.VDDE.n13 pmos_current_bgr_2_0.vdde 0.189773
R293 digital_0.VDDE.n0 digital_0.VDDE.n118 0.130524
R294 digital_0.VDDE.n38 digital_0.VDDE.n30 0.0937836
R295 digital_0.VDDE.n7 digital_0.VDDE.n94 0.0875991
R296 digital_0.VDDE.n98 digital_0.VDDE.n6 0.0875991
R297 digital_0.VDDE.n2 digital_0.VDDE.n1 0.0618269
R298 digital_0.VDDE.n73 digital_0.VDDE.n0 0.0816518
R299 digital_0.VDDE.n73 digital_0.VDDE.n64 0.0775833
R300 pmos_current_bgr_2_0.D3.n3 pmos_current_bgr_2_0.D3.t1 1051.12
R301 pmos_current_bgr_2_0.D3.n5 pmos_current_bgr_2_0.D3.n4 1051.12
R302 pmos_current_bgr_2_0.D3.t3 pmos_current_bgr_2_0.D3.n6 1051.12
R303 pmos_current_bgr_2_0.D3.n8 pmos_current_bgr_2_0.D3.t5 402.695
R304 pmos_current_bgr_2_0.D3.n11 pmos_current_bgr_2_0.D3.t11 402.695
R305 pmos_current_bgr_2_0.D3.n7 pmos_current_bgr_2_0.D3.t13 387.759
R306 pmos_current_bgr_2_0.D3.n2 pmos_current_bgr_2_0.D3.t8 387.759
R307 pmos_current_bgr_2_0.D3.n8 pmos_current_bgr_2_0.D3.t7 227.323
R308 pmos_current_bgr_2_0.D3.t12 pmos_current_bgr_2_0.D3.n11 227.323
R309 pmos_current_bgr_2_0.D3.n10 pmos_current_bgr_2_0.D3.n9 199.65
R310 pmos_current_bgr_2_0.D3.n13 pmos_current_bgr_2_0.D3.n12 199.65
R311 pmos_current_bgr_2_0.D3.n0 pmos_current_bgr_2_0.D3.t14 83.7172
R312 pmos_current_bgr_2_0.D3.n0 pmos_current_bgr_2_0.D3.t4 83.7172
R313 pmos_current_bgr_2_0.D3.n1 pmos_current_bgr_2_0.D3.t2 83.7172
R314 pmos_current_bgr_2_0.D3.n1 pmos_current_bgr_2_0.D3.t10 83.7172
R315 pmos_current_bgr_2_0.D3.n2 pmos_current_bgr_2_0.D3.t9 82.8128
R316 pmos_current_bgr_2_0.D3.n7 pmos_current_bgr_2_0.D3.t15 82.8128
R317 pmos_current_bgr_2_0.D3.n9 pmos_current_bgr_2_0.D3.t0 28.5655
R318 pmos_current_bgr_2_0.D3.n9 pmos_current_bgr_2_0.D3.t6 28.5655
R319 pmos_current_bgr_2_0.D3.n12 pmos_current_bgr_2_0.D3.t12 28.5655
R320 pmos_current_bgr_2_0.D3.n12 pmos_current_bgr_2_0.D3.t16 28.5655
R321 pmos_current_bgr_2_0.D3.n0 pmos_current_bgr_2_0.D3.n14 12.1496
R322 pmos_current_bgr_2_0.D3.t1 pmos_current_bgr_2_0.D3.n1 11.2067
R323 pmos_current_bgr_2_0.D3.n0 pmos_current_bgr_2_0.D3.t3 11.1977
R324 pmos_current_bgr_2_0.D3.n14 pmos_current_bgr_2_0.D3.n13 4.29736
R325 pmos_current_bgr_2_0.D3.n14 pmos_current_bgr_2_0.D3 4.21562
R326 pmos_current_bgr_2_0.D3 pmos_current_bgr_2_0.D3.n10 4.03965
R327 pmos_current_bgr_2_0.D3.n3 pmos_current_bgr_2_0.D3.t20 1.2055
R328 pmos_current_bgr_2_0.D3.t1 pmos_current_bgr_2_0.D3.t19 1.2055
R329 pmos_current_bgr_2_0.D3.n5 pmos_current_bgr_2_0.D3.t19 1.2055
R330 pmos_current_bgr_2_0.D3.t22 pmos_current_bgr_2_0.D3.n3 1.2055
R331 pmos_current_bgr_2_0.D3.n4 pmos_current_bgr_2_0.D3.t22 1.2055
R332 pmos_current_bgr_2_0.D3.n4 pmos_current_bgr_2_0.D3.t18 1.2055
R333 pmos_current_bgr_2_0.D3.t3 pmos_current_bgr_2_0.D3.t18 1.2055
R334 pmos_current_bgr_2_0.D3.t21 pmos_current_bgr_2_0.D3.n5 1.2055
R335 pmos_current_bgr_2_0.D3.n6 pmos_current_bgr_2_0.D3.t21 1.2055
R336 pmos_current_bgr_2_0.D3.n6 pmos_current_bgr_2_0.D3.t17 1.2055
R337 pmos_current_bgr_2_0.D3.n1 pmos_current_bgr_2_0.D3.n2 0.732467
R338 pmos_current_bgr_2_0.D3.n0 pmos_current_bgr_2_0.D3.n7 0.732467
R339 pmos_current_bgr_2_0.D3.n10 pmos_current_bgr_2_0.D3.n8 0.610083
R340 pmos_current_bgr_2_0.D3.n13 pmos_current_bgr_2_0.D3.n11 0.610083
R341 AVSS.n6055 AVSS.n5928 135808
R342 AVSS.n5990 AVSS.n5967 80943.8
R343 AVSS.n5990 AVSS.n295 80943.8
R344 AVSS.n5967 AVSS.n5965 80938
R345 AVSS.n5965 AVSS.n295 80938
R346 AVSS.n5980 AVSS.n293 67287.1
R347 AVSS.n6059 AVSS.n293 67287.1
R348 AVSS.n5980 AVSS.n294 67287.1
R349 AVSS.n6059 AVSS.n294 67287.1
R350 AVSS.n5993 AVSS.n5961 49951.1
R351 AVSS.n5993 AVSS.n5962 49951.1
R352 AVSS.n5997 AVSS.n5961 49951.1
R353 AVSS.n5997 AVSS.n5962 49951.1
R354 AVSS.n6056 AVSS.n6055 34523.1
R355 AVSS.n6032 AVSS.n5938 30453.9
R356 AVSS.n6035 AVSS.n5938 30453.9
R357 AVSS.n6032 AVSS.n5939 30326.4
R358 AVSS.n6035 AVSS.n5939 30326.4
R359 AVSS.n6015 AVSS.n6012 19445.1
R360 AVSS.n6015 AVSS.n6008 19445.1
R361 AVSS.n6022 AVSS.n6012 19445.1
R362 AVSS.n6022 AVSS.n6008 19445.1
R363 AVSS.n6162 AVSS.n6161 18756
R364 AVSS.n6057 AVSS.n6056 18401.6
R365 AVSS.n5674 AVSS.n5673 15929.3
R366 AVSS.n6017 AVSS.n5929 14213
R367 AVSS.n6053 AVSS.n5929 14213
R368 AVSS.n6017 AVSS.n5930 14213
R369 AVSS.n6053 AVSS.n5930 14213
R370 AVSS.n5989 AVSS.n5968 5259.29
R371 AVSS.n5989 AVSS.n5988 5259.29
R372 AVSS.n5987 AVSS.n5968 5258.92
R373 AVSS.n5988 AVSS.n5987 5258.92
R374 AVSS.n5947 AVSS.n5943 4797.53
R375 AVSS.n5959 AVSS.n5943 4768.56
R376 AVSS.n5959 AVSS.n5944 4768.56
R377 AVSS.n5947 AVSS.n5944 4739.59
R378 AVSS.n5981 AVSS.n291 4371.95
R379 AVSS.n6060 AVSS.n291 4371.95
R380 AVSS.n5981 AVSS.n292 4371.95
R381 AVSS.n6060 AVSS.n292 4371.95
R382 AVSS.n5994 AVSS.n5963 3245.55
R383 AVSS.n5995 AVSS.n5994 3245.55
R384 AVSS.n5996 AVSS.n5963 3245.55
R385 AVSS.n5996 AVSS.n5995 3245.55
R386 AVSS.n5966 AVSS.t16 3243.42
R387 AVSS.n3591 AVSS.n3575 2225.3
R388 AVSS.n5675 AVSS.n5674 2157.28
R389 AVSS.n5701 AVSS.n399 2157.28
R390 AVSS.n859 AVSS.n858 2157.28
R391 AVSS.n886 AVSS.n885 2157.28
R392 AVSS.n1320 AVSS.n1319 2157.28
R393 AVSS.n1345 AVSS.n1132 2157.28
R394 AVSS.n3244 AVSS.n3243 2157.28
R395 AVSS.n3270 AVSS.n2982 2157.28
R396 AVSS.n6186 AVSS.n161 2157.28
R397 AVSS.n858 AVSS.n399 2135.92
R398 AVSS.n1319 AVSS.n886 2135.92
R399 AVSS.n3243 AVSS.n1132 2135.92
R400 AVSS.n2982 AVSS.n161 2135.92
R401 AVSS.n5701 AVSS.n5700 2050.49
R402 AVSS.n885 AVSS.n668 2050.49
R403 AVSS.n1345 AVSS.n1344 2050.49
R404 AVSS.n3270 AVSS.n3269 2050.49
R405 AVSS.n6162 AVSS.n173 2050.49
R406 AVSS.n6030 AVSS.n5936 1974.59
R407 AVSS.n6037 AVSS.n5936 1974.59
R408 AVSS.n6031 AVSS.n5937 1970.45
R409 AVSS.n6036 AVSS.n5937 1970.45
R410 AVSS.n6058 AVSS.t16 1925.32
R411 AVSS.n5675 AVSS.n5639 1922.33
R412 AVSS.n5681 AVSS.n5639 1922.33
R413 AVSS.n5682 AVSS.n5681 1922.33
R414 AVSS.n5684 AVSS.n5682 1922.33
R415 AVSS.n5684 AVSS.n5683 1922.33
R416 AVSS.n5691 AVSS.n5690 1922.33
R417 AVSS.n5692 AVSS.n5691 1922.33
R418 AVSS.n5692 AVSS.n5632 1922.33
R419 AVSS.n5699 AVSS.n5632 1922.33
R420 AVSS.n5700 AVSS.n5699 1922.33
R421 AVSS.n860 AVSS.n859 1922.33
R422 AVSS.n860 AVSS.n678 1922.33
R423 AVSS.n867 AVSS.n678 1922.33
R424 AVSS.n868 AVSS.n867 1922.33
R425 AVSS.n869 AVSS.n868 1922.33
R426 AVSS.n871 AVSS.n674 1922.33
R427 AVSS.n877 AVSS.n674 1922.33
R428 AVSS.n878 AVSS.n877 1922.33
R429 AVSS.n879 AVSS.n878 1922.33
R430 AVSS.n879 AVSS.n668 1922.33
R431 AVSS.n1320 AVSS.n1156 1922.33
R432 AVSS.n1326 AVSS.n1156 1922.33
R433 AVSS.n1327 AVSS.n1326 1922.33
R434 AVSS.n1329 AVSS.n1327 1922.33
R435 AVSS.n1329 AVSS.n1328 1922.33
R436 AVSS.n1336 AVSS.n297 1922.33
R437 AVSS.n1336 AVSS.n1150 1922.33
R438 AVSS.n1343 AVSS.n1150 1922.33
R439 AVSS.n1344 AVSS.n1343 1922.33
R440 AVSS.n3244 AVSS.n3082 1922.33
R441 AVSS.n3250 AVSS.n3082 1922.33
R442 AVSS.n3251 AVSS.n3250 1922.33
R443 AVSS.n3253 AVSS.n3251 1922.33
R444 AVSS.n3253 AVSS.n3252 1922.33
R445 AVSS.n3260 AVSS.n3259 1922.33
R446 AVSS.n3261 AVSS.n3260 1922.33
R447 AVSS.n3261 AVSS.n3075 1922.33
R448 AVSS.n3268 AVSS.n3075 1922.33
R449 AVSS.n3269 AVSS.n3268 1922.33
R450 AVSS.n6186 AVSS.n6185 1922.33
R451 AVSS.n6185 AVSS.n6184 1922.33
R452 AVSS.n6184 AVSS.n162 1922.33
R453 AVSS.n6178 AVSS.n162 1922.33
R454 AVSS.n6178 AVSS.n6177 1922.33
R455 AVSS.n6176 AVSS.n169 1922.33
R456 AVSS.n6170 AVSS.n169 1922.33
R457 AVSS.n6170 AVSS.n6169 1922.33
R458 AVSS.n6169 AVSS.n6168 1922.33
R459 AVSS.n6168 AVSS.n173 1922.33
R460 AVSS.n6058 AVSS.t17 1819.95
R461 AVSS.n5927 AVSS.n296 1794.17
R462 AVSS.t17 AVSS.n6057 1712.84
R463 AVSS.n6011 AVSS.n6007 1263.44
R464 AVSS.n6024 AVSS.n6007 1263.44
R465 AVSS.n6023 AVSS.n6011 1263.44
R466 AVSS.n6024 AVSS.n6023 1263.44
R467 AVSS.n5991 AVSS.t13 1191.99
R468 AVSS.t10 AVSS.n5991 1067.61
R469 AVSS.n5690 AVSS.t90 1003.88
R470 AVSS.n871 AVSS.t80 1003.88
R471 AVSS.t78 AVSS.n296 1003.88
R472 AVSS.n3259 AVSS.t76 1003.88
R473 AVSS.t85 AVSS.n6176 1003.88
R474 AVSS.n5933 AVSS.n5931 923.482
R475 AVSS.n6052 AVSS.n5931 923.482
R476 AVSS.n6051 AVSS.n5933 923.482
R477 AVSS.n6052 AVSS.n6051 923.482
R478 AVSS.n5683 AVSS.t90 918.447
R479 AVSS.n869 AVSS.t80 918.447
R480 AVSS.n1328 AVSS.t78 918.447
R481 AVSS.n3252 AVSS.t76 918.447
R482 AVSS.n6177 AVSS.t85 918.447
R483 AVSS.n5926 AVSS.n5925 684.131
R484 AVSS.t13 AVSS.t6 680.644
R485 AVSS.t117 AVSS.t123 663.428
R486 AVSS.n6056 AVSS.n5927 597.168
R487 AVSS.n5912 AVSS.n5911 589.519
R488 AVSS.n5569 AVSS.n5447 585
R489 AVSS.n5568 AVSS.n5567 585
R490 AVSS.n5449 AVSS.n5448 585
R491 AVSS.n5563 AVSS.n5562 585
R492 AVSS.n5561 AVSS.n5454 585
R493 AVSS.n5560 AVSS.n5559 585
R494 AVSS.n5558 AVSS.n5557 585
R495 AVSS.n5556 AVSS.n5555 585
R496 AVSS.n5554 AVSS.n5553 585
R497 AVSS.n5552 AVSS.n5551 585
R498 AVSS.n5550 AVSS.n5549 585
R499 AVSS.n5257 AVSS.n5255 585
R500 AVSS.n5420 AVSS.n5419 585
R501 AVSS.n5422 AVSS.n5299 585
R502 AVSS.n5425 AVSS.n5424 585
R503 AVSS.n5426 AVSS.n5298 585
R504 AVSS.n5428 AVSS.n5427 585
R505 AVSS.n5430 AVSS.n5297 585
R506 AVSS.n5433 AVSS.n5432 585
R507 AVSS.n5434 AVSS.n5296 585
R508 AVSS.n5436 AVSS.n5435 585
R509 AVSS.n5438 AVSS.n5295 585
R510 AVSS.n5441 AVSS.n5440 585
R511 AVSS.n5442 AVSS.n5281 585
R512 AVSS.n6279 AVSS.n6278 585
R513 AVSS.n6281 AVSS.n10 585
R514 AVSS.n6284 AVSS.n6283 585
R515 AVSS.n6285 AVSS.n9 585
R516 AVSS.n6287 AVSS.n6286 585
R517 AVSS.n6289 AVSS.n8 585
R518 AVSS.n6292 AVSS.n6291 585
R519 AVSS.n6293 AVSS.n7 585
R520 AVSS.n6295 AVSS.n6294 585
R521 AVSS.n6297 AVSS.n6 585
R522 AVSS.n6298 AVSS.n2 585
R523 AVSS.n6301 AVSS.n6300 585
R524 AVSS.n5223 AVSS.n409 585
R525 AVSS.n5197 AVSS.n410 585
R526 AVSS.n5199 AVSS.n5198 585
R527 AVSS.n5201 AVSS.n5200 585
R528 AVSS.n5203 AVSS.n5202 585
R529 AVSS.n5205 AVSS.n5204 585
R530 AVSS.n5207 AVSS.n5206 585
R531 AVSS.n5209 AVSS.n5208 585
R532 AVSS.n5211 AVSS.n5210 585
R533 AVSS.n5213 AVSS.n5212 585
R534 AVSS.n5215 AVSS.n5214 585
R535 AVSS.n5216 AVSS.n418 585
R536 AVSS.n5879 AVSS.n5878 585
R537 AVSS.n5881 AVSS.n322 585
R538 AVSS.n5883 AVSS.n5882 585
R539 AVSS.n5884 AVSS.n321 585
R540 AVSS.n5886 AVSS.n5885 585
R541 AVSS.n5888 AVSS.n319 585
R542 AVSS.n5890 AVSS.n5889 585
R543 AVSS.n5891 AVSS.n318 585
R544 AVSS.n5893 AVSS.n5892 585
R545 AVSS.n5895 AVSS.n315 585
R546 AVSS.n5897 AVSS.n5896 585
R547 AVSS.n5898 AVSS.n314 585
R548 AVSS.n5093 AVSS.n5092 585
R549 AVSS.n5091 AVSS.n427 585
R550 AVSS.n5090 AVSS.n5089 585
R551 AVSS.n5088 AVSS.n5087 585
R552 AVSS.n5086 AVSS.n5085 585
R553 AVSS.n5084 AVSS.n5083 585
R554 AVSS.n5082 AVSS.n5081 585
R555 AVSS.n5080 AVSS.n5079 585
R556 AVSS.n5078 AVSS.n5077 585
R557 AVSS.n422 AVSS.n421 585
R558 AVSS.n5098 AVSS.n5097 585
R559 AVSS.n408 AVSS.n406 585
R560 AVSS.n5900 AVSS.n5899 585
R561 AVSS.n5901 AVSS.n5900 585
R562 AVSS.n312 AVSS.n311 585
R563 AVSS.n5902 AVSS.n312 585
R564 AVSS.n5905 AVSS.n5904 585
R565 AVSS.n5904 AVSS.n5903 585
R566 AVSS.n5906 AVSS.n310 585
R567 AVSS.n310 AVSS.n309 585
R568 AVSS.n5908 AVSS.n5907 585
R569 AVSS.n5909 AVSS.n5908 585
R570 AVSS.n308 AVSS.n307 585
R571 AVSS.n5910 AVSS.n308 585
R572 AVSS.n5218 AVSS.n5217 585
R573 AVSS.n5219 AVSS.n5218 585
R574 AVSS.n419 AVSS.n417 585
R575 AVSS.n417 AVSS.n416 585
R576 AVSS.n439 AVSS.n438 585
R577 AVSS.n440 AVSS.n439 585
R578 AVSS.n443 AVSS.n442 585
R579 AVSS.n442 AVSS.n441 585
R580 AVSS.n444 AVSS.n437 585
R581 AVSS.n437 AVSS.n436 585
R582 AVSS.n446 AVSS.n445 585
R583 AVSS.n447 AVSS.n446 585
R584 AVSS.n435 AVSS.n434 585
R585 AVSS.n448 AVSS.n435 585
R586 AVSS.n5067 AVSS.n5066 585
R587 AVSS.n5066 AVSS.n5065 585
R588 AVSS.n5068 AVSS.n433 585
R589 AVSS.n433 AVSS.n432 585
R590 AVSS.n5070 AVSS.n5069 585
R591 AVSS.n5071 AVSS.n5070 585
R592 AVSS.n430 AVSS.n429 585
R593 AVSS.n5072 AVSS.n430 585
R594 AVSS.n5075 AVSS.n5074 585
R595 AVSS.n5074 AVSS.n5073 585
R596 AVSS.n5076 AVSS.n428 585
R597 AVSS.n431 AVSS.n428 585
R598 AVSS.n5444 AVSS.n5443 585
R599 AVSS.n5445 AVSS.n5444 585
R600 AVSS.n5294 AVSS.n5280 585
R601 AVSS.n5280 AVSS.n5279 585
R602 AVSS.n5293 AVSS.n5292 585
R603 AVSS.n5292 AVSS.n5291 585
R604 AVSS.n5283 AVSS.n5282 585
R605 AVSS.n5290 AVSS.n5283 585
R606 AVSS.n5288 AVSS.n5287 585
R607 AVSS.n5289 AVSS.n5288 585
R608 AVSS.n5286 AVSS.n5285 585
R609 AVSS.n5285 AVSS.n5284 585
R610 AVSS.n18 AVSS.n17 585
R611 AVSS.n19 AVSS.n18 585
R612 AVSS.n6268 AVSS.n6267 585
R613 AVSS.n6267 AVSS.n6266 585
R614 AVSS.n6269 AVSS.n16 585
R615 AVSS.n16 AVSS.n15 585
R616 AVSS.n6271 AVSS.n6270 585
R617 AVSS.n6272 AVSS.n6271 585
R618 AVSS.n13 AVSS.n12 585
R619 AVSS.n6273 AVSS.n13 585
R620 AVSS.n6276 AVSS.n6275 585
R621 AVSS.n6275 AVSS.n6274 585
R622 AVSS.n6277 AVSS.n11 585
R623 AVSS.n14 AVSS.n11 585
R624 AVSS.n5615 AVSS.n5614 585
R625 AVSS.n5616 AVSS.n5615 585
R626 AVSS.n5593 AVSS.n5266 585
R627 AVSS.n5266 AVSS.n5265 585
R628 AVSS.n5592 AVSS.n5591 585
R629 AVSS.n5591 AVSS.n5590 585
R630 AVSS.n5269 AVSS.n5268 585
R631 AVSS.n5589 AVSS.n5269 585
R632 AVSS.n5587 AVSS.n5586 585
R633 AVSS.n5588 AVSS.n5587 585
R634 AVSS.n5585 AVSS.n5271 585
R635 AVSS.n5271 AVSS.n5270 585
R636 AVSS.n5584 AVSS.n5583 585
R637 AVSS.n5583 AVSS.n5582 585
R638 AVSS.n5273 AVSS.n5272 585
R639 AVSS.n5581 AVSS.n5273 585
R640 AVSS.n5579 AVSS.n5578 585
R641 AVSS.n5580 AVSS.n5579 585
R642 AVSS.n5577 AVSS.n5275 585
R643 AVSS.n5275 AVSS.n5274 585
R644 AVSS.n5576 AVSS.n5575 585
R645 AVSS.n5575 AVSS.n5574 585
R646 AVSS.n5277 AVSS.n5276 585
R647 AVSS.n5573 AVSS.n5277 585
R648 AVSS.n5571 AVSS.n5570 585
R649 AVSS.n5572 AVSS.n5571 585
R650 AVSS.n5847 AVSS.n5258 585
R651 AVSS.n5594 AVSS.n5259 585
R652 AVSS.n5596 AVSS.n5595 585
R653 AVSS.n5598 AVSS.n5597 585
R654 AVSS.n5600 AVSS.n5599 585
R655 AVSS.n5602 AVSS.n5601 585
R656 AVSS.n5604 AVSS.n5603 585
R657 AVSS.n5606 AVSS.n5605 585
R658 AVSS.n5608 AVSS.n5607 585
R659 AVSS.n5610 AVSS.n5609 585
R660 AVSS.n5612 AVSS.n5611 585
R661 AVSS.n5613 AVSS.n5267 585
R662 AVSS.n5841 AVSS.n5840 585
R663 AVSS.n5839 AVSS.n5623 585
R664 AVSS.n5838 AVSS.n5837 585
R665 AVSS.n5836 AVSS.n5835 585
R666 AVSS.n5834 AVSS.n5833 585
R667 AVSS.n5832 AVSS.n5831 585
R668 AVSS.n5830 AVSS.n5829 585
R669 AVSS.n5828 AVSS.n5827 585
R670 AVSS.n5826 AVSS.n5825 585
R671 AVSS.n5824 AVSS.n5823 585
R672 AVSS.n5822 AVSS.n5821 585
R673 AVSS.n5627 AVSS.n5626 585
R674 AVSS.n5672 AVSS.n5671 585
R675 AVSS.n5673 AVSS.n5672 585
R676 AVSS.n5670 AVSS.n5644 585
R677 AVSS.n5644 AVSS.n5643 585
R678 AVSS.n5669 AVSS.n5668 585
R679 AVSS.n5668 AVSS.n5667 585
R680 AVSS.n5646 AVSS.n5645 585
R681 AVSS.n5666 AVSS.n5646 585
R682 AVSS.n5664 AVSS.n5663 585
R683 AVSS.n5665 AVSS.n5664 585
R684 AVSS.n5662 AVSS.n5647 585
R685 AVSS.n5647 AVSS.n37 585
R686 AVSS.n5661 AVSS.n5660 585
R687 AVSS.n5660 AVSS.n36 585
R688 AVSS.n5659 AVSS.n5648 585
R689 AVSS.n5659 AVSS.n5658 585
R690 AVSS.n5653 AVSS.n5649 585
R691 AVSS.n5657 AVSS.n5649 585
R692 AVSS.n5655 AVSS.n5654 585
R693 AVSS.n5656 AVSS.n5655 585
R694 AVSS.n5652 AVSS.n5651 585
R695 AVSS.n5651 AVSS.n5650 585
R696 AVSS.n5625 AVSS.n5624 585
R697 AVSS.n5624 AVSS.n5617 585
R698 AVSS.n1587 AVSS.n1384 585
R699 AVSS.n1585 AVSS.n1584 585
R700 AVSS.n1583 AVSS.n1385 585
R701 AVSS.n1582 AVSS.n1581 585
R702 AVSS.n1579 AVSS.n1386 585
R703 AVSS.n1577 AVSS.n1576 585
R704 AVSS.n1575 AVSS.n1387 585
R705 AVSS.n1574 AVSS.n1573 585
R706 AVSS.n1571 AVSS.n1388 585
R707 AVSS.n1569 AVSS.n1568 585
R708 AVSS.n1567 AVSS.n1389 585
R709 AVSS.n1566 AVSS.n1565 585
R710 AVSS.n2363 AVSS.n2362 585
R711 AVSS.n2360 AVSS.n2310 585
R712 AVSS.n2359 AVSS.n2358 585
R713 AVSS.n2357 AVSS.n2356 585
R714 AVSS.n2355 AVSS.n2312 585
R715 AVSS.n2353 AVSS.n2352 585
R716 AVSS.n2351 AVSS.n2313 585
R717 AVSS.n2350 AVSS.n2349 585
R718 AVSS.n2347 AVSS.n2314 585
R719 AVSS.n2345 AVSS.n2344 585
R720 AVSS.n2343 AVSS.n2315 585
R721 AVSS.n2341 AVSS.n2340 585
R722 AVSS.n2413 AVSS.n2412 585
R723 AVSS.n2409 AVSS.n2303 585
R724 AVSS.n2408 AVSS.n2407 585
R725 AVSS.n2406 AVSS.n2405 585
R726 AVSS.n2404 AVSS.n2306 585
R727 AVSS.n2402 AVSS.n2401 585
R728 AVSS.n2400 AVSS.n2307 585
R729 AVSS.n2399 AVSS.n2398 585
R730 AVSS.n2396 AVSS.n2308 585
R731 AVSS.n2394 AVSS.n2393 585
R732 AVSS.n2392 AVSS.n2309 585
R733 AVSS.n2391 AVSS.n2390 585
R734 AVSS.n2279 AVSS.n2278 585
R735 AVSS.n2281 AVSS.n2200 585
R736 AVSS.n2284 AVSS.n2283 585
R737 AVSS.n2285 AVSS.n2199 585
R738 AVSS.n2287 AVSS.n2286 585
R739 AVSS.n2289 AVSS.n2198 585
R740 AVSS.n2292 AVSS.n2291 585
R741 AVSS.n2293 AVSS.n2197 585
R742 AVSS.n2295 AVSS.n2294 585
R743 AVSS.n2297 AVSS.n2196 585
R744 AVSS.n2300 AVSS.n2299 585
R745 AVSS.n973 AVSS.n971 585
R746 AVSS.n2233 AVSS.n2232 585
R747 AVSS.n2234 AVSS.n2208 585
R748 AVSS.n2236 AVSS.n2235 585
R749 AVSS.n2238 AVSS.n2206 585
R750 AVSS.n2240 AVSS.n2239 585
R751 AVSS.n2241 AVSS.n2205 585
R752 AVSS.n2243 AVSS.n2242 585
R753 AVSS.n2245 AVSS.n2203 585
R754 AVSS.n2247 AVSS.n2246 585
R755 AVSS.n2248 AVSS.n2202 585
R756 AVSS.n2250 AVSS.n2249 585
R757 AVSS.n2252 AVSS.n2201 585
R758 AVSS.n693 AVSS.n692 585
R759 AVSS.n694 AVSS.n689 585
R760 AVSS.n696 AVSS.n695 585
R761 AVSS.n698 AVSS.n688 585
R762 AVSS.n701 AVSS.n700 585
R763 AVSS.n702 AVSS.n687 585
R764 AVSS.n704 AVSS.n703 585
R765 AVSS.n706 AVSS.n686 585
R766 AVSS.n709 AVSS.n708 585
R767 AVSS.n710 AVSS.n685 585
R768 AVSS.n712 AVSS.n711 585
R769 AVSS.n714 AVSS.n684 585
R770 AVSS.n1563 AVSS.n1562 585
R771 AVSS.n1561 AVSS.n1560 585
R772 AVSS.n1559 AVSS.n1558 585
R773 AVSS.n1557 AVSS.n1556 585
R774 AVSS.n1555 AVSS.n1554 585
R775 AVSS.n1553 AVSS.n1552 585
R776 AVSS.n1551 AVSS.n1550 585
R777 AVSS.n1549 AVSS.n1548 585
R778 AVSS.n1547 AVSS.n1546 585
R779 AVSS.n1545 AVSS.n1544 585
R780 AVSS.n1543 AVSS.n1542 585
R781 AVSS.n1541 AVSS.n1540 585
R782 AVSS.n1539 AVSS.n613 585
R783 AVSS.n5016 AVSS.n613 585
R784 AVSS.n2388 AVSS.n2387 585
R785 AVSS.n2386 AVSS.n2385 585
R786 AVSS.n2384 AVSS.n2383 585
R787 AVSS.n2382 AVSS.n2381 585
R788 AVSS.n2380 AVSS.n2379 585
R789 AVSS.n2378 AVSS.n2377 585
R790 AVSS.n2376 AVSS.n2375 585
R791 AVSS.n2374 AVSS.n2373 585
R792 AVSS.n2372 AVSS.n2371 585
R793 AVSS.n2370 AVSS.n2369 585
R794 AVSS.n2368 AVSS.n2367 585
R795 AVSS.n2366 AVSS.n2365 585
R796 AVSS.n2364 AVSS.n626 585
R797 AVSS.n5016 AVSS.n626 585
R798 AVSS.n2254 AVSS.n2253 585
R799 AVSS.n2256 AVSS.n2255 585
R800 AVSS.n2258 AVSS.n2257 585
R801 AVSS.n2260 AVSS.n2259 585
R802 AVSS.n2262 AVSS.n2261 585
R803 AVSS.n2264 AVSS.n2263 585
R804 AVSS.n2266 AVSS.n2265 585
R805 AVSS.n2268 AVSS.n2267 585
R806 AVSS.n2270 AVSS.n2269 585
R807 AVSS.n2272 AVSS.n2271 585
R808 AVSS.n2274 AVSS.n2273 585
R809 AVSS.n2276 AVSS.n2275 585
R810 AVSS.n2277 AVSS.n606 585
R811 AVSS.n5016 AVSS.n606 585
R812 AVSS.n855 AVSS.n682 585
R813 AVSS.n854 AVSS.n853 585
R814 AVSS.n852 AVSS.n851 585
R815 AVSS.n850 AVSS.n849 585
R816 AVSS.n848 AVSS.n847 585
R817 AVSS.n846 AVSS.n845 585
R818 AVSS.n844 AVSS.n843 585
R819 AVSS.n842 AVSS.n841 585
R820 AVSS.n840 AVSS.n839 585
R821 AVSS.n838 AVSS.n837 585
R822 AVSS.n836 AVSS.n835 585
R823 AVSS.n690 AVSS.n683 585
R824 AVSS.n5877 AVSS.n324 585
R825 AVSS.n5876 AVSS.n5875 585
R826 AVSS.n376 AVSS.n327 585
R827 AVSS.n378 AVSS.n377 585
R828 AVSS.n380 AVSS.n379 585
R829 AVSS.n382 AVSS.n381 585
R830 AVSS.n384 AVSS.n383 585
R831 AVSS.n386 AVSS.n385 585
R832 AVSS.n388 AVSS.n387 585
R833 AVSS.n390 AVSS.n389 585
R834 AVSS.n392 AVSS.n391 585
R835 AVSS.n394 AVSS.n393 585
R836 AVSS.n395 AVSS.n340 585
R837 AVSS.n5873 AVSS.n340 585
R838 AVSS.n5225 AVSS.n5224 585
R839 AVSS.n5227 AVSS.n5226 585
R840 AVSS.n5229 AVSS.n5228 585
R841 AVSS.n5231 AVSS.n5230 585
R842 AVSS.n5233 AVSS.n5232 585
R843 AVSS.n5235 AVSS.n5234 585
R844 AVSS.n5237 AVSS.n5236 585
R845 AVSS.n5239 AVSS.n5238 585
R846 AVSS.n5241 AVSS.n5240 585
R847 AVSS.n5243 AVSS.n5242 585
R848 AVSS.n5245 AVSS.n5244 585
R849 AVSS.n5246 AVSS.n407 585
R850 AVSS.n5248 AVSS.n5247 585
R851 AVSS.n5873 AVSS.n5248 585
R852 AVSS.n5418 AVSS.n5300 585
R853 AVSS.n5417 AVSS.n5416 585
R854 AVSS.n5415 AVSS.n5414 585
R855 AVSS.n5413 AVSS.n5412 585
R856 AVSS.n5411 AVSS.n5410 585
R857 AVSS.n5409 AVSS.n5408 585
R858 AVSS.n5407 AVSS.n5406 585
R859 AVSS.n5405 AVSS.n5404 585
R860 AVSS.n5403 AVSS.n5402 585
R861 AVSS.n5401 AVSS.n5400 585
R862 AVSS.n5399 AVSS.n5398 585
R863 AVSS.n5397 AVSS.n5396 585
R864 AVSS.n4 AVSS.n3 585
R865 AVSS.n5873 AVSS.n4 585
R866 AVSS.n5849 AVSS.n5848 585
R867 AVSS.n5851 AVSS.n5850 585
R868 AVSS.n5853 AVSS.n5852 585
R869 AVSS.n5855 AVSS.n5854 585
R870 AVSS.n5857 AVSS.n5856 585
R871 AVSS.n5859 AVSS.n5858 585
R872 AVSS.n5861 AVSS.n5860 585
R873 AVSS.n5863 AVSS.n5862 585
R874 AVSS.n5865 AVSS.n5864 585
R875 AVSS.n5867 AVSS.n5866 585
R876 AVSS.n5869 AVSS.n5868 585
R877 AVSS.n5870 AVSS.n5256 585
R878 AVSS.n5872 AVSS.n5871 585
R879 AVSS.n5873 AVSS.n5872 585
R880 AVSS.n5704 AVSS.n5703 585
R881 AVSS.n5706 AVSS.n5705 585
R882 AVSS.n5708 AVSS.n5707 585
R883 AVSS.n5710 AVSS.n5709 585
R884 AVSS.n5712 AVSS.n5711 585
R885 AVSS.n5714 AVSS.n5713 585
R886 AVSS.n5716 AVSS.n5715 585
R887 AVSS.n5718 AVSS.n5717 585
R888 AVSS.n5720 AVSS.n5719 585
R889 AVSS.n5722 AVSS.n5721 585
R890 AVSS.n5724 AVSS.n5723 585
R891 AVSS.n5629 AVSS.n5628 585
R892 AVSS.n5015 AVSS.n5014 585
R893 AVSS.n5016 AVSS.n5015 585
R894 AVSS.n635 AVSS.n633 585
R895 AVSS.n901 AVSS.n900 585
R896 AVSS.n903 AVSS.n902 585
R897 AVSS.n905 AVSS.n904 585
R898 AVSS.n907 AVSS.n906 585
R899 AVSS.n909 AVSS.n908 585
R900 AVSS.n911 AVSS.n910 585
R901 AVSS.n913 AVSS.n912 585
R902 AVSS.n915 AVSS.n914 585
R903 AVSS.n917 AVSS.n916 585
R904 AVSS.n919 AVSS.n918 585
R905 AVSS.n920 AVSS.n899 585
R906 AVSS.n922 AVSS.n921 585
R907 AVSS.n924 AVSS.n898 585
R908 AVSS.n927 AVSS.n926 585
R909 AVSS.n928 AVSS.n897 585
R910 AVSS.n930 AVSS.n929 585
R911 AVSS.n932 AVSS.n896 585
R912 AVSS.n935 AVSS.n934 585
R913 AVSS.n936 AVSS.n895 585
R914 AVSS.n938 AVSS.n937 585
R915 AVSS.n940 AVSS.n894 585
R916 AVSS.n943 AVSS.n942 585
R917 AVSS.n944 AVSS.n892 585
R918 AVSS.n4994 AVSS.n4993 585
R919 AVSS.n4996 AVSS.n642 585
R920 AVSS.n4998 AVSS.n4997 585
R921 AVSS.n4999 AVSS.n641 585
R922 AVSS.n5001 AVSS.n5000 585
R923 AVSS.n5003 AVSS.n639 585
R924 AVSS.n5005 AVSS.n5004 585
R925 AVSS.n5006 AVSS.n638 585
R926 AVSS.n5008 AVSS.n5007 585
R927 AVSS.n5010 AVSS.n636 585
R928 AVSS.n5012 AVSS.n5011 585
R929 AVSS.n5013 AVSS.n634 585
R930 AVSS.n3121 AVSS.n3091 585
R931 AVSS.n3120 AVSS.n3119 585
R932 AVSS.n3117 AVSS.n3092 585
R933 AVSS.n3115 AVSS.n3114 585
R934 AVSS.n3113 AVSS.n3093 585
R935 AVSS.n3112 AVSS.n3111 585
R936 AVSS.n3109 AVSS.n3094 585
R937 AVSS.n3107 AVSS.n3106 585
R938 AVSS.n3105 AVSS.n3095 585
R939 AVSS.n3104 AVSS.n3103 585
R940 AVSS.n3101 AVSS.n3096 585
R941 AVSS.n3099 AVSS.n3098 585
R942 AVSS.n2898 AVSS.n2836 585
R943 AVSS.n2897 AVSS.n2896 585
R944 AVSS.n2895 AVSS.n2894 585
R945 AVSS.n2893 AVSS.n2892 585
R946 AVSS.n2891 AVSS.n2890 585
R947 AVSS.n2889 AVSS.n2888 585
R948 AVSS.n2887 AVSS.n2886 585
R949 AVSS.n2885 AVSS.n2884 585
R950 AVSS.n2883 AVSS.n2882 585
R951 AVSS.n2791 AVSS.n2790 585
R952 AVSS.n4501 AVSS.n4500 585
R953 AVSS.n4502 AVSS.n2789 585
R954 AVSS.n4674 AVSS.n2776 585
R955 AVSS.n4677 AVSS.n4676 585
R956 AVSS.n2778 AVSS.n2777 585
R957 AVSS.n2843 AVSS.n2842 585
R958 AVSS.n2845 AVSS.n2844 585
R959 AVSS.n2847 AVSS.n2840 585
R960 AVSS.n2850 AVSS.n2849 585
R961 AVSS.n2851 AVSS.n2839 585
R962 AVSS.n2853 AVSS.n2852 585
R963 AVSS.n2855 AVSS.n2838 585
R964 AVSS.n2856 AVSS.n2837 585
R965 AVSS.n2859 AVSS.n2858 585
R966 AVSS.n3039 AVSS.n3013 585
R967 AVSS.n3037 AVSS.n3036 585
R968 AVSS.n3035 AVSS.n3014 585
R969 AVSS.n3034 AVSS.n3033 585
R970 AVSS.n3031 AVSS.n3015 585
R971 AVSS.n3029 AVSS.n3028 585
R972 AVSS.n3027 AVSS.n3016 585
R973 AVSS.n3026 AVSS.n3025 585
R974 AVSS.n3023 AVSS.n3017 585
R975 AVSS.n3021 AVSS.n3020 585
R976 AVSS.n3019 AVSS.n1737 585
R977 AVSS.n4682 AVSS.n1736 585
R978 AVSS.n4706 AVSS.n1723 585
R979 AVSS.n4709 AVSS.n4708 585
R980 AVSS.n1725 AVSS.n1724 585
R981 AVSS.n2996 AVSS.n2995 585
R982 AVSS.n2998 AVSS.n2997 585
R983 AVSS.n3000 AVSS.n2993 585
R984 AVSS.n3003 AVSS.n3002 585
R985 AVSS.n3004 AVSS.n2992 585
R986 AVSS.n3006 AVSS.n3005 585
R987 AVSS.n3008 AVSS.n2991 585
R988 AVSS.n3011 AVSS.n3010 585
R989 AVSS.n3012 AVSS.n2989 585
R990 AVSS.n4474 AVSS.n4473 585
R991 AVSS.n2826 AVSS.n2807 585
R992 AVSS.n2825 AVSS.n2824 585
R993 AVSS.n2823 AVSS.n2822 585
R994 AVSS.n2821 AVSS.n2820 585
R995 AVSS.n2819 AVSS.n2818 585
R996 AVSS.n2817 AVSS.n2816 585
R997 AVSS.n2815 AVSS.n2814 585
R998 AVSS.n2813 AVSS.n2812 585
R999 AVSS.n2811 AVSS.n2810 585
R1000 AVSS.n2809 AVSS.n1721 585
R1001 AVSS.n4715 AVSS.n4714 585
R1002 AVSS.n2941 AVSS.n2940 585
R1003 AVSS.n2942 AVSS.n2913 585
R1004 AVSS.n2944 AVSS.n2943 585
R1005 AVSS.n2946 AVSS.n2912 585
R1006 AVSS.n2949 AVSS.n2948 585
R1007 AVSS.n2950 AVSS.n2911 585
R1008 AVSS.n2952 AVSS.n2951 585
R1009 AVSS.n2954 AVSS.n2910 585
R1010 AVSS.n2956 AVSS.n2955 585
R1011 AVSS.n2958 AVSS.n2957 585
R1012 AVSS.n2959 AVSS.n2908 585
R1013 AVSS.n2962 AVSS.n2961 585
R1014 AVSS.n4716 AVSS.n1717 585
R1015 AVSS.n4719 AVSS.n4718 585
R1016 AVSS.n1718 AVSS.n1716 585
R1017 AVSS.n2923 AVSS.n2920 585
R1018 AVSS.n2925 AVSS.n2924 585
R1019 AVSS.n2926 AVSS.n2919 585
R1020 AVSS.n2928 AVSS.n2927 585
R1021 AVSS.n2930 AVSS.n2917 585
R1022 AVSS.n2932 AVSS.n2931 585
R1023 AVSS.n2933 AVSS.n2916 585
R1024 AVSS.n2935 AVSS.n2934 585
R1025 AVSS.n2937 AVSS.n2915 585
R1026 AVSS.n2938 AVSS.n2914 585
R1027 AVSS.n2938 AVSS.n1719 585
R1028 AVSS.n4684 AVSS.n4683 585
R1029 AVSS.n4686 AVSS.n1734 585
R1030 AVSS.n4688 AVSS.n4687 585
R1031 AVSS.n4689 AVSS.n1733 585
R1032 AVSS.n4691 AVSS.n4690 585
R1033 AVSS.n4693 AVSS.n1731 585
R1034 AVSS.n4695 AVSS.n4694 585
R1035 AVSS.n4696 AVSS.n1730 585
R1036 AVSS.n4698 AVSS.n4697 585
R1037 AVSS.n4700 AVSS.n1728 585
R1038 AVSS.n4702 AVSS.n4701 585
R1039 AVSS.n4703 AVSS.n1727 585
R1040 AVSS.n4705 AVSS.n4704 585
R1041 AVSS.n4705 AVSS.n1719 585
R1042 AVSS.n4504 AVSS.n4503 585
R1043 AVSS.n4506 AVSS.n2787 585
R1044 AVSS.n4508 AVSS.n4507 585
R1045 AVSS.n4509 AVSS.n2786 585
R1046 AVSS.n4511 AVSS.n4510 585
R1047 AVSS.n4513 AVSS.n2784 585
R1048 AVSS.n4515 AVSS.n4514 585
R1049 AVSS.n4516 AVSS.n2783 585
R1050 AVSS.n4518 AVSS.n4517 585
R1051 AVSS.n4520 AVSS.n2781 585
R1052 AVSS.n4522 AVSS.n4521 585
R1053 AVSS.n4523 AVSS.n2780 585
R1054 AVSS.n4673 AVSS.n4672 585
R1055 AVSS.n4673 AVSS.n1719 585
R1056 AVSS.n3241 AVSS.n3240 585
R1057 AVSS.n3239 AVSS.n3238 585
R1058 AVSS.n3237 AVSS.n3086 585
R1059 AVSS.n3235 AVSS.n3234 585
R1060 AVSS.n3233 AVSS.n3087 585
R1061 AVSS.n3232 AVSS.n3231 585
R1062 AVSS.n3229 AVSS.n3088 585
R1063 AVSS.n3227 AVSS.n3226 585
R1064 AVSS.n3225 AVSS.n3089 585
R1065 AVSS.n3224 AVSS.n3223 585
R1066 AVSS.n3221 AVSS.n3090 585
R1067 AVSS.n3219 AVSS.n3218 585
R1068 AVSS.n2163 AVSS.n2161 585
R1069 AVSS.n2160 AVSS.n2159 585
R1070 AVSS.n2158 AVSS.n2157 585
R1071 AVSS.n2156 AVSS.n2155 585
R1072 AVSS.n2154 AVSS.n2153 585
R1073 AVSS.n2152 AVSS.n2151 585
R1074 AVSS.n2150 AVSS.n2149 585
R1075 AVSS.n2148 AVSS.n2147 585
R1076 AVSS.n2146 AVSS.n2145 585
R1077 AVSS.n2144 AVSS.n2143 585
R1078 AVSS.n2142 AVSS.n2141 585
R1079 AVSS.n2140 AVSS.n2139 585
R1080 AVSS.n2138 AVSS.n1139 585
R1081 AVSS.n4933 AVSS.n1139 585
R1082 AVSS.n4937 AVSS.n1089 585
R1083 AVSS.n4936 AVSS.n4935 585
R1084 AVSS.n1091 AVSS.n1090 585
R1085 AVSS.n4650 AVSS.n4649 585
R1086 AVSS.n4652 AVSS.n4651 585
R1087 AVSS.n4654 AVSS.n4653 585
R1088 AVSS.n4656 AVSS.n4655 585
R1089 AVSS.n4658 AVSS.n4657 585
R1090 AVSS.n4660 AVSS.n4659 585
R1091 AVSS.n4662 AVSS.n4661 585
R1092 AVSS.n4664 AVSS.n4663 585
R1093 AVSS.n4666 AVSS.n4665 585
R1094 AVSS.n4648 AVSS.n1126 585
R1095 AVSS.n4933 AVSS.n1126 585
R1096 AVSS.n1348 AVSS.n1347 585
R1097 AVSS.n1350 AVSS.n1349 585
R1098 AVSS.n1352 AVSS.n1351 585
R1099 AVSS.n1354 AVSS.n1353 585
R1100 AVSS.n1356 AVSS.n1355 585
R1101 AVSS.n1358 AVSS.n1357 585
R1102 AVSS.n1360 AVSS.n1359 585
R1103 AVSS.n1362 AVSS.n1361 585
R1104 AVSS.n1364 AVSS.n1363 585
R1105 AVSS.n1365 AVSS.n1146 585
R1106 AVSS.n1367 AVSS.n1366 585
R1107 AVSS.n1173 AVSS.n1145 585
R1108 AVSS.n4932 AVSS.n4931 585
R1109 AVSS.n4933 AVSS.n4932 585
R1110 AVSS.n1371 AVSS.n1369 585
R1111 AVSS.n4806 AVSS.n4805 585
R1112 AVSS.n4804 AVSS.n4803 585
R1113 AVSS.n4802 AVSS.n4801 585
R1114 AVSS.n4800 AVSS.n4799 585
R1115 AVSS.n4798 AVSS.n4797 585
R1116 AVSS.n4796 AVSS.n4795 585
R1117 AVSS.n4794 AVSS.n4793 585
R1118 AVSS.n4792 AVSS.n4791 585
R1119 AVSS.n4790 AVSS.n4789 585
R1120 AVSS.n4788 AVSS.n4787 585
R1121 AVSS.n4786 AVSS.n4785 585
R1122 AVSS.n4930 AVSS.n1370 585
R1123 AVSS.n4929 AVSS.n4928 585
R1124 AVSS.n1373 AVSS.n1372 585
R1125 AVSS.n4924 AVSS.n4923 585
R1126 AVSS.n4922 AVSS.n1378 585
R1127 AVSS.n4921 AVSS.n4920 585
R1128 AVSS.n4919 AVSS.n4918 585
R1129 AVSS.n4917 AVSS.n4916 585
R1130 AVSS.n4915 AVSS.n4914 585
R1131 AVSS.n4913 AVSS.n4912 585
R1132 AVSS.n4911 AVSS.n4910 585
R1133 AVSS.n4909 AVSS.n4908 585
R1134 AVSS.n2115 AVSS.n2114 585
R1135 AVSS.n2117 AVSS.n2088 585
R1136 AVSS.n2120 AVSS.n2119 585
R1137 AVSS.n2121 AVSS.n2087 585
R1138 AVSS.n2123 AVSS.n2122 585
R1139 AVSS.n2125 AVSS.n2086 585
R1140 AVSS.n2128 AVSS.n2127 585
R1141 AVSS.n2129 AVSS.n2085 585
R1142 AVSS.n2131 AVSS.n2130 585
R1143 AVSS.n2133 AVSS.n2084 585
R1144 AVSS.n2134 AVSS.n2082 585
R1145 AVSS.n2137 AVSS.n2136 585
R1146 AVSS.n2165 AVSS.n2164 585
R1147 AVSS.n2166 AVSS.n2080 585
R1148 AVSS.n2168 AVSS.n2167 585
R1149 AVSS.n2170 AVSS.n2078 585
R1150 AVSS.n2172 AVSS.n2171 585
R1151 AVSS.n2173 AVSS.n2077 585
R1152 AVSS.n2175 AVSS.n2174 585
R1153 AVSS.n2177 AVSS.n2075 585
R1154 AVSS.n2179 AVSS.n2178 585
R1155 AVSS.n2180 AVSS.n2074 585
R1156 AVSS.n2182 AVSS.n2181 585
R1157 AVSS.n2184 AVSS.n2072 585
R1158 AVSS.n4625 AVSS.n4624 585
R1159 AVSS.n4627 AVSS.n4623 585
R1160 AVSS.n4630 AVSS.n4629 585
R1161 AVSS.n4631 AVSS.n4622 585
R1162 AVSS.n4633 AVSS.n4632 585
R1163 AVSS.n4635 AVSS.n4621 585
R1164 AVSS.n4638 AVSS.n4637 585
R1165 AVSS.n4639 AVSS.n4620 585
R1166 AVSS.n4641 AVSS.n4640 585
R1167 AVSS.n4643 AVSS.n4619 585
R1168 AVSS.n4644 AVSS.n4617 585
R1169 AVSS.n4647 AVSS.n4646 585
R1170 AVSS.n4939 AVSS.n4938 585
R1171 AVSS.n4941 AVSS.n1087 585
R1172 AVSS.n4943 AVSS.n4942 585
R1173 AVSS.n4944 AVSS.n1086 585
R1174 AVSS.n4946 AVSS.n4945 585
R1175 AVSS.n4948 AVSS.n1084 585
R1176 AVSS.n4950 AVSS.n4949 585
R1177 AVSS.n4951 AVSS.n1083 585
R1178 AVSS.n4953 AVSS.n4952 585
R1179 AVSS.n4955 AVSS.n1080 585
R1180 AVSS.n4957 AVSS.n4956 585
R1181 AVSS.n4958 AVSS.n1079 585
R1182 AVSS.n1196 AVSS.n1165 585
R1183 AVSS.n1195 AVSS.n1194 585
R1184 AVSS.n1167 AVSS.n1166 585
R1185 AVSS.n1190 AVSS.n1189 585
R1186 AVSS.n1188 AVSS.n1172 585
R1187 AVSS.n1187 AVSS.n1186 585
R1188 AVSS.n1185 AVSS.n1184 585
R1189 AVSS.n1183 AVSS.n1182 585
R1190 AVSS.n1181 AVSS.n1180 585
R1191 AVSS.n1179 AVSS.n1178 585
R1192 AVSS.n1177 AVSS.n1176 585
R1193 AVSS.n1175 AVSS.n1174 585
R1194 AVSS.n4907 AVSS.n1379 585
R1195 AVSS.n4905 AVSS.n4904 585
R1196 AVSS.n1381 AVSS.n1380 585
R1197 AVSS.n4742 AVSS.n4741 585
R1198 AVSS.n4744 AVSS.n4743 585
R1199 AVSS.n4746 AVSS.n4738 585
R1200 AVSS.n4748 AVSS.n4747 585
R1201 AVSS.n4749 AVSS.n4737 585
R1202 AVSS.n4751 AVSS.n4750 585
R1203 AVSS.n4753 AVSS.n4735 585
R1204 AVSS.n4755 AVSS.n4754 585
R1205 AVSS.n4756 AVSS.n4734 585
R1206 AVSS.n4758 AVSS.n4757 585
R1207 AVSS.n4758 AVSS.n1071 585
R1208 AVSS.n2185 AVSS.n2070 585
R1209 AVSS.n2188 AVSS.n2187 585
R1210 AVSS.n2071 AVSS.n2069 585
R1211 AVSS.n2097 AVSS.n2096 585
R1212 AVSS.n2099 AVSS.n2098 585
R1213 AVSS.n2101 AVSS.n2093 585
R1214 AVSS.n2103 AVSS.n2102 585
R1215 AVSS.n2104 AVSS.n2092 585
R1216 AVSS.n2106 AVSS.n2105 585
R1217 AVSS.n2108 AVSS.n2091 585
R1218 AVSS.n2109 AVSS.n2090 585
R1219 AVSS.n2112 AVSS.n2111 585
R1220 AVSS.n2113 AVSS.n2089 585
R1221 AVSS.n2089 AVSS.n1071 585
R1222 AVSS.n4960 AVSS.n4959 585
R1223 AVSS.n4962 AVSS.n1077 585
R1224 AVSS.n4964 AVSS.n4963 585
R1225 AVSS.n4965 AVSS.n1076 585
R1226 AVSS.n4967 AVSS.n4966 585
R1227 AVSS.n4969 AVSS.n1074 585
R1228 AVSS.n4971 AVSS.n4970 585
R1229 AVSS.n4972 AVSS.n1073 585
R1230 AVSS.n4974 AVSS.n4973 585
R1231 AVSS.n4976 AVSS.n1072 585
R1232 AVSS.n4977 AVSS.n1069 585
R1233 AVSS.n4980 AVSS.n4979 585
R1234 AVSS.n1070 AVSS.n1068 585
R1235 AVSS.n1071 AVSS.n1070 585
R1236 AVSS.n1317 AVSS.n1316 585
R1237 AVSS.n1315 AVSS.n1314 585
R1238 AVSS.n1313 AVSS.n1160 585
R1239 AVSS.n1311 AVSS.n1310 585
R1240 AVSS.n1309 AVSS.n1161 585
R1241 AVSS.n1308 AVSS.n1307 585
R1242 AVSS.n1305 AVSS.n1162 585
R1243 AVSS.n1303 AVSS.n1302 585
R1244 AVSS.n1301 AVSS.n1163 585
R1245 AVSS.n1300 AVSS.n1299 585
R1246 AVSS.n1297 AVSS.n1164 585
R1247 AVSS.n1295 AVSS.n1294 585
R1248 AVSS.n1589 AVSS.n1588 585
R1249 AVSS.n1592 AVSS.n1591 585
R1250 AVSS.n1590 AVSS.n1383 585
R1251 AVSS.n1495 AVSS.n1494 585
R1252 AVSS.n1497 AVSS.n1496 585
R1253 AVSS.n1499 AVSS.n1498 585
R1254 AVSS.n1501 AVSS.n1500 585
R1255 AVSS.n1503 AVSS.n1502 585
R1256 AVSS.n1505 AVSS.n1504 585
R1257 AVSS.n1507 AVSS.n1506 585
R1258 AVSS.n1509 AVSS.n1508 585
R1259 AVSS.n1511 AVSS.n1510 585
R1260 AVSS.n1512 AVSS.n661 585
R1261 AVSS.n4988 AVSS.n661 585
R1262 AVSS.n4992 AVSS.n644 585
R1263 AVSS.n4991 AVSS.n4990 585
R1264 AVSS.n945 AVSS.n647 585
R1265 AVSS.n947 AVSS.n946 585
R1266 AVSS.n949 AVSS.n948 585
R1267 AVSS.n951 AVSS.n950 585
R1268 AVSS.n953 AVSS.n952 585
R1269 AVSS.n955 AVSS.n954 585
R1270 AVSS.n957 AVSS.n956 585
R1271 AVSS.n959 AVSS.n958 585
R1272 AVSS.n961 AVSS.n960 585
R1273 AVSS.n962 AVSS.n893 585
R1274 AVSS.n964 AVSS.n963 585
R1275 AVSS.n4988 AVSS.n964 585
R1276 AVSS.n2411 AVSS.n2304 585
R1277 AVSS.n2317 AVSS.n2316 585
R1278 AVSS.n2319 AVSS.n2318 585
R1279 AVSS.n2321 AVSS.n2320 585
R1280 AVSS.n2323 AVSS.n2322 585
R1281 AVSS.n2325 AVSS.n2324 585
R1282 AVSS.n2327 AVSS.n2326 585
R1283 AVSS.n2329 AVSS.n2328 585
R1284 AVSS.n2331 AVSS.n2330 585
R1285 AVSS.n2333 AVSS.n2332 585
R1286 AVSS.n2335 AVSS.n2334 585
R1287 AVSS.n2337 AVSS.n2336 585
R1288 AVSS.n2338 AVSS.n654 585
R1289 AVSS.n4988 AVSS.n654 585
R1290 AVSS.n2231 AVSS.n2229 585
R1291 AVSS.n2228 AVSS.n2227 585
R1292 AVSS.n2226 AVSS.n2225 585
R1293 AVSS.n2224 AVSS.n2223 585
R1294 AVSS.n2222 AVSS.n2221 585
R1295 AVSS.n2220 AVSS.n2219 585
R1296 AVSS.n2218 AVSS.n2217 585
R1297 AVSS.n2216 AVSS.n2215 585
R1298 AVSS.n2214 AVSS.n2213 585
R1299 AVSS.n2212 AVSS.n2211 585
R1300 AVSS.n2210 AVSS.n2209 585
R1301 AVSS.n974 AVSS.n972 585
R1302 AVSS.n4987 AVSS.n4986 585
R1303 AVSS.n4988 AVSS.n4987 585
R1304 AVSS.n671 AVSS.n669 585
R1305 AVSS.n718 AVSS.n717 585
R1306 AVSS.n720 AVSS.n719 585
R1307 AVSS.n722 AVSS.n721 585
R1308 AVSS.n724 AVSS.n723 585
R1309 AVSS.n726 AVSS.n725 585
R1310 AVSS.n728 AVSS.n727 585
R1311 AVSS.n730 AVSS.n729 585
R1312 AVSS.n732 AVSS.n731 585
R1313 AVSS.n734 AVSS.n733 585
R1314 AVSS.n736 AVSS.n735 585
R1315 AVSS.n716 AVSS.n715 585
R1316 AVSS.n1862 AVSS.n1860 585
R1317 AVSS.n1860 AVSS.n1071 585
R1318 AVSS.n1864 AVSS.n1863 585
R1319 AVSS.n1866 AVSS.n1858 585
R1320 AVSS.n1869 AVSS.n1868 585
R1321 AVSS.n1870 AVSS.n1857 585
R1322 AVSS.n1872 AVSS.n1871 585
R1323 AVSS.n1874 AVSS.n1856 585
R1324 AVSS.n1877 AVSS.n1876 585
R1325 AVSS.n1878 AVSS.n1855 585
R1326 AVSS.n1880 AVSS.n1879 585
R1327 AVSS.n1882 AVSS.n1854 585
R1328 AVSS.n1885 AVSS.n1884 585
R1329 AVSS.n2512 AVSS.n1853 585
R1330 AVSS.n2585 AVSS.n2584 585
R1331 AVSS.n2578 AVSS.n1741 585
R1332 AVSS.n2580 AVSS.n2579 585
R1333 AVSS.n2577 AVSS.n1746 585
R1334 AVSS.n2576 AVSS.n2575 585
R1335 AVSS.n2574 AVSS.n2573 585
R1336 AVSS.n2572 AVSS.n2571 585
R1337 AVSS.n2570 AVSS.n2569 585
R1338 AVSS.n2568 AVSS.n2567 585
R1339 AVSS.n2566 AVSS.n2565 585
R1340 AVSS.n2564 AVSS.n2563 585
R1341 AVSS.n1859 AVSS.n1747 585
R1342 AVSS.n2586 AVSS.n1119 585
R1343 AVSS.n4933 AVSS.n1119 585
R1344 AVSS.n2588 AVSS.n2587 585
R1345 AVSS.n1825 AVSS.n1739 585
R1346 AVSS.n1827 AVSS.n1826 585
R1347 AVSS.n1829 AVSS.n1828 585
R1348 AVSS.n1831 AVSS.n1830 585
R1349 AVSS.n1833 AVSS.n1832 585
R1350 AVSS.n1835 AVSS.n1834 585
R1351 AVSS.n1837 AVSS.n1836 585
R1352 AVSS.n1839 AVSS.n1838 585
R1353 AVSS.n1841 AVSS.n1840 585
R1354 AVSS.n1843 AVSS.n1842 585
R1355 AVSS.n1846 AVSS.n1845 585
R1356 AVSS.n2515 AVSS.n2514 585
R1357 AVSS.n2517 AVSS.n1852 585
R1358 AVSS.n2520 AVSS.n2519 585
R1359 AVSS.n2521 AVSS.n1851 585
R1360 AVSS.n2523 AVSS.n2522 585
R1361 AVSS.n2525 AVSS.n1850 585
R1362 AVSS.n2528 AVSS.n2527 585
R1363 AVSS.n2529 AVSS.n1849 585
R1364 AVSS.n2531 AVSS.n2530 585
R1365 AVSS.n2533 AVSS.n1848 585
R1366 AVSS.n2534 AVSS.n1824 585
R1367 AVSS.n2537 AVSS.n2536 585
R1368 AVSS.n3968 AVSS.n3967 585
R1369 AVSS.n3970 AVSS.n3906 585
R1370 AVSS.n3973 AVSS.n3972 585
R1371 AVSS.n3974 AVSS.n3905 585
R1372 AVSS.n3976 AVSS.n3975 585
R1373 AVSS.n3978 AVSS.n3904 585
R1374 AVSS.n3981 AVSS.n3980 585
R1375 AVSS.n3982 AVSS.n3903 585
R1376 AVSS.n3984 AVSS.n3983 585
R1377 AVSS.n3986 AVSS.n3902 585
R1378 AVSS.n3989 AVSS.n3988 585
R1379 AVSS.n4269 AVSS.n3901 585
R1380 AVSS.n4293 AVSS.n3889 585
R1381 AVSS.n4296 AVSS.n4295 585
R1382 AVSS.n3891 AVSS.n3890 585
R1383 AVSS.n3925 AVSS.n3924 585
R1384 AVSS.n3927 AVSS.n3926 585
R1385 AVSS.n3929 AVSS.n3922 585
R1386 AVSS.n3932 AVSS.n3931 585
R1387 AVSS.n3933 AVSS.n3921 585
R1388 AVSS.n3935 AVSS.n3934 585
R1389 AVSS.n3937 AVSS.n3920 585
R1390 AVSS.n3938 AVSS.n3919 585
R1391 AVSS.n3941 AVSS.n3940 585
R1392 AVSS.n3757 AVSS.n3756 585
R1393 AVSS.n3759 AVSS.n3695 585
R1394 AVSS.n3762 AVSS.n3761 585
R1395 AVSS.n3763 AVSS.n3694 585
R1396 AVSS.n3765 AVSS.n3764 585
R1397 AVSS.n3767 AVSS.n3693 585
R1398 AVSS.n3770 AVSS.n3769 585
R1399 AVSS.n3771 AVSS.n3692 585
R1400 AVSS.n3773 AVSS.n3772 585
R1401 AVSS.n3775 AVSS.n3691 585
R1402 AVSS.n3778 AVSS.n3777 585
R1403 AVSS.n4302 AVSS.n3690 585
R1404 AVSS.n4326 AVSS.n3678 585
R1405 AVSS.n4329 AVSS.n4328 585
R1406 AVSS.n3680 AVSS.n3679 585
R1407 AVSS.n3714 AVSS.n3713 585
R1408 AVSS.n3716 AVSS.n3715 585
R1409 AVSS.n3718 AVSS.n3711 585
R1410 AVSS.n3721 AVSS.n3720 585
R1411 AVSS.n3722 AVSS.n3710 585
R1412 AVSS.n3724 AVSS.n3723 585
R1413 AVSS.n3726 AVSS.n3709 585
R1414 AVSS.n3727 AVSS.n3708 585
R1415 AVSS.n3730 AVSS.n3729 585
R1416 AVSS.n3620 AVSS.n3619 585
R1417 AVSS.n3622 AVSS.n3519 585
R1418 AVSS.n3625 AVSS.n3624 585
R1419 AVSS.n3626 AVSS.n3518 585
R1420 AVSS.n3628 AVSS.n3627 585
R1421 AVSS.n3630 AVSS.n3517 585
R1422 AVSS.n3633 AVSS.n3632 585
R1423 AVSS.n3634 AVSS.n3516 585
R1424 AVSS.n3636 AVSS.n3635 585
R1425 AVSS.n3638 AVSS.n3515 585
R1426 AVSS.n3640 AVSS.n3639 585
R1427 AVSS.n4336 AVSS.n4335 585
R1428 AVSS.n4337 AVSS.n3512 585
R1429 AVSS.n4340 AVSS.n4339 585
R1430 AVSS.n3513 AVSS.n3511 585
R1431 AVSS.n3545 AVSS.n3542 585
R1432 AVSS.n3547 AVSS.n3546 585
R1433 AVSS.n3548 AVSS.n3541 585
R1434 AVSS.n3550 AVSS.n3549 585
R1435 AVSS.n3552 AVSS.n3539 585
R1436 AVSS.n3554 AVSS.n3553 585
R1437 AVSS.n3555 AVSS.n3538 585
R1438 AVSS.n3557 AVSS.n3556 585
R1439 AVSS.n3559 AVSS.n3537 585
R1440 AVSS.n3560 AVSS.n3536 585
R1441 AVSS.n3560 AVSS.n151 585
R1442 AVSS.n4304 AVSS.n4303 585
R1443 AVSS.n4306 AVSS.n3688 585
R1444 AVSS.n4308 AVSS.n4307 585
R1445 AVSS.n4309 AVSS.n3687 585
R1446 AVSS.n4311 AVSS.n4310 585
R1447 AVSS.n4313 AVSS.n3685 585
R1448 AVSS.n4315 AVSS.n4314 585
R1449 AVSS.n4316 AVSS.n3684 585
R1450 AVSS.n4318 AVSS.n4317 585
R1451 AVSS.n4320 AVSS.n3682 585
R1452 AVSS.n4322 AVSS.n4321 585
R1453 AVSS.n4323 AVSS.n3681 585
R1454 AVSS.n4325 AVSS.n4324 585
R1455 AVSS.n4325 AVSS.n151 585
R1456 AVSS.n4271 AVSS.n4270 585
R1457 AVSS.n4273 AVSS.n3899 585
R1458 AVSS.n4275 AVSS.n4274 585
R1459 AVSS.n4276 AVSS.n3898 585
R1460 AVSS.n4278 AVSS.n4277 585
R1461 AVSS.n4280 AVSS.n3896 585
R1462 AVSS.n4282 AVSS.n4281 585
R1463 AVSS.n4283 AVSS.n3895 585
R1464 AVSS.n4285 AVSS.n4284 585
R1465 AVSS.n4287 AVSS.n3893 585
R1466 AVSS.n4289 AVSS.n4288 585
R1467 AVSS.n4290 AVSS.n3892 585
R1468 AVSS.n4292 AVSS.n4291 585
R1469 AVSS.n4292 AVSS.n151 585
R1470 AVSS.n6191 AVSS.n6190 585
R1471 AVSS.n6193 AVSS.n156 585
R1472 AVSS.n6195 AVSS.n6194 585
R1473 AVSS.n6196 AVSS.n155 585
R1474 AVSS.n6198 AVSS.n6197 585
R1475 AVSS.n6200 AVSS.n153 585
R1476 AVSS.n6202 AVSS.n6201 585
R1477 AVSS.n6203 AVSS.n152 585
R1478 AVSS.n6205 AVSS.n6204 585
R1479 AVSS.n6207 AVSS.n149 585
R1480 AVSS.n6209 AVSS.n6208 585
R1481 AVSS.n256 AVSS.n148 585
R1482 AVSS.n4472 AVSS.n2808 585
R1483 AVSS.n4471 AVSS.n4470 585
R1484 AVSS.n2828 AVSS.n2827 585
R1485 AVSS.n2980 AVSS.n2979 585
R1486 AVSS.n2978 AVSS.n2907 585
R1487 AVSS.n2977 AVSS.n2976 585
R1488 AVSS.n2975 AVSS.n2974 585
R1489 AVSS.n2973 AVSS.n2972 585
R1490 AVSS.n2971 AVSS.n2970 585
R1491 AVSS.n2969 AVSS.n2968 585
R1492 AVSS.n2967 AVSS.n2966 585
R1493 AVSS.n2965 AVSS.n2964 585
R1494 AVSS.n2963 AVSS.n2902 585
R1495 AVSS.n4468 AVSS.n2902 585
R1496 AVSS.n3041 AVSS.n3040 585
R1497 AVSS.n3043 AVSS.n3042 585
R1498 AVSS.n3045 AVSS.n3044 585
R1499 AVSS.n3047 AVSS.n3046 585
R1500 AVSS.n3049 AVSS.n3048 585
R1501 AVSS.n3051 AVSS.n3050 585
R1502 AVSS.n3053 AVSS.n3052 585
R1503 AVSS.n3055 AVSS.n3054 585
R1504 AVSS.n3057 AVSS.n3056 585
R1505 AVSS.n3059 AVSS.n3058 585
R1506 AVSS.n3061 AVSS.n3060 585
R1507 AVSS.n3062 AVSS.n2990 585
R1508 AVSS.n3064 AVSS.n3063 585
R1509 AVSS.n4468 AVSS.n3064 585
R1510 AVSS.n2900 AVSS.n2899 585
R1511 AVSS.n2881 AVSS.n2835 585
R1512 AVSS.n2880 AVSS.n2879 585
R1513 AVSS.n2878 AVSS.n2877 585
R1514 AVSS.n2876 AVSS.n2875 585
R1515 AVSS.n2874 AVSS.n2873 585
R1516 AVSS.n2872 AVSS.n2871 585
R1517 AVSS.n2870 AVSS.n2869 585
R1518 AVSS.n2868 AVSS.n2867 585
R1519 AVSS.n2866 AVSS.n2865 585
R1520 AVSS.n2864 AVSS.n2863 585
R1521 AVSS.n2862 AVSS.n2861 585
R1522 AVSS.n2860 AVSS.n2829 585
R1523 AVSS.n4468 AVSS.n2829 585
R1524 AVSS.n3273 AVSS.n3272 585
R1525 AVSS.n3275 AVSS.n3274 585
R1526 AVSS.n3277 AVSS.n3276 585
R1527 AVSS.n3279 AVSS.n3278 585
R1528 AVSS.n3281 AVSS.n3280 585
R1529 AVSS.n3283 AVSS.n3282 585
R1530 AVSS.n3285 AVSS.n3284 585
R1531 AVSS.n3287 AVSS.n3286 585
R1532 AVSS.n3289 AVSS.n3288 585
R1533 AVSS.n3290 AVSS.n3071 585
R1534 AVSS.n3292 AVSS.n3291 585
R1535 AVSS.n3097 AVSS.n3070 585
R1536 AVSS.n230 AVSS.n229 585
R1537 AVSS.n229 AVSS.n151 585
R1538 AVSS.n4237 AVSS.n4236 585
R1539 AVSS.n4239 AVSS.n4235 585
R1540 AVSS.n4242 AVSS.n4241 585
R1541 AVSS.n4243 AVSS.n4234 585
R1542 AVSS.n4245 AVSS.n4244 585
R1543 AVSS.n4247 AVSS.n4233 585
R1544 AVSS.n4250 AVSS.n4249 585
R1545 AVSS.n4251 AVSS.n4232 585
R1546 AVSS.n4253 AVSS.n4252 585
R1547 AVSS.n4255 AVSS.n4231 585
R1548 AVSS.n4257 AVSS.n4256 585
R1549 AVSS.n4259 AVSS.n4258 585
R1550 AVSS.n4260 AVSS.n4206 585
R1551 AVSS.n4263 AVSS.n4262 585
R1552 AVSS.n4229 AVSS.n4207 585
R1553 AVSS.n4227 AVSS.n4226 585
R1554 AVSS.n4225 AVSS.n4208 585
R1555 AVSS.n4224 AVSS.n4223 585
R1556 AVSS.n4221 AVSS.n4209 585
R1557 AVSS.n4219 AVSS.n4218 585
R1558 AVSS.n4217 AVSS.n4210 585
R1559 AVSS.n4216 AVSS.n4215 585
R1560 AVSS.n4213 AVSS.n4211 585
R1561 AVSS.n213 AVSS.n211 585
R1562 AVSS.n6110 AVSS.n223 585
R1563 AVSS.n6109 AVSS.n6108 585
R1564 AVSS.n6106 AVSS.n224 585
R1565 AVSS.n6104 AVSS.n6103 585
R1566 AVSS.n6102 AVSS.n225 585
R1567 AVSS.n6101 AVSS.n6100 585
R1568 AVSS.n6098 AVSS.n226 585
R1569 AVSS.n6096 AVSS.n6095 585
R1570 AVSS.n6094 AVSS.n227 585
R1571 AVSS.n6093 AVSS.n6092 585
R1572 AVSS.n6090 AVSS.n228 585
R1573 AVSS.n6088 AVSS.n6087 585
R1574 AVSS.n257 AVSS.n232 585
R1575 AVSS.n260 AVSS.n259 585
R1576 AVSS.n255 AVSS.n233 585
R1577 AVSS.n253 AVSS.n252 585
R1578 AVSS.n251 AVSS.n234 585
R1579 AVSS.n250 AVSS.n249 585
R1580 AVSS.n247 AVSS.n235 585
R1581 AVSS.n245 AVSS.n244 585
R1582 AVSS.n243 AVSS.n236 585
R1583 AVSS.n242 AVSS.n241 585
R1584 AVSS.n239 AVSS.n237 585
R1585 AVSS.n186 AVSS.n185 585
R1586 AVSS.n3618 AVSS.n3520 585
R1587 AVSS.n3520 AVSS.n205 585
R1588 AVSS.n3617 AVSS.n3616 585
R1589 AVSS.n3616 AVSS.n3615 585
R1590 AVSS.n3522 AVSS.n3521 585
R1591 AVSS.n3614 AVSS.n3522 585
R1592 AVSS.n3612 AVSS.n3611 585
R1593 AVSS.n3613 AVSS.n3612 585
R1594 AVSS.n3610 AVSS.n3524 585
R1595 AVSS.n3524 AVSS.n3523 585
R1596 AVSS.n3609 AVSS.n3608 585
R1597 AVSS.n3608 AVSS.n3607 585
R1598 AVSS.n3526 AVSS.n3525 585
R1599 AVSS.n3606 AVSS.n3526 585
R1600 AVSS.n3582 AVSS.n3581 585
R1601 AVSS.n3582 AVSS.n3527 585
R1602 AVSS.n3585 AVSS.n3584 585
R1603 AVSS.n3584 AVSS.n3583 585
R1604 AVSS.n3586 AVSS.n3580 585
R1605 AVSS.n3580 AVSS.n3579 585
R1606 AVSS.n3588 AVSS.n3587 585
R1607 AVSS.n3589 AVSS.n3588 585
R1608 AVSS.n3578 AVSS.n3577 585
R1609 AVSS.n3590 AVSS.n3578 585
R1610 AVSS.n3593 AVSS.n3592 585
R1611 AVSS.n3592 AVSS.n3591 585
R1612 AVSS.n3755 AVSS.n3696 585
R1613 AVSS.n3696 AVSS.n199 585
R1614 AVSS.n3754 AVSS.n3753 585
R1615 AVSS.n3753 AVSS.n3752 585
R1616 AVSS.n3698 AVSS.n3697 585
R1617 AVSS.n3751 AVSS.n3698 585
R1618 AVSS.n3749 AVSS.n3748 585
R1619 AVSS.n3750 AVSS.n3749 585
R1620 AVSS.n3747 AVSS.n3700 585
R1621 AVSS.n3700 AVSS.n3699 585
R1622 AVSS.n3746 AVSS.n3745 585
R1623 AVSS.n3745 AVSS.n3744 585
R1624 AVSS.n3702 AVSS.n3701 585
R1625 AVSS.n3743 AVSS.n3702 585
R1626 AVSS.n3741 AVSS.n3740 585
R1627 AVSS.n3742 AVSS.n3741 585
R1628 AVSS.n3739 AVSS.n3704 585
R1629 AVSS.n3704 AVSS.n3703 585
R1630 AVSS.n3738 AVSS.n3737 585
R1631 AVSS.n3737 AVSS.n3736 585
R1632 AVSS.n3706 AVSS.n3705 585
R1633 AVSS.n3735 AVSS.n3706 585
R1634 AVSS.n3733 AVSS.n3732 585
R1635 AVSS.n3734 AVSS.n3733 585
R1636 AVSS.n3731 AVSS.n3707 585
R1637 AVSS.n3707 AVSS.n206 585
R1638 AVSS.n3966 AVSS.n3907 585
R1639 AVSS.n3907 AVSS.n209 585
R1640 AVSS.n3965 AVSS.n3964 585
R1641 AVSS.n3964 AVSS.n3963 585
R1642 AVSS.n3909 AVSS.n3908 585
R1643 AVSS.n3962 AVSS.n3909 585
R1644 AVSS.n3960 AVSS.n3959 585
R1645 AVSS.n3961 AVSS.n3960 585
R1646 AVSS.n3958 AVSS.n3911 585
R1647 AVSS.n3911 AVSS.n3910 585
R1648 AVSS.n3957 AVSS.n3956 585
R1649 AVSS.n3956 AVSS.n3955 585
R1650 AVSS.n3913 AVSS.n3912 585
R1651 AVSS.n3954 AVSS.n3913 585
R1652 AVSS.n3952 AVSS.n3951 585
R1653 AVSS.n3953 AVSS.n3952 585
R1654 AVSS.n3950 AVSS.n3915 585
R1655 AVSS.n3915 AVSS.n3914 585
R1656 AVSS.n3949 AVSS.n3948 585
R1657 AVSS.n3948 AVSS.n3947 585
R1658 AVSS.n3917 AVSS.n3916 585
R1659 AVSS.n3946 AVSS.n3917 585
R1660 AVSS.n3944 AVSS.n3943 585
R1661 AVSS.n3945 AVSS.n3944 585
R1662 AVSS.n3942 AVSS.n3918 585
R1663 AVSS.n3918 AVSS.n198 585
R1664 AVSS.n6112 AVSS.n6111 585
R1665 AVSS.n6112 AVSS.n202 585
R1666 AVSS.n6113 AVSS.n222 585
R1667 AVSS.n6114 AVSS.n6113 585
R1668 AVSS.n6117 AVSS.n6116 585
R1669 AVSS.n6116 AVSS.n6115 585
R1670 AVSS.n6118 AVSS.n221 585
R1671 AVSS.n221 AVSS.n220 585
R1672 AVSS.n6120 AVSS.n6119 585
R1673 AVSS.n6121 AVSS.n6120 585
R1674 AVSS.n219 AVSS.n218 585
R1675 AVSS.n6122 AVSS.n219 585
R1676 AVSS.n6125 AVSS.n6124 585
R1677 AVSS.n6124 AVSS.n6123 585
R1678 AVSS.n6126 AVSS.n217 585
R1679 AVSS.n217 AVSS.n216 585
R1680 AVSS.n6128 AVSS.n6127 585
R1681 AVSS.n6129 AVSS.n6128 585
R1682 AVSS.n215 AVSS.n214 585
R1683 AVSS.n6130 AVSS.n215 585
R1684 AVSS.n6133 AVSS.n6132 585
R1685 AVSS.n6132 AVSS.n6131 585
R1686 AVSS.n6134 AVSS.n212 585
R1687 AVSS.n212 AVSS.n210 585
R1688 AVSS.n6136 AVSS.n6135 585
R1689 AVSS.n6137 AVSS.n6136 585
R1690 AVSS.n176 AVSS.n175 585
R1691 AVSS.n6161 AVSS.n176 585
R1692 AVSS.n6159 AVSS.n6158 585
R1693 AVSS.n6160 AVSS.n6159 585
R1694 AVSS.n6157 AVSS.n178 585
R1695 AVSS.n178 AVSS.n177 585
R1696 AVSS.n6156 AVSS.n6155 585
R1697 AVSS.n6155 AVSS.n6154 585
R1698 AVSS.n6152 AVSS.n179 585
R1699 AVSS.n6153 AVSS.n6152 585
R1700 AVSS.n6151 AVSS.n6150 585
R1701 AVSS.n6151 AVSS.n168 585
R1702 AVSS.n6149 AVSS.n180 585
R1703 AVSS.n180 AVSS.n167 585
R1704 AVSS.n6148 AVSS.n6147 585
R1705 AVSS.n6147 AVSS.n6146 585
R1706 AVSS.n182 AVSS.n181 585
R1707 AVSS.n6145 AVSS.n182 585
R1708 AVSS.n6143 AVSS.n6142 585
R1709 AVSS.n6144 AVSS.n6143 585
R1710 AVSS.n6141 AVSS.n184 585
R1711 AVSS.n184 AVSS.n183 585
R1712 AVSS.n6140 AVSS.n6139 585
R1713 AVSS.n6139 AVSS.n6138 585
R1714 AVSS.n6189 AVSS.n158 585
R1715 AVSS.n161 AVSS.n158 585
R1716 AVSS.n6165 AVSS.n174 585
R1717 AVSS.n174 AVSS.n173 585
R1718 AVSS.n6167 AVSS.n6166 585
R1719 AVSS.n6168 AVSS.n6167 585
R1720 AVSS.n172 AVSS.n171 585
R1721 AVSS.n6169 AVSS.n172 585
R1722 AVSS.n6172 AVSS.n6171 585
R1723 AVSS.n6171 AVSS.n6170 585
R1724 AVSS.n6173 AVSS.n170 585
R1725 AVSS.n170 AVSS.n169 585
R1726 AVSS.n6175 AVSS.n6174 585
R1727 AVSS.n6176 AVSS.n6175 585
R1728 AVSS.n165 AVSS.n164 585
R1729 AVSS.n6177 AVSS.n165 585
R1730 AVSS.n6180 AVSS.n6179 585
R1731 AVSS.n6179 AVSS.n6178 585
R1732 AVSS.n6181 AVSS.n163 585
R1733 AVSS.n163 AVSS.n162 585
R1734 AVSS.n6183 AVSS.n6182 585
R1735 AVSS.n6184 AVSS.n6183 585
R1736 AVSS.n160 AVSS.n159 585
R1737 AVSS.n6185 AVSS.n160 585
R1738 AVSS.n6188 AVSS.n6187 585
R1739 AVSS.n6187 AVSS.n6186 585
R1740 AVSS.n6164 AVSS.n6163 585
R1741 AVSS.n6163 AVSS.n6162 585
R1742 AVSS.n3242 AVSS.n3084 585
R1743 AVSS.n3243 AVSS.n3242 585
R1744 AVSS.n3265 AVSS.n3074 585
R1745 AVSS.n3269 AVSS.n3074 585
R1746 AVSS.n3267 AVSS.n3266 585
R1747 AVSS.n3268 AVSS.n3267 585
R1748 AVSS.n3264 AVSS.n3076 585
R1749 AVSS.n3076 AVSS.n3075 585
R1750 AVSS.n3263 AVSS.n3262 585
R1751 AVSS.n3262 AVSS.n3261 585
R1752 AVSS.n3078 AVSS.n3077 585
R1753 AVSS.n3260 AVSS.n3078 585
R1754 AVSS.n3258 AVSS.n3257 585
R1755 AVSS.n3259 AVSS.n3258 585
R1756 AVSS.n3256 AVSS.n3079 585
R1757 AVSS.n3252 AVSS.n3079 585
R1758 AVSS.n3255 AVSS.n3254 585
R1759 AVSS.n3254 AVSS.n3253 585
R1760 AVSS.n3081 AVSS.n3080 585
R1761 AVSS.n3251 AVSS.n3081 585
R1762 AVSS.n3249 AVSS.n3248 585
R1763 AVSS.n3250 AVSS.n3249 585
R1764 AVSS.n3247 AVSS.n3083 585
R1765 AVSS.n3083 AVSS.n3082 585
R1766 AVSS.n3246 AVSS.n3245 585
R1767 AVSS.n3245 AVSS.n3244 585
R1768 AVSS.n3271 AVSS.n3073 585
R1769 AVSS.n3271 AVSS.n3270 585
R1770 AVSS.n1318 AVSS.n1158 585
R1771 AVSS.n1319 AVSS.n1318 585
R1772 AVSS.n1340 AVSS.n1149 585
R1773 AVSS.n1344 AVSS.n1149 585
R1774 AVSS.n1342 AVSS.n1341 585
R1775 AVSS.n1343 AVSS.n1342 585
R1776 AVSS.n1339 AVSS.n1151 585
R1777 AVSS.n1151 AVSS.n1150 585
R1778 AVSS.n1338 AVSS.n1337 585
R1779 AVSS.n1337 AVSS.n1336 585
R1780 AVSS.n1335 AVSS.n1152 585
R1781 AVSS.n1335 AVSS.n297 585
R1782 AVSS.n1334 AVSS.n1333 585
R1783 AVSS.n1334 AVSS.n296 585
R1784 AVSS.n1332 AVSS.n1153 585
R1785 AVSS.n1328 AVSS.n1153 585
R1786 AVSS.n1331 AVSS.n1330 585
R1787 AVSS.n1330 AVSS.n1329 585
R1788 AVSS.n1155 AVSS.n1154 585
R1789 AVSS.n1327 AVSS.n1155 585
R1790 AVSS.n1325 AVSS.n1324 585
R1791 AVSS.n1326 AVSS.n1325 585
R1792 AVSS.n1323 AVSS.n1157 585
R1793 AVSS.n1157 AVSS.n1156 585
R1794 AVSS.n1322 AVSS.n1321 585
R1795 AVSS.n1321 AVSS.n1320 585
R1796 AVSS.n1346 AVSS.n1148 585
R1797 AVSS.n1346 AVSS.n1345 585
R1798 AVSS.n857 AVSS.n856 585
R1799 AVSS.n858 AVSS.n857 585
R1800 AVSS.n882 AVSS.n670 585
R1801 AVSS.n670 AVSS.n668 585
R1802 AVSS.n881 AVSS.n880 585
R1803 AVSS.n880 AVSS.n879 585
R1804 AVSS.n673 AVSS.n672 585
R1805 AVSS.n878 AVSS.n673 585
R1806 AVSS.n876 AVSS.n875 585
R1807 AVSS.n877 AVSS.n876 585
R1808 AVSS.n874 AVSS.n675 585
R1809 AVSS.n675 AVSS.n674 585
R1810 AVSS.n873 AVSS.n872 585
R1811 AVSS.n872 AVSS.n871 585
R1812 AVSS.n870 AVSS.n676 585
R1813 AVSS.n870 AVSS.n869 585
R1814 AVSS.n864 AVSS.n677 585
R1815 AVSS.n868 AVSS.n677 585
R1816 AVSS.n866 AVSS.n865 585
R1817 AVSS.n867 AVSS.n866 585
R1818 AVSS.n863 AVSS.n679 585
R1819 AVSS.n679 AVSS.n678 585
R1820 AVSS.n862 AVSS.n861 585
R1821 AVSS.n861 AVSS.n860 585
R1822 AVSS.n681 AVSS.n680 585
R1823 AVSS.n859 AVSS.n681 585
R1824 AVSS.n884 AVSS.n883 585
R1825 AVSS.n885 AVSS.n884 585
R1826 AVSS.n5642 AVSS.n5641 585
R1827 AVSS.n5674 AVSS.n5642 585
R1828 AVSS.n5696 AVSS.n5631 585
R1829 AVSS.n5700 AVSS.n5631 585
R1830 AVSS.n5698 AVSS.n5697 585
R1831 AVSS.n5699 AVSS.n5698 585
R1832 AVSS.n5695 AVSS.n5633 585
R1833 AVSS.n5633 AVSS.n5632 585
R1834 AVSS.n5694 AVSS.n5693 585
R1835 AVSS.n5693 AVSS.n5692 585
R1836 AVSS.n5635 AVSS.n5634 585
R1837 AVSS.n5691 AVSS.n5635 585
R1838 AVSS.n5689 AVSS.n5688 585
R1839 AVSS.n5690 AVSS.n5689 585
R1840 AVSS.n5687 AVSS.n5636 585
R1841 AVSS.n5683 AVSS.n5636 585
R1842 AVSS.n5686 AVSS.n5685 585
R1843 AVSS.n5685 AVSS.n5684 585
R1844 AVSS.n5638 AVSS.n5637 585
R1845 AVSS.n5682 AVSS.n5638 585
R1846 AVSS.n5680 AVSS.n5679 585
R1847 AVSS.n5681 AVSS.n5680 585
R1848 AVSS.n5678 AVSS.n5640 585
R1849 AVSS.n5640 AVSS.n5639 585
R1850 AVSS.n5677 AVSS.n5676 585
R1851 AVSS.n5676 AVSS.n5675 585
R1852 AVSS.n5702 AVSS.n5630 585
R1853 AVSS.n5702 AVSS.n5701 585
R1854 AVSS.n5913 AVSS.n5912 585
R1855 AVSS.n5914 AVSS.n306 585
R1856 AVSS.n306 AVSS.n305 585
R1857 AVSS.n5916 AVSS.n5915 585
R1858 AVSS.n5917 AVSS.n5916 585
R1859 AVSS.n304 AVSS.n303 585
R1860 AVSS.n5918 AVSS.n304 585
R1861 AVSS.n5921 AVSS.n5920 585
R1862 AVSS.n5920 AVSS.n5919 585
R1863 AVSS.n5922 AVSS.n301 585
R1864 AVSS.n301 AVSS.n299 585
R1865 AVSS.n5924 AVSS.n5923 585
R1866 AVSS.n5925 AVSS.n5924 585
R1867 AVSS.n3563 AVSS.n3562 585
R1868 AVSS.n3562 AVSS.n3561 585
R1869 AVSS.n3564 AVSS.n3535 585
R1870 AVSS.n3535 AVSS.n3534 585
R1871 AVSS.n3566 AVSS.n3565 585
R1872 AVSS.n3567 AVSS.n3566 585
R1873 AVSS.n3533 AVSS.n3532 585
R1874 AVSS.n3568 AVSS.n3533 585
R1875 AVSS.n3571 AVSS.n3570 585
R1876 AVSS.n3570 AVSS.n3569 585
R1877 AVSS.n3572 AVSS.n3530 585
R1878 AVSS.n3530 AVSS.n3528 585
R1879 AVSS.n3604 AVSS.n3603 585
R1880 AVSS.n3605 AVSS.n3604 585
R1881 AVSS.n3602 AVSS.n3531 585
R1882 AVSS.n3531 AVSS.n3529 585
R1883 AVSS.n3601 AVSS.n3600 585
R1884 AVSS.n3600 AVSS.n3599 585
R1885 AVSS.n3574 AVSS.n3573 585
R1886 AVSS.n3598 AVSS.n3574 585
R1887 AVSS.n3596 AVSS.n3595 585
R1888 AVSS.n3597 AVSS.n3596 585
R1889 AVSS.n3594 AVSS.n3576 585
R1890 AVSS.n3576 AVSS.n3575 585
R1891 AVSS.n4759 AVSS.n4733 585
R1892 AVSS.n4760 AVSS.n4759 585
R1893 AVSS.n4763 AVSS.n4762 585
R1894 AVSS.n4762 AVSS.n4761 585
R1895 AVSS.n4764 AVSS.n4732 585
R1896 AVSS.n4732 AVSS.n4731 585
R1897 AVSS.n4767 AVSS.n4766 585
R1898 AVSS.n4768 AVSS.n4767 585
R1899 AVSS.n4765 AVSS.n4729 585
R1900 AVSS.n4769 AVSS.n4729 585
R1901 AVSS.n4771 AVSS.n4730 585
R1902 AVSS.n4771 AVSS.n4770 585
R1903 AVSS.n4772 AVSS.n4728 585
R1904 AVSS.n4773 AVSS.n4772 585
R1905 AVSS.n4776 AVSS.n4775 585
R1906 AVSS.n4775 AVSS.n4774 585
R1907 AVSS.n4777 AVSS.n4727 585
R1908 AVSS.n4727 AVSS.n4726 585
R1909 AVSS.n4780 AVSS.n4779 585
R1910 AVSS.n4781 AVSS.n4780 585
R1911 AVSS.n4778 AVSS.n4725 585
R1912 AVSS.n4782 AVSS.n4725 585
R1913 AVSS.n4784 AVSS.n4724 585
R1914 AVSS.n4784 AVSS.n4783 585
R1915 AVSS.n1538 AVSS.n1537 585
R1916 AVSS.n1537 AVSS.n1536 585
R1917 AVSS.n1485 AVSS.n1484 585
R1918 AVSS.n1535 AVSS.n1485 585
R1919 AVSS.n1533 AVSS.n1532 585
R1920 AVSS.n1534 AVSS.n1533 585
R1921 AVSS.n1531 AVSS.n1487 585
R1922 AVSS.n1487 AVSS.n1486 585
R1923 AVSS.n1530 AVSS.n1529 585
R1924 AVSS.n1529 AVSS.n1528 585
R1925 AVSS.n1526 AVSS.n1488 585
R1926 AVSS.n1527 AVSS.n1526 585
R1927 AVSS.n1525 AVSS.n1490 585
R1928 AVSS.n1525 AVSS.n1524 585
R1929 AVSS.n1493 AVSS.n1489 585
R1930 AVSS.n1523 AVSS.n1489 585
R1931 AVSS.n1521 AVSS.n1520 585
R1932 AVSS.n1522 AVSS.n1521 585
R1933 AVSS.n1519 AVSS.n1492 585
R1934 AVSS.n1492 AVSS.n1491 585
R1935 AVSS.n1518 AVSS.n1517 585
R1936 AVSS.n1517 AVSS.n1516 585
R1937 AVSS.n1514 AVSS.n1513 585
R1938 AVSS.n1515 AVSS.n1514 585
R1939 AVSS.n302 AVSS.n300 585
R1940 AVSS.n300 AVSS.n298 585
R1941 AVSS.n358 AVSS.n357 585
R1942 AVSS.n357 AVSS.n356 585
R1943 AVSS.n359 AVSS.n355 585
R1944 AVSS.n355 AVSS.n354 585
R1945 AVSS.n361 AVSS.n360 585
R1946 AVSS.n362 AVSS.n361 585
R1947 AVSS.n353 AVSS.n352 585
R1948 AVSS.n363 AVSS.n353 585
R1949 AVSS.n366 AVSS.n365 585
R1950 AVSS.n365 AVSS.n364 585
R1951 AVSS.n367 AVSS.n351 585
R1952 AVSS.n351 AVSS.n350 585
R1953 AVSS.n369 AVSS.n368 585
R1954 AVSS.n370 AVSS.n369 585
R1955 AVSS.n349 AVSS.n348 585
R1956 AVSS.n371 AVSS.n349 585
R1957 AVSS.n374 AVSS.n373 585
R1958 AVSS.n373 AVSS.n372 585
R1959 AVSS.n375 AVSS.n347 585
R1960 AVSS.n347 AVSS.n346 585
R1961 AVSS.n397 AVSS.n396 585
R1962 AVSS.n398 AVSS.n397 585
R1963 AVSS.n4392 AVSS.n4360 585
R1964 AVSS.n4392 AVSS.n4391 585
R1965 AVSS.n4363 AVSS.n4359 585
R1966 AVSS.n4390 AVSS.n4359 585
R1967 AVSS.n4388 AVSS.n4387 585
R1968 AVSS.n4389 AVSS.n4388 585
R1969 AVSS.n4386 AVSS.n4362 585
R1970 AVSS.n4362 AVSS.n4361 585
R1971 AVSS.n4385 AVSS.n4384 585
R1972 AVSS.n4384 AVSS.n4383 585
R1973 AVSS.n4381 AVSS.n4364 585
R1974 AVSS.n4382 AVSS.n4381 585
R1975 AVSS.n4380 AVSS.n4366 585
R1976 AVSS.n4380 AVSS.n4379 585
R1977 AVSS.n4369 AVSS.n4365 585
R1978 AVSS.n4378 AVSS.n4365 585
R1979 AVSS.n4376 AVSS.n4375 585
R1980 AVSS.n4377 AVSS.n4376 585
R1981 AVSS.n4374 AVSS.n4368 585
R1982 AVSS.n4368 AVSS.n4367 585
R1983 AVSS.n4373 AVSS.n4372 585
R1984 AVSS.n4372 AVSS.n4371 585
R1985 AVSS.n3302 AVSS.n3300 585
R1986 AVSS.n4370 AVSS.n3300 585
R1987 AVSS.n4418 AVSS.n4352 585
R1988 AVSS.n4416 AVSS.n4415 585
R1989 AVSS.n4413 AVSS.n4353 585
R1990 AVSS.n4412 AVSS.n4411 585
R1991 AVSS.n4409 AVSS.n4354 585
R1992 AVSS.n4407 AVSS.n4406 585
R1993 AVSS.n4405 AVSS.n4355 585
R1994 AVSS.n4404 AVSS.n4403 585
R1995 AVSS.n4401 AVSS.n4356 585
R1996 AVSS.n4399 AVSS.n4398 585
R1997 AVSS.n4397 AVSS.n4357 585
R1998 AVSS.n4396 AVSS.n4395 585
R1999 AVSS.n4393 AVSS.n4358 585
R2000 AVSS.n4393 AVSS.n1719 585
R2001 AVSS.n4442 AVSS.n4346 585
R2002 AVSS.n4440 AVSS.n4439 585
R2003 AVSS.n4438 AVSS.n4347 585
R2004 AVSS.n4437 AVSS.n4436 585
R2005 AVSS.n4434 AVSS.n4348 585
R2006 AVSS.n4432 AVSS.n4431 585
R2007 AVSS.n4430 AVSS.n4349 585
R2008 AVSS.n4429 AVSS.n4428 585
R2009 AVSS.n4426 AVSS.n4350 585
R2010 AVSS.n4424 AVSS.n4423 585
R2011 AVSS.n4422 AVSS.n4351 585
R2012 AVSS.n4421 AVSS.n4420 585
R2013 AVSS.n4444 AVSS.n4443 585
R2014 AVSS.n4446 AVSS.n4445 585
R2015 AVSS.n4448 AVSS.n4447 585
R2016 AVSS.n4450 AVSS.n4449 585
R2017 AVSS.n4452 AVSS.n4451 585
R2018 AVSS.n4454 AVSS.n4453 585
R2019 AVSS.n4456 AVSS.n4455 585
R2020 AVSS.n4458 AVSS.n4457 585
R2021 AVSS.n4460 AVSS.n4459 585
R2022 AVSS.n4462 AVSS.n4461 585
R2023 AVSS.n4464 AVSS.n4463 585
R2024 AVSS.n4465 AVSS.n3301 585
R2025 AVSS.n4467 AVSS.n4466 585
R2026 AVSS.n4468 AVSS.n4467 585
R2027 AVSS.t15 AVSS.t117 540.062
R2028 AVSS.n5928 AVSS.n5927 512.543
R2029 AVSS.t6 AVSS.n5966 501.846
R2030 AVSS.n5927 AVSS.n5926 499.428
R2031 AVSS.n431 AVSS.n313 491.875
R2032 AVSS.n5220 AVSS.n14 491.875
R2033 AVSS.n5572 AVSS.n5446 491.875
R2034 AVSS.n5844 AVSS.n5617 491.875
R2035 AVSS.n1536 AVSS.n399 458.238
R2036 AVSS.n4760 AVSS.n886 458.238
R2037 AVSS.n4391 AVSS.n1132 458.238
R2038 AVSS.n3561 AVSS.n2982 458.238
R2039 AVSS.n399 AVSS.n398 449.12
R2040 AVSS.n1515 AVSS.n886 449.12
R2041 AVSS.n4783 AVSS.n1132 449.12
R2042 AVSS.n4370 AVSS.n2982 449.12
R2043 AVSS.n5446 AVSS.n5278 434.043
R2044 AVSS.n5221 AVSS.n5220 434.043
R2045 AVSS.n317 AVSS.n313 434.043
R2046 AVSS.n5845 AVSS.n5844 434.043
R2047 AVSS.t84 AVSS.n197 434.043
R2048 AVSS.t84 AVSS.n207 434.043
R2049 AVSS.t84 AVSS.n201 434.043
R2050 AVSS.t84 AVSS.n203 434.043
R2051 AVSS.t10 AVSS.n5941 429.034
R2052 AVSS.t84 AVSS.n206 424.014
R2053 AVSS.t84 AVSS.n198 424.014
R2054 AVSS.t84 AVSS.n6137 424.014
R2055 AVSS.n6138 AVSS.t84 424.014
R2056 AVSS.n5565 AVSS.n5446 421.277
R2057 AVSS.n5220 AVSS.n5 421.277
R2058 AVSS.n5095 AVSS.n313 421.277
R2059 AVSS.n5844 AVSS.n5843 421.277
R2060 AVSS.t84 AVSS.n208 421.277
R2061 AVSS.t84 AVSS.n200 421.277
R2062 AVSS.t84 AVSS.n204 421.277
R2063 AVSS.t84 AVSS.n166 421.277
R2064 AVSS.n5926 AVSS.n298 348.923
R2065 AVSS.n5901 AVSS.n313 335.981
R2066 AVSS.n5220 AVSS.n5219 335.981
R2067 AVSS.n5446 AVSS.n5445 335.981
R2068 AVSS.n5844 AVSS.n5616 335.981
R2069 AVSS.n5565 AVSS.t90 331.916
R2070 AVSS.t90 AVSS.n5 331.916
R2071 AVSS.n5095 AVSS.t90 331.916
R2072 AVSS.n5843 AVSS.t90 331.916
R2073 AVSS.t80 AVSS.n593 185.648
R2074 AVSS.t80 AVSS.n595 185.648
R2075 AVSS.t80 AVSS.n597 185.648
R2076 AVSS.t80 AVSS.n599 185.648
R2077 AVSS.n2800 AVSS.t76 185.648
R2078 AVSS.n2801 AVSS.t76 185.648
R2079 AVSS.t76 AVSS.n2779 185.648
R2080 AVSS.t76 AVSS.n1726 185.648
R2081 AVSS.t102 AVSS.n208 331.916
R2082 AVSS.t95 AVSS.n200 331.916
R2083 AVSS.t108 AVSS.n204 331.916
R2084 AVSS.t85 AVSS.n166 331.916
R2085 AVSS.n5278 AVSS.t90 319.149
R2086 AVSS.n5221 AVSS.t90 319.149
R2087 AVSS.t90 AVSS.n317 319.149
R2088 AVSS.n5845 AVSS.t90 319.149
R2089 AVSS.t80 AVSS.n592 183.917
R2090 AVSS.t80 AVSS.n594 183.917
R2091 AVSS.t80 AVSS.n596 183.917
R2092 AVSS.t80 AVSS.n598 183.917
R2093 AVSS.n2799 AVSS.t76 183.917
R2094 AVSS.n4498 AVSS.t76 183.917
R2095 AVSS.n2802 AVSS.t76 183.917
R2096 AVSS.n4476 AVSS.t76 183.917
R2097 AVSS.t95 AVSS.n197 319.149
R2098 AVSS.t108 AVSS.n207 319.149
R2099 AVSS.t110 AVSS.n201 319.149
R2100 AVSS.t102 AVSS.n203 319.149
R2101 AVSS.t5 AVSS.n5941 311.154
R2102 AVSS.n5954 AVSS.n5945 309.836
R2103 AVSS.n5958 AVSS.n5945 309.836
R2104 AVSS.n5958 AVSS.n5957 309.836
R2105 AVSS.n5957 AVSS.n5948 307.954
R2106 AVSS.t84 AVSS.n205 289.627
R2107 AVSS.t84 AVSS.n199 289.627
R2108 AVSS.t84 AVSS.n209 289.627
R2109 AVSS.t84 AVSS.n202 289.627
R2110 AVSS.n6055 AVSS.t20 260.437
R2111 AVSS.n546 AVSS.n484 258.334
R2112 AVSS.n1476 AVSS.n1412 258.334
R2113 AVSS.n4896 AVSS.n4832 258.334
R2114 AVSS.n2063 AVSS.n1999 258.334
R2115 AVSS.n1970 AVSS.n1908 258.334
R2116 AVSS.n3389 AVSS.n3326 258.334
R2117 AVSS.n257 AVSS.n256 257.466
R2118 AVSS.n1295 AVSS.n1165 257.466
R2119 AVSS.n4625 AVSS.n1070 257.466
R2120 AVSS.n2115 AVSS.n2089 257.466
R2121 AVSS.n692 AVSS.n690 257.466
R2122 AVSS.n5571 AVSS.n5447 257.466
R2123 AVSS.n6279 AVSS.n11 257.466
R2124 AVSS.n5093 AVSS.n428 257.466
R2125 AVSS.n5924 AVSS.n300 257.466
R2126 AVSS.n5841 AVSS.n5624 257.466
R2127 AVSS.n2279 AVSS.n606 257.466
R2128 AVSS.n2362 AVSS.n626 257.466
R2129 AVSS.n1537 AVSS.n613 257.466
R2130 AVSS.n922 AVSS.n899 257.466
R2131 AVSS.n3219 AVSS.n3091 257.466
R2132 AVSS.n4674 AVSS.n4673 257.466
R2133 AVSS.n4706 AVSS.n4705 257.466
R2134 AVSS.n2940 AVSS.n2938 257.466
R2135 AVSS.n4759 AVSS.n4758 257.466
R2136 AVSS.n2515 AVSS.n1853 257.466
R2137 AVSS.n4293 AVSS.n4292 257.466
R2138 AVSS.n4326 AVSS.n4325 257.466
R2139 AVSS.n3562 AVSS.n3560 257.466
R2140 AVSS.n4260 AVSS.n4259 257.466
R2141 AVSS.n4393 AVSS.n4392 257.466
R2142 AVSS.n6034 AVSS.t15 254.953
R2143 AVSS.n5566 AVSS.n5565 254.34
R2144 AVSS.n5565 AVSS.n5564 254.34
R2145 AVSS.n5565 AVSS.n5453 254.34
R2146 AVSS.n5565 AVSS.n5452 254.34
R2147 AVSS.n5565 AVSS.n5451 254.34
R2148 AVSS.n5565 AVSS.n5450 254.34
R2149 AVSS.n5421 AVSS.n5278 254.34
R2150 AVSS.n5423 AVSS.n5278 254.34
R2151 AVSS.n5429 AVSS.n5278 254.34
R2152 AVSS.n5431 AVSS.n5278 254.34
R2153 AVSS.n5437 AVSS.n5278 254.34
R2154 AVSS.n5439 AVSS.n5278 254.34
R2155 AVSS.n6280 AVSS.n5 254.34
R2156 AVSS.n6282 AVSS.n5 254.34
R2157 AVSS.n6288 AVSS.n5 254.34
R2158 AVSS.n6290 AVSS.n5 254.34
R2159 AVSS.n6296 AVSS.n5 254.34
R2160 AVSS.n6299 AVSS.n5 254.34
R2161 AVSS.n5222 AVSS.n5221 254.34
R2162 AVSS.n5221 AVSS.n415 254.34
R2163 AVSS.n5221 AVSS.n414 254.34
R2164 AVSS.n5221 AVSS.n413 254.34
R2165 AVSS.n5221 AVSS.n412 254.34
R2166 AVSS.n5221 AVSS.n411 254.34
R2167 AVSS.n5880 AVSS.n317 254.34
R2168 AVSS.n323 AVSS.n317 254.34
R2169 AVSS.n5887 AVSS.n317 254.34
R2170 AVSS.n320 AVSS.n317 254.34
R2171 AVSS.n5894 AVSS.n317 254.34
R2172 AVSS.n317 AVSS.n316 254.34
R2173 AVSS.n5095 AVSS.n5094 254.34
R2174 AVSS.n5095 AVSS.n426 254.34
R2175 AVSS.n5095 AVSS.n425 254.34
R2176 AVSS.n5095 AVSS.n424 254.34
R2177 AVSS.n5095 AVSS.n423 254.34
R2178 AVSS.n5096 AVSS.n5095 254.34
R2179 AVSS.n5846 AVSS.n5845 254.34
R2180 AVSS.n5845 AVSS.n5264 254.34
R2181 AVSS.n5845 AVSS.n5263 254.34
R2182 AVSS.n5845 AVSS.n5262 254.34
R2183 AVSS.n5845 AVSS.n5261 254.34
R2184 AVSS.n5845 AVSS.n5260 254.34
R2185 AVSS.n5843 AVSS.n5842 254.34
R2186 AVSS.n5843 AVSS.n5622 254.34
R2187 AVSS.n5843 AVSS.n5621 254.34
R2188 AVSS.n5843 AVSS.n5620 254.34
R2189 AVSS.n5843 AVSS.n5619 254.34
R2190 AVSS.n5843 AVSS.n5618 254.34
R2191 AVSS.n1586 AVSS.n592 254.34
R2192 AVSS.n1580 AVSS.n592 254.34
R2193 AVSS.n1578 AVSS.n592 254.34
R2194 AVSS.n1572 AVSS.n592 254.34
R2195 AVSS.n1570 AVSS.n592 254.34
R2196 AVSS.n1564 AVSS.n592 254.34
R2197 AVSS.n2361 AVSS.n595 254.34
R2198 AVSS.n2311 AVSS.n595 254.34
R2199 AVSS.n2354 AVSS.n595 254.34
R2200 AVSS.n2348 AVSS.n595 254.34
R2201 AVSS.n2346 AVSS.n595 254.34
R2202 AVSS.n2339 AVSS.n595 254.34
R2203 AVSS.n2410 AVSS.n596 254.34
R2204 AVSS.n2305 AVSS.n596 254.34
R2205 AVSS.n2403 AVSS.n596 254.34
R2206 AVSS.n2397 AVSS.n596 254.34
R2207 AVSS.n2395 AVSS.n596 254.34
R2208 AVSS.n2389 AVSS.n596 254.34
R2209 AVSS.n2280 AVSS.n597 254.34
R2210 AVSS.n2282 AVSS.n597 254.34
R2211 AVSS.n2288 AVSS.n597 254.34
R2212 AVSS.n2290 AVSS.n597 254.34
R2213 AVSS.n2296 AVSS.n597 254.34
R2214 AVSS.n2298 AVSS.n597 254.34
R2215 AVSS.n2230 AVSS.n598 254.34
R2216 AVSS.n2237 AVSS.n598 254.34
R2217 AVSS.n2207 AVSS.n598 254.34
R2218 AVSS.n2244 AVSS.n598 254.34
R2219 AVSS.n2204 AVSS.n598 254.34
R2220 AVSS.n2251 AVSS.n598 254.34
R2221 AVSS.n691 AVSS.n599 254.34
R2222 AVSS.n697 AVSS.n599 254.34
R2223 AVSS.n699 AVSS.n599 254.34
R2224 AVSS.n705 AVSS.n599 254.34
R2225 AVSS.n707 AVSS.n599 254.34
R2226 AVSS.n713 AVSS.n599 254.34
R2227 AVSS.n5016 AVSS.n619 254.34
R2228 AVSS.n5016 AVSS.n618 254.34
R2229 AVSS.n5016 AVSS.n617 254.34
R2230 AVSS.n5016 AVSS.n616 254.34
R2231 AVSS.n5016 AVSS.n615 254.34
R2232 AVSS.n5016 AVSS.n614 254.34
R2233 AVSS.n5016 AVSS.n620 254.34
R2234 AVSS.n5016 AVSS.n621 254.34
R2235 AVSS.n5016 AVSS.n622 254.34
R2236 AVSS.n5016 AVSS.n623 254.34
R2237 AVSS.n5016 AVSS.n624 254.34
R2238 AVSS.n5016 AVSS.n625 254.34
R2239 AVSS.n5016 AVSS.n612 254.34
R2240 AVSS.n5016 AVSS.n611 254.34
R2241 AVSS.n5016 AVSS.n610 254.34
R2242 AVSS.n5016 AVSS.n609 254.34
R2243 AVSS.n5016 AVSS.n608 254.34
R2244 AVSS.n5016 AVSS.n607 254.34
R2245 AVSS.n5016 AVSS.n627 254.34
R2246 AVSS.n5016 AVSS.n628 254.34
R2247 AVSS.n5016 AVSS.n629 254.34
R2248 AVSS.n5016 AVSS.n630 254.34
R2249 AVSS.n5016 AVSS.n631 254.34
R2250 AVSS.n5016 AVSS.n632 254.34
R2251 AVSS.n5874 AVSS.n5873 254.34
R2252 AVSS.n5873 AVSS.n345 254.34
R2253 AVSS.n5873 AVSS.n344 254.34
R2254 AVSS.n5873 AVSS.n343 254.34
R2255 AVSS.n5873 AVSS.n342 254.34
R2256 AVSS.n5873 AVSS.n341 254.34
R2257 AVSS.n5873 AVSS.n400 254.34
R2258 AVSS.n5873 AVSS.n401 254.34
R2259 AVSS.n5873 AVSS.n402 254.34
R2260 AVSS.n5873 AVSS.n403 254.34
R2261 AVSS.n5873 AVSS.n404 254.34
R2262 AVSS.n5873 AVSS.n405 254.34
R2263 AVSS.n5873 AVSS.n339 254.34
R2264 AVSS.n5873 AVSS.n338 254.34
R2265 AVSS.n5873 AVSS.n337 254.34
R2266 AVSS.n5873 AVSS.n336 254.34
R2267 AVSS.n5873 AVSS.n335 254.34
R2268 AVSS.n5873 AVSS.n334 254.34
R2269 AVSS.n5873 AVSS.n5249 254.34
R2270 AVSS.n5873 AVSS.n5250 254.34
R2271 AVSS.n5873 AVSS.n5251 254.34
R2272 AVSS.n5873 AVSS.n5252 254.34
R2273 AVSS.n5873 AVSS.n5253 254.34
R2274 AVSS.n5873 AVSS.n5254 254.34
R2275 AVSS.n5873 AVSS.n333 254.34
R2276 AVSS.n5873 AVSS.n332 254.34
R2277 AVSS.n5873 AVSS.n331 254.34
R2278 AVSS.n5873 AVSS.n330 254.34
R2279 AVSS.n5873 AVSS.n329 254.34
R2280 AVSS.n5873 AVSS.n328 254.34
R2281 AVSS.n5016 AVSS.n605 254.34
R2282 AVSS.n5016 AVSS.n604 254.34
R2283 AVSS.n5016 AVSS.n603 254.34
R2284 AVSS.n5016 AVSS.n602 254.34
R2285 AVSS.n5016 AVSS.n601 254.34
R2286 AVSS.n5016 AVSS.n600 254.34
R2287 AVSS.n923 AVSS.n593 254.34
R2288 AVSS.n925 AVSS.n593 254.34
R2289 AVSS.n931 AVSS.n593 254.34
R2290 AVSS.n933 AVSS.n593 254.34
R2291 AVSS.n939 AVSS.n593 254.34
R2292 AVSS.n941 AVSS.n593 254.34
R2293 AVSS.n4995 AVSS.n594 254.34
R2294 AVSS.n643 AVSS.n594 254.34
R2295 AVSS.n5002 AVSS.n594 254.34
R2296 AVSS.n640 AVSS.n594 254.34
R2297 AVSS.n5009 AVSS.n594 254.34
R2298 AVSS.n637 AVSS.n594 254.34
R2299 AVSS.n3118 AVSS.n2801 254.34
R2300 AVSS.n3116 AVSS.n2801 254.34
R2301 AVSS.n3110 AVSS.n2801 254.34
R2302 AVSS.n3108 AVSS.n2801 254.34
R2303 AVSS.n3102 AVSS.n2801 254.34
R2304 AVSS.n3100 AVSS.n2801 254.34
R2305 AVSS.n4498 AVSS.n2796 254.34
R2306 AVSS.n4498 AVSS.n2795 254.34
R2307 AVSS.n4498 AVSS.n2794 254.34
R2308 AVSS.n4498 AVSS.n2793 254.34
R2309 AVSS.n4498 AVSS.n2792 254.34
R2310 AVSS.n4499 AVSS.n4498 254.34
R2311 AVSS.n4675 AVSS.n2779 254.34
R2312 AVSS.n2841 AVSS.n2779 254.34
R2313 AVSS.n2846 AVSS.n2779 254.34
R2314 AVSS.n2848 AVSS.n2779 254.34
R2315 AVSS.n2854 AVSS.n2779 254.34
R2316 AVSS.n2857 AVSS.n2779 254.34
R2317 AVSS.n3038 AVSS.n2802 254.34
R2318 AVSS.n3032 AVSS.n2802 254.34
R2319 AVSS.n3030 AVSS.n2802 254.34
R2320 AVSS.n3024 AVSS.n2802 254.34
R2321 AVSS.n3022 AVSS.n2802 254.34
R2322 AVSS.n3018 AVSS.n2802 254.34
R2323 AVSS.n4707 AVSS.n1726 254.34
R2324 AVSS.n2994 AVSS.n1726 254.34
R2325 AVSS.n2999 AVSS.n1726 254.34
R2326 AVSS.n3001 AVSS.n1726 254.34
R2327 AVSS.n3007 AVSS.n1726 254.34
R2328 AVSS.n3009 AVSS.n1726 254.34
R2329 AVSS.n4476 AVSS.n4475 254.34
R2330 AVSS.n4476 AVSS.n2806 254.34
R2331 AVSS.n4476 AVSS.n2805 254.34
R2332 AVSS.n4476 AVSS.n2804 254.34
R2333 AVSS.n4476 AVSS.n2803 254.34
R2334 AVSS.n4476 AVSS.n1720 254.34
R2335 AVSS.n2939 AVSS.n2800 254.34
R2336 AVSS.n2945 AVSS.n2800 254.34
R2337 AVSS.n2947 AVSS.n2800 254.34
R2338 AVSS.n2953 AVSS.n2800 254.34
R2339 AVSS.n2909 AVSS.n2800 254.34
R2340 AVSS.n2960 AVSS.n2800 254.34
R2341 AVSS.n4717 AVSS.n1719 254.34
R2342 AVSS.n2922 AVSS.n1719 254.34
R2343 AVSS.n2921 AVSS.n1719 254.34
R2344 AVSS.n2929 AVSS.n1719 254.34
R2345 AVSS.n2918 AVSS.n1719 254.34
R2346 AVSS.n2936 AVSS.n1719 254.34
R2347 AVSS.n4685 AVSS.n1719 254.34
R2348 AVSS.n1735 AVSS.n1719 254.34
R2349 AVSS.n4692 AVSS.n1719 254.34
R2350 AVSS.n1732 AVSS.n1719 254.34
R2351 AVSS.n4699 AVSS.n1719 254.34
R2352 AVSS.n1729 AVSS.n1719 254.34
R2353 AVSS.n4505 AVSS.n1719 254.34
R2354 AVSS.n2788 AVSS.n1719 254.34
R2355 AVSS.n4512 AVSS.n1719 254.34
R2356 AVSS.n2785 AVSS.n1719 254.34
R2357 AVSS.n4519 AVSS.n1719 254.34
R2358 AVSS.n2782 AVSS.n1719 254.34
R2359 AVSS.n3085 AVSS.n1719 254.34
R2360 AVSS.n3236 AVSS.n1719 254.34
R2361 AVSS.n3230 AVSS.n1719 254.34
R2362 AVSS.n3228 AVSS.n1719 254.34
R2363 AVSS.n3222 AVSS.n1719 254.34
R2364 AVSS.n3220 AVSS.n1719 254.34
R2365 AVSS.n4933 AVSS.n1133 254.34
R2366 AVSS.n4933 AVSS.n1134 254.34
R2367 AVSS.n4933 AVSS.n1135 254.34
R2368 AVSS.n4933 AVSS.n1136 254.34
R2369 AVSS.n4933 AVSS.n1137 254.34
R2370 AVSS.n4933 AVSS.n1138 254.34
R2371 AVSS.n4934 AVSS.n4933 254.34
R2372 AVSS.n4933 AVSS.n1131 254.34
R2373 AVSS.n4933 AVSS.n1130 254.34
R2374 AVSS.n4933 AVSS.n1129 254.34
R2375 AVSS.n4933 AVSS.n1128 254.34
R2376 AVSS.n4933 AVSS.n1127 254.34
R2377 AVSS.n4933 AVSS.n1140 254.34
R2378 AVSS.n4933 AVSS.n1141 254.34
R2379 AVSS.n4933 AVSS.n1142 254.34
R2380 AVSS.n4933 AVSS.n1143 254.34
R2381 AVSS.n4933 AVSS.n1144 254.34
R2382 AVSS.n4933 AVSS.n1368 254.34
R2383 AVSS.n4933 AVSS.n1125 254.34
R2384 AVSS.n4933 AVSS.n1124 254.34
R2385 AVSS.n4933 AVSS.n1123 254.34
R2386 AVSS.n4933 AVSS.n1122 254.34
R2387 AVSS.n4933 AVSS.n1121 254.34
R2388 AVSS.n4933 AVSS.n1120 254.34
R2389 AVSS.n4927 AVSS.n4926 254.34
R2390 AVSS.n4926 AVSS.n4925 254.34
R2391 AVSS.n4926 AVSS.n1377 254.34
R2392 AVSS.n4926 AVSS.n1376 254.34
R2393 AVSS.n4926 AVSS.n1375 254.34
R2394 AVSS.n4926 AVSS.n1374 254.34
R2395 AVSS.n2116 AVSS.n2083 254.34
R2396 AVSS.n2118 AVSS.n2083 254.34
R2397 AVSS.n2124 AVSS.n2083 254.34
R2398 AVSS.n2126 AVSS.n2083 254.34
R2399 AVSS.n2132 AVSS.n2083 254.34
R2400 AVSS.n2135 AVSS.n2083 254.34
R2401 AVSS.n2162 AVSS.n2073 254.34
R2402 AVSS.n2169 AVSS.n2073 254.34
R2403 AVSS.n2079 AVSS.n2073 254.34
R2404 AVSS.n2176 AVSS.n2073 254.34
R2405 AVSS.n2076 AVSS.n2073 254.34
R2406 AVSS.n2183 AVSS.n2073 254.34
R2407 AVSS.n4626 AVSS.n4618 254.34
R2408 AVSS.n4628 AVSS.n4618 254.34
R2409 AVSS.n4634 AVSS.n4618 254.34
R2410 AVSS.n4636 AVSS.n4618 254.34
R2411 AVSS.n4642 AVSS.n4618 254.34
R2412 AVSS.n4645 AVSS.n4618 254.34
R2413 AVSS.n4940 AVSS.n1082 254.34
R2414 AVSS.n1088 AVSS.n1082 254.34
R2415 AVSS.n4947 AVSS.n1082 254.34
R2416 AVSS.n1085 AVSS.n1082 254.34
R2417 AVSS.n4954 AVSS.n1082 254.34
R2418 AVSS.n1082 AVSS.n1081 254.34
R2419 AVSS.n1193 AVSS.n1192 254.34
R2420 AVSS.n1192 AVSS.n1191 254.34
R2421 AVSS.n1192 AVSS.n1171 254.34
R2422 AVSS.n1192 AVSS.n1170 254.34
R2423 AVSS.n1192 AVSS.n1169 254.34
R2424 AVSS.n1192 AVSS.n1168 254.34
R2425 AVSS.n4906 AVSS.n1071 254.34
R2426 AVSS.n4740 AVSS.n1071 254.34
R2427 AVSS.n4745 AVSS.n1071 254.34
R2428 AVSS.n4739 AVSS.n1071 254.34
R2429 AVSS.n4752 AVSS.n1071 254.34
R2430 AVSS.n4736 AVSS.n1071 254.34
R2431 AVSS.n2186 AVSS.n1071 254.34
R2432 AVSS.n2095 AVSS.n1071 254.34
R2433 AVSS.n2100 AVSS.n1071 254.34
R2434 AVSS.n2094 AVSS.n1071 254.34
R2435 AVSS.n2107 AVSS.n1071 254.34
R2436 AVSS.n2110 AVSS.n1071 254.34
R2437 AVSS.n4961 AVSS.n1071 254.34
R2438 AVSS.n1078 AVSS.n1071 254.34
R2439 AVSS.n4968 AVSS.n1071 254.34
R2440 AVSS.n1075 AVSS.n1071 254.34
R2441 AVSS.n4975 AVSS.n1071 254.34
R2442 AVSS.n4978 AVSS.n1071 254.34
R2443 AVSS.n1159 AVSS.n1071 254.34
R2444 AVSS.n1312 AVSS.n1071 254.34
R2445 AVSS.n1306 AVSS.n1071 254.34
R2446 AVSS.n1304 AVSS.n1071 254.34
R2447 AVSS.n1298 AVSS.n1071 254.34
R2448 AVSS.n1296 AVSS.n1071 254.34
R2449 AVSS.n4988 AVSS.n667 254.34
R2450 AVSS.n4988 AVSS.n666 254.34
R2451 AVSS.n4988 AVSS.n665 254.34
R2452 AVSS.n4988 AVSS.n664 254.34
R2453 AVSS.n4988 AVSS.n663 254.34
R2454 AVSS.n4988 AVSS.n662 254.34
R2455 AVSS.n4989 AVSS.n4988 254.34
R2456 AVSS.n4988 AVSS.n887 254.34
R2457 AVSS.n4988 AVSS.n888 254.34
R2458 AVSS.n4988 AVSS.n889 254.34
R2459 AVSS.n4988 AVSS.n890 254.34
R2460 AVSS.n4988 AVSS.n891 254.34
R2461 AVSS.n4988 AVSS.n660 254.34
R2462 AVSS.n4988 AVSS.n659 254.34
R2463 AVSS.n4988 AVSS.n658 254.34
R2464 AVSS.n4988 AVSS.n657 254.34
R2465 AVSS.n4988 AVSS.n656 254.34
R2466 AVSS.n4988 AVSS.n655 254.34
R2467 AVSS.n4988 AVSS.n965 254.34
R2468 AVSS.n4988 AVSS.n966 254.34
R2469 AVSS.n4988 AVSS.n967 254.34
R2470 AVSS.n4988 AVSS.n968 254.34
R2471 AVSS.n4988 AVSS.n969 254.34
R2472 AVSS.n4988 AVSS.n970 254.34
R2473 AVSS.n4988 AVSS.n653 254.34
R2474 AVSS.n4988 AVSS.n652 254.34
R2475 AVSS.n4988 AVSS.n651 254.34
R2476 AVSS.n4988 AVSS.n650 254.34
R2477 AVSS.n4988 AVSS.n649 254.34
R2478 AVSS.n4988 AVSS.n648 254.34
R2479 AVSS.n1865 AVSS.n1071 254.34
R2480 AVSS.n1867 AVSS.n1071 254.34
R2481 AVSS.n1873 AVSS.n1071 254.34
R2482 AVSS.n1875 AVSS.n1071 254.34
R2483 AVSS.n1881 AVSS.n1071 254.34
R2484 AVSS.n1883 AVSS.n1071 254.34
R2485 AVSS.n2583 AVSS.n2582 254.34
R2486 AVSS.n2582 AVSS.n2581 254.34
R2487 AVSS.n2582 AVSS.n1745 254.34
R2488 AVSS.n2582 AVSS.n1744 254.34
R2489 AVSS.n2582 AVSS.n1743 254.34
R2490 AVSS.n2582 AVSS.n1742 254.34
R2491 AVSS.n4933 AVSS.n1118 254.34
R2492 AVSS.n4933 AVSS.n1117 254.34
R2493 AVSS.n4933 AVSS.n1116 254.34
R2494 AVSS.n4933 AVSS.n1115 254.34
R2495 AVSS.n4933 AVSS.n1114 254.34
R2496 AVSS.n4933 AVSS.n1113 254.34
R2497 AVSS.n2516 AVSS.n1847 254.34
R2498 AVSS.n2518 AVSS.n1847 254.34
R2499 AVSS.n2524 AVSS.n1847 254.34
R2500 AVSS.n2526 AVSS.n1847 254.34
R2501 AVSS.n2532 AVSS.n1847 254.34
R2502 AVSS.n2535 AVSS.n1847 254.34
R2503 AVSS.n3969 AVSS.n197 254.34
R2504 AVSS.n3971 AVSS.n197 254.34
R2505 AVSS.n3977 AVSS.n197 254.34
R2506 AVSS.n3979 AVSS.n197 254.34
R2507 AVSS.n3985 AVSS.n197 254.34
R2508 AVSS.n3987 AVSS.n197 254.34
R2509 AVSS.n4294 AVSS.n200 254.34
R2510 AVSS.n3923 AVSS.n200 254.34
R2511 AVSS.n3928 AVSS.n200 254.34
R2512 AVSS.n3930 AVSS.n200 254.34
R2513 AVSS.n3936 AVSS.n200 254.34
R2514 AVSS.n3939 AVSS.n200 254.34
R2515 AVSS.n3758 AVSS.n207 254.34
R2516 AVSS.n3760 AVSS.n207 254.34
R2517 AVSS.n3766 AVSS.n207 254.34
R2518 AVSS.n3768 AVSS.n207 254.34
R2519 AVSS.n3774 AVSS.n207 254.34
R2520 AVSS.n3776 AVSS.n207 254.34
R2521 AVSS.n4327 AVSS.n204 254.34
R2522 AVSS.n3712 AVSS.n204 254.34
R2523 AVSS.n3717 AVSS.n204 254.34
R2524 AVSS.n3719 AVSS.n204 254.34
R2525 AVSS.n3725 AVSS.n204 254.34
R2526 AVSS.n3728 AVSS.n204 254.34
R2527 AVSS.n3621 AVSS.n201 254.34
R2528 AVSS.n3623 AVSS.n201 254.34
R2529 AVSS.n3629 AVSS.n201 254.34
R2530 AVSS.n3631 AVSS.n201 254.34
R2531 AVSS.n3637 AVSS.n201 254.34
R2532 AVSS.n3514 AVSS.n201 254.34
R2533 AVSS.n4338 AVSS.n151 254.34
R2534 AVSS.n3544 AVSS.n151 254.34
R2535 AVSS.n3543 AVSS.n151 254.34
R2536 AVSS.n3551 AVSS.n151 254.34
R2537 AVSS.n3540 AVSS.n151 254.34
R2538 AVSS.n3558 AVSS.n151 254.34
R2539 AVSS.n4305 AVSS.n151 254.34
R2540 AVSS.n3689 AVSS.n151 254.34
R2541 AVSS.n4312 AVSS.n151 254.34
R2542 AVSS.n3686 AVSS.n151 254.34
R2543 AVSS.n4319 AVSS.n151 254.34
R2544 AVSS.n3683 AVSS.n151 254.34
R2545 AVSS.n4272 AVSS.n151 254.34
R2546 AVSS.n3900 AVSS.n151 254.34
R2547 AVSS.n4279 AVSS.n151 254.34
R2548 AVSS.n3897 AVSS.n151 254.34
R2549 AVSS.n4286 AVSS.n151 254.34
R2550 AVSS.n3894 AVSS.n151 254.34
R2551 AVSS.n6192 AVSS.n151 254.34
R2552 AVSS.n157 AVSS.n151 254.34
R2553 AVSS.n6199 AVSS.n151 254.34
R2554 AVSS.n154 AVSS.n151 254.34
R2555 AVSS.n6206 AVSS.n151 254.34
R2556 AVSS.n151 AVSS.n150 254.34
R2557 AVSS.n4469 AVSS.n4468 254.34
R2558 AVSS.n4468 AVSS.n2981 254.34
R2559 AVSS.n4468 AVSS.n2906 254.34
R2560 AVSS.n4468 AVSS.n2905 254.34
R2561 AVSS.n4468 AVSS.n2904 254.34
R2562 AVSS.n4468 AVSS.n2903 254.34
R2563 AVSS.n4468 AVSS.n2983 254.34
R2564 AVSS.n4468 AVSS.n2984 254.34
R2565 AVSS.n4468 AVSS.n2985 254.34
R2566 AVSS.n4468 AVSS.n2986 254.34
R2567 AVSS.n4468 AVSS.n2987 254.34
R2568 AVSS.n4468 AVSS.n2988 254.34
R2569 AVSS.n4468 AVSS.n2901 254.34
R2570 AVSS.n4468 AVSS.n2834 254.34
R2571 AVSS.n4468 AVSS.n2833 254.34
R2572 AVSS.n4468 AVSS.n2832 254.34
R2573 AVSS.n4468 AVSS.n2831 254.34
R2574 AVSS.n4468 AVSS.n2830 254.34
R2575 AVSS.n4468 AVSS.n3065 254.34
R2576 AVSS.n4468 AVSS.n3066 254.34
R2577 AVSS.n4468 AVSS.n3067 254.34
R2578 AVSS.n4468 AVSS.n3068 254.34
R2579 AVSS.n4468 AVSS.n3069 254.34
R2580 AVSS.n4468 AVSS.n3293 254.34
R2581 AVSS.n4238 AVSS.n151 254.34
R2582 AVSS.n4240 AVSS.n151 254.34
R2583 AVSS.n4246 AVSS.n151 254.34
R2584 AVSS.n4248 AVSS.n151 254.34
R2585 AVSS.n4254 AVSS.n151 254.34
R2586 AVSS.n4230 AVSS.n151 254.34
R2587 AVSS.n4261 AVSS.n208 254.34
R2588 AVSS.n4228 AVSS.n208 254.34
R2589 AVSS.n4222 AVSS.n208 254.34
R2590 AVSS.n4220 AVSS.n208 254.34
R2591 AVSS.n4214 AVSS.n208 254.34
R2592 AVSS.n4212 AVSS.n208 254.34
R2593 AVSS.n6107 AVSS.n203 254.34
R2594 AVSS.n6105 AVSS.n203 254.34
R2595 AVSS.n6099 AVSS.n203 254.34
R2596 AVSS.n6097 AVSS.n203 254.34
R2597 AVSS.n6091 AVSS.n203 254.34
R2598 AVSS.n6089 AVSS.n203 254.34
R2599 AVSS.n258 AVSS.n166 254.34
R2600 AVSS.n254 AVSS.n166 254.34
R2601 AVSS.n248 AVSS.n166 254.34
R2602 AVSS.n246 AVSS.n166 254.34
R2603 AVSS.n240 AVSS.n166 254.34
R2604 AVSS.n238 AVSS.n166 254.34
R2605 AVSS.n4417 AVSS.n1719 254.34
R2606 AVSS.n4410 AVSS.n1719 254.34
R2607 AVSS.n4408 AVSS.n1719 254.34
R2608 AVSS.n4402 AVSS.n1719 254.34
R2609 AVSS.n4400 AVSS.n1719 254.34
R2610 AVSS.n4394 AVSS.n1719 254.34
R2611 AVSS.n4441 AVSS.n2799 254.34
R2612 AVSS.n4435 AVSS.n2799 254.34
R2613 AVSS.n4433 AVSS.n2799 254.34
R2614 AVSS.n4427 AVSS.n2799 254.34
R2615 AVSS.n4425 AVSS.n2799 254.34
R2616 AVSS.n4419 AVSS.n2799 254.34
R2617 AVSS.n4468 AVSS.n3294 254.34
R2618 AVSS.n4468 AVSS.n3295 254.34
R2619 AVSS.n4468 AVSS.n3296 254.34
R2620 AVSS.n4468 AVSS.n3297 254.34
R2621 AVSS.n4468 AVSS.n3298 254.34
R2622 AVSS.n4468 AVSS.n3299 254.34
R2623 AVSS.n144 AVSS.n58 250
R2624 AVSS.n4202 AVSS.n4116 250
R2625 AVSS.n4060 AVSS.n3996 250
R2626 AVSS.n3849 AVSS.n3785 250
R2627 AVSS.n3490 AVSS.n3426 250
R2628 AVSS.n5795 AVSS.n5746 250
R2629 AVSS.n5523 AVSS.n5474 250
R2630 AVSS.n5356 AVSS.n5354 250
R2631 AVSS.n5157 AVSS.n5155 250
R2632 AVSS.n3212 AVSS.n3125 250
R2633 AVSS.n1288 AVSS.n1201 250
R2634 AVSS.n4592 AVSS.n4543 250
R2635 AVSS.n2772 AVSS.n2686 250
R2636 AVSS.n2662 AVSS.n2598 250
R2637 AVSS.n1695 AVSS.n1631 250
R2638 AVSS.n829 AVSS.n742 250
R2639 AVSS.n1043 AVSS.n994 250
R2640 AVSS.n2489 AVSS.n2487 250
R2641 AVSS.n1784 AVSS.n1770 250
R2642 AVSS.n6139 AVSS.n186 249.663
R2643 AVSS.n1174 AVSS.n1145 249.663
R2644 AVSS.n4646 AVSS.n1126 249.663
R2645 AVSS.n2136 AVSS.n1139 249.663
R2646 AVSS.n715 AVSS.n714 249.663
R2647 AVSS.n5872 AVSS.n5255 249.663
R2648 AVSS.n6300 AVSS.n4 249.663
R2649 AVSS.n5248 AVSS.n406 249.663
R2650 AVSS.n397 AVSS.n340 249.663
R2651 AVSS.n5628 AVSS.n5627 249.663
R2652 AVSS.n4987 AVSS.n971 249.663
R2653 AVSS.n2340 AVSS.n654 249.663
R2654 AVSS.n1514 AVSS.n661 249.663
R2655 AVSS.n964 AVSS.n892 249.663
R2656 AVSS.n3099 AVSS.n3070 249.663
R2657 AVSS.n2858 AVSS.n2829 249.663
R2658 AVSS.n3064 AVSS.n2989 249.663
R2659 AVSS.n2961 AVSS.n2902 249.663
R2660 AVSS.n4785 AVSS.n4784 249.663
R2661 AVSS.n2536 AVSS.n1846 249.663
R2662 AVSS.n3940 AVSS.n3918 249.663
R2663 AVSS.n3729 AVSS.n3707 249.663
R2664 AVSS.n3592 AVSS.n3576 249.663
R2665 AVSS.n6136 AVSS.n211 249.663
R2666 AVSS.n4467 AVSS.n3300 249.663
R2667 AVSS.n6057 AVSS.n295 248.843
R2668 AVSS.n5910 AVSS.n5909 241.906
R2669 AVSS.n5909 AVSS.n309 241.906
R2670 AVSS.n5903 AVSS.n309 241.906
R2671 AVSS.n5903 AVSS.n5902 241.906
R2672 AVSS.n5902 AVSS.n5901 241.906
R2673 AVSS.n5073 AVSS.n431 241.906
R2674 AVSS.n5073 AVSS.n5072 241.906
R2675 AVSS.n5072 AVSS.n5071 241.906
R2676 AVSS.n5071 AVSS.n432 241.906
R2677 AVSS.n5065 AVSS.n432 241.906
R2678 AVSS.n448 AVSS.n447 241.906
R2679 AVSS.n447 AVSS.n436 241.906
R2680 AVSS.n441 AVSS.n436 241.906
R2681 AVSS.n441 AVSS.n440 241.906
R2682 AVSS.n440 AVSS.n416 241.906
R2683 AVSS.n5219 AVSS.n416 241.906
R2684 AVSS.n6274 AVSS.n14 241.906
R2685 AVSS.n6274 AVSS.n6273 241.906
R2686 AVSS.n6273 AVSS.n6272 241.906
R2687 AVSS.n6272 AVSS.n15 241.906
R2688 AVSS.n6266 AVSS.n15 241.906
R2689 AVSS.n5284 AVSS.n19 241.906
R2690 AVSS.n5289 AVSS.n5284 241.906
R2691 AVSS.n5290 AVSS.n5289 241.906
R2692 AVSS.n5291 AVSS.n5290 241.906
R2693 AVSS.n5291 AVSS.n5279 241.906
R2694 AVSS.n5445 AVSS.n5279 241.906
R2695 AVSS.n5573 AVSS.n5572 241.906
R2696 AVSS.n5574 AVSS.n5573 241.906
R2697 AVSS.n5574 AVSS.n5274 241.906
R2698 AVSS.n5580 AVSS.n5274 241.906
R2699 AVSS.n5581 AVSS.n5580 241.906
R2700 AVSS.n5582 AVSS.n5270 241.906
R2701 AVSS.n5588 AVSS.n5270 241.906
R2702 AVSS.n5589 AVSS.n5588 241.906
R2703 AVSS.n5590 AVSS.n5589 241.906
R2704 AVSS.n5590 AVSS.n5265 241.906
R2705 AVSS.n5616 AVSS.n5265 241.906
R2706 AVSS.n5650 AVSS.n5617 241.906
R2707 AVSS.n5656 AVSS.n5650 241.906
R2708 AVSS.n5657 AVSS.n5656 241.906
R2709 AVSS.n5658 AVSS.n5657 241.906
R2710 AVSS.n5658 AVSS.n36 241.906
R2711 AVSS.n5665 AVSS.n37 241.906
R2712 AVSS.n5666 AVSS.n5665 241.906
R2713 AVSS.n5667 AVSS.n5666 241.906
R2714 AVSS.n5667 AVSS.n5643 241.906
R2715 AVSS.n5673 AVSS.n5643 241.906
R2716 AVSS.t47 AVSS.n5940 228.911
R2717 AVSS.t123 AVSS.t37 227.54
R2718 AVSS.t37 AVSS.t51 227.54
R2719 AVSS.t128 AVSS.t25 227.54
R2720 AVSS.t20 AVSS.t128 227.54
R2721 AVSS.n119 AVSS.n118 221.667
R2722 AVSS.n5761 AVSS.n5760 221.667
R2723 AVSS.n5489 AVSS.n5488 221.667
R2724 AVSS.n5390 AVSS.n5303 221.667
R2725 AVSS.n5191 AVSS.n5104 221.667
R2726 AVSS.n3193 AVSS.n3192 221.667
R2727 AVSS.n1269 AVSS.n1268 221.667
R2728 AVSS.n4558 AVSS.n4557 221.667
R2729 AVSS.n2747 AVSS.n2746 221.667
R2730 AVSS.n810 AVSS.n809 221.667
R2731 AVSS.n1009 AVSS.n1008 221.667
R2732 AVSS.n2455 AVSS.n2435 221.667
R2733 AVSS.n1805 AVSS.n1804 221.667
R2734 AVSS.t2 AVSS.n5960 212.462
R2735 AVSS.n3591 AVSS.n3590 208.531
R2736 AVSS.n3590 AVSS.n3589 208.531
R2737 AVSS.n3589 AVSS.n3579 208.531
R2738 AVSS.n3583 AVSS.n3579 208.531
R2739 AVSS.n3583 AVSS.n3527 208.531
R2740 AVSS.n3607 AVSS.n3606 208.531
R2741 AVSS.n3607 AVSS.n3523 208.531
R2742 AVSS.n3613 AVSS.n3523 208.531
R2743 AVSS.n3614 AVSS.n3613 208.531
R2744 AVSS.n3615 AVSS.n3614 208.531
R2745 AVSS.n3615 AVSS.n205 208.531
R2746 AVSS.n3734 AVSS.n206 208.531
R2747 AVSS.n3735 AVSS.n3734 208.531
R2748 AVSS.n3736 AVSS.n3735 208.531
R2749 AVSS.n3736 AVSS.n3703 208.531
R2750 AVSS.n3742 AVSS.n3703 208.531
R2751 AVSS.n3744 AVSS.n3743 208.531
R2752 AVSS.n3744 AVSS.n3699 208.531
R2753 AVSS.n3750 AVSS.n3699 208.531
R2754 AVSS.n3751 AVSS.n3750 208.531
R2755 AVSS.n3752 AVSS.n3751 208.531
R2756 AVSS.n3752 AVSS.n199 208.531
R2757 AVSS.n3945 AVSS.n198 208.531
R2758 AVSS.n3946 AVSS.n3945 208.531
R2759 AVSS.n3947 AVSS.n3946 208.531
R2760 AVSS.n3947 AVSS.n3914 208.531
R2761 AVSS.n3953 AVSS.n3914 208.531
R2762 AVSS.n3955 AVSS.n3954 208.531
R2763 AVSS.n3955 AVSS.n3910 208.531
R2764 AVSS.n3961 AVSS.n3910 208.531
R2765 AVSS.n3962 AVSS.n3961 208.531
R2766 AVSS.n3963 AVSS.n3962 208.531
R2767 AVSS.n3963 AVSS.n209 208.531
R2768 AVSS.n6137 AVSS.n210 208.531
R2769 AVSS.n6131 AVSS.n210 208.531
R2770 AVSS.n6131 AVSS.n6130 208.531
R2771 AVSS.n6130 AVSS.n6129 208.531
R2772 AVSS.n6129 AVSS.n216 208.531
R2773 AVSS.n6123 AVSS.n6122 208.531
R2774 AVSS.n6122 AVSS.n6121 208.531
R2775 AVSS.n6121 AVSS.n220 208.531
R2776 AVSS.n6115 AVSS.n220 208.531
R2777 AVSS.n6115 AVSS.n6114 208.531
R2778 AVSS.n6114 AVSS.n202 208.531
R2779 AVSS.n6138 AVSS.n183 208.531
R2780 AVSS.n6144 AVSS.n183 208.531
R2781 AVSS.n6145 AVSS.n6144 208.531
R2782 AVSS.n6146 AVSS.n6145 208.531
R2783 AVSS.n6146 AVSS.n167 208.531
R2784 AVSS.n6153 AVSS.n168 208.531
R2785 AVSS.n6154 AVSS.n6153 208.531
R2786 AVSS.n6154 AVSS.n177 208.531
R2787 AVSS.n6160 AVSS.n177 208.531
R2788 AVSS.n6161 AVSS.n6160 208.531
R2789 AVSS.n5942 AVSS.t0 205.607
R2790 AVSS.n356 AVSS.n298 205.181
R2791 AVSS.n356 AVSS.n354 205.181
R2792 AVSS.n362 AVSS.n354 205.181
R2793 AVSS.n363 AVSS.n362 205.181
R2794 AVSS.n364 AVSS.n363 205.181
R2795 AVSS.n370 AVSS.n350 205.181
R2796 AVSS.n371 AVSS.n370 205.181
R2797 AVSS.n372 AVSS.n371 205.181
R2798 AVSS.n372 AVSS.n346 205.181
R2799 AVSS.n398 AVSS.n346 205.181
R2800 AVSS.n1536 AVSS.n1535 205.181
R2801 AVSS.n1535 AVSS.n1534 205.181
R2802 AVSS.n1534 AVSS.n1486 205.181
R2803 AVSS.n1528 AVSS.n1486 205.181
R2804 AVSS.n1528 AVSS.n1527 205.181
R2805 AVSS.n1524 AVSS.n1523 205.181
R2806 AVSS.n1523 AVSS.n1522 205.181
R2807 AVSS.n1522 AVSS.n1491 205.181
R2808 AVSS.n1516 AVSS.n1491 205.181
R2809 AVSS.n1516 AVSS.n1515 205.181
R2810 AVSS.n4761 AVSS.n4760 205.181
R2811 AVSS.n4761 AVSS.n4731 205.181
R2812 AVSS.n4768 AVSS.n4731 205.181
R2813 AVSS.n4769 AVSS.n4768 205.181
R2814 AVSS.n4770 AVSS.n4769 205.181
R2815 AVSS.n4774 AVSS.n4773 205.181
R2816 AVSS.n4774 AVSS.n4726 205.181
R2817 AVSS.n4781 AVSS.n4726 205.181
R2818 AVSS.n4782 AVSS.n4781 205.181
R2819 AVSS.n4783 AVSS.n4782 205.181
R2820 AVSS.n4391 AVSS.n4390 205.181
R2821 AVSS.n4390 AVSS.n4389 205.181
R2822 AVSS.n4389 AVSS.n4361 205.181
R2823 AVSS.n4383 AVSS.n4361 205.181
R2824 AVSS.n4383 AVSS.n4382 205.181
R2825 AVSS.n4379 AVSS.n4378 205.181
R2826 AVSS.n4378 AVSS.n4377 205.181
R2827 AVSS.n4377 AVSS.n4367 205.181
R2828 AVSS.n4371 AVSS.n4367 205.181
R2829 AVSS.n4371 AVSS.n4370 205.181
R2830 AVSS.n3561 AVSS.n3534 205.181
R2831 AVSS.n3567 AVSS.n3534 205.181
R2832 AVSS.n3568 AVSS.n3567 205.181
R2833 AVSS.n3569 AVSS.n3568 205.181
R2834 AVSS.n3569 AVSS.n3528 205.181
R2835 AVSS.n3605 AVSS.n3529 205.181
R2836 AVSS.n3599 AVSS.n3529 205.181
R2837 AVSS.n3599 AVSS.n3598 205.181
R2838 AVSS.n3598 AVSS.n3597 205.181
R2839 AVSS.n3597 AVSS.n3575 205.181
R2840 AVSS.t44 AVSS.t7 202.798
R2841 AVSS.t47 AVSS.t5 198.762
R2842 AVSS.t15 AVSS.t117 198.762
R2843 AVSS.n2083 AVSS.t78 185.648
R2844 AVSS.n1847 AVSS.t78 185.648
R2845 AVSS.n4618 AVSS.t78 185.648
R2846 AVSS.n1192 AVSS.t78 185.648
R2847 AVSS.n58 AVSS.n56 185
R2848 AVSS.n79 AVSS.n78 185
R2849 AVSS.n81 AVSS.n80 185
R2850 AVSS.n83 AVSS.n82 185
R2851 AVSS.n85 AVSS.n84 185
R2852 AVSS.n86 AVSS.n77 185
R2853 AVSS.n141 AVSS.n140 185
R2854 AVSS.n139 AVSS.n76 185
R2855 AVSS.n138 AVSS.n137 185
R2856 AVSS.n120 AVSS.n119 185
R2857 AVSS.n122 AVSS.n121 185
R2858 AVSS.n124 AVSS.n123 185
R2859 AVSS.n126 AVSS.n125 185
R2860 AVSS.n128 AVSS.n127 185
R2861 AVSS.n130 AVSS.n129 185
R2862 AVSS.n132 AVSS.n131 185
R2863 AVSS.n134 AVSS.n133 185
R2864 AVSS.n136 AVSS.n135 185
R2865 AVSS.n118 AVSS.n117 185
R2866 AVSS.n116 AVSS.n115 185
R2867 AVSS.n114 AVSS.n113 185
R2868 AVSS.n112 AVSS.n111 185
R2869 AVSS.n110 AVSS.n109 185
R2870 AVSS.n108 AVSS.n107 185
R2871 AVSS.n106 AVSS.n105 185
R2872 AVSS.n104 AVSS.n103 185
R2873 AVSS.n102 AVSS.n101 185
R2874 AVSS.n100 AVSS.n99 185
R2875 AVSS.n98 AVSS.n97 185
R2876 AVSS.n96 AVSS.n95 185
R2877 AVSS.n94 AVSS.n93 185
R2878 AVSS.n92 AVSS.n91 185
R2879 AVSS.n90 AVSS.n89 185
R2880 AVSS.n88 AVSS.n87 185
R2881 AVSS.n59 AVSS.n57 185
R2882 AVSS.n145 AVSS.n144 185
R2883 AVSS.n4168 AVSS.n4167 185
R2884 AVSS.n4166 AVSS.n4165 185
R2885 AVSS.n4164 AVSS.n4163 185
R2886 AVSS.n4162 AVSS.n4161 185
R2887 AVSS.n4160 AVSS.n4159 185
R2888 AVSS.n4158 AVSS.n4157 185
R2889 AVSS.n4156 AVSS.n4155 185
R2890 AVSS.n4154 AVSS.n4153 185
R2891 AVSS.n4152 AVSS.n4151 185
R2892 AVSS.n4170 AVSS.n4169 185
R2893 AVSS.n4171 AVSS.n4124 185
R2894 AVSS.t101 AVSS.n4124 185
R2895 AVSS.n4173 AVSS.n4172 185
R2896 AVSS.n4175 AVSS.n4174 185
R2897 AVSS.n4177 AVSS.n4176 185
R2898 AVSS.n4179 AVSS.n4178 185
R2899 AVSS.n4181 AVSS.n4180 185
R2900 AVSS.n4183 AVSS.n4182 185
R2901 AVSS.n4185 AVSS.n4184 185
R2902 AVSS.n4116 AVSS.n4114 185
R2903 AVSS.n4200 AVSS.n4199 185
R2904 AVSS.n4198 AVSS.n4135 185
R2905 AVSS.n4197 AVSS.n4196 185
R2906 AVSS.n4195 AVSS.n4194 185
R2907 AVSS.n4193 AVSS.n4192 185
R2908 AVSS.n4191 AVSS.n4190 185
R2909 AVSS.n4189 AVSS.n4188 185
R2910 AVSS.n4187 AVSS.n4186 185
R2911 AVSS.n4150 AVSS.n4149 185
R2912 AVSS.n4148 AVSS.n4147 185
R2913 AVSS.n4146 AVSS.n4145 185
R2914 AVSS.n4144 AVSS.n4143 185
R2915 AVSS.n4142 AVSS.n4141 185
R2916 AVSS.n4140 AVSS.n4139 185
R2917 AVSS.n4138 AVSS.n4137 185
R2918 AVSS.n4117 AVSS.n4115 185
R2919 AVSS.n4203 AVSS.n4202 185
R2920 AVSS.n4202 AVSS.t101 185
R2921 AVSS.n4026 AVSS.n4025 185
R2922 AVSS.n4024 AVSS.n4007 185
R2923 AVSS.n4022 AVSS.n4021 185
R2924 AVSS.n4020 AVSS.n4008 185
R2925 AVSS.n4019 AVSS.n4018 185
R2926 AVSS.n4016 AVSS.n4009 185
R2927 AVSS.n4014 AVSS.n4013 185
R2928 AVSS.n4012 AVSS.n4011 185
R2929 AVSS.n3992 AVSS.n3990 185
R2930 AVSS.n4028 AVSS.n4027 185
R2931 AVSS.n4029 AVSS.n4005 185
R2932 AVSS.n4029 AVSS.t94 185
R2933 AVSS.n4032 AVSS.n4031 185
R2934 AVSS.n4033 AVSS.n4004 185
R2935 AVSS.n4035 AVSS.n4034 185
R2936 AVSS.n4037 AVSS.n4003 185
R2937 AVSS.n4040 AVSS.n4039 185
R2938 AVSS.n4041 AVSS.n4002 185
R2939 AVSS.n4043 AVSS.n4042 185
R2940 AVSS.n4061 AVSS.n4060 185
R2941 AVSS.n4058 AVSS.n3997 185
R2942 AVSS.n4057 AVSS.n4056 185
R2943 AVSS.n4055 AVSS.n4054 185
R2944 AVSS.n4053 AVSS.n3999 185
R2945 AVSS.n4051 AVSS.n4050 185
R2946 AVSS.n4049 AVSS.n4000 185
R2947 AVSS.n4048 AVSS.n4047 185
R2948 AVSS.n4045 AVSS.n4001 185
R2949 AVSS.n4079 AVSS.n4078 185
R2950 AVSS.n4076 AVSS.n3991 185
R2951 AVSS.n4075 AVSS.n3993 185
R2952 AVSS.n4073 AVSS.n4072 185
R2953 AVSS.n4071 AVSS.n3994 185
R2954 AVSS.n4070 AVSS.n4069 185
R2955 AVSS.n4067 AVSS.n3995 185
R2956 AVSS.n4065 AVSS.n4064 185
R2957 AVSS.n4063 AVSS.n3996 185
R2958 AVSS.n3996 AVSS.t94 185
R2959 AVSS.n3815 AVSS.n3814 185
R2960 AVSS.n3813 AVSS.n3796 185
R2961 AVSS.n3811 AVSS.n3810 185
R2962 AVSS.n3809 AVSS.n3797 185
R2963 AVSS.n3808 AVSS.n3807 185
R2964 AVSS.n3805 AVSS.n3798 185
R2965 AVSS.n3803 AVSS.n3802 185
R2966 AVSS.n3801 AVSS.n3800 185
R2967 AVSS.n3781 AVSS.n3779 185
R2968 AVSS.n3817 AVSS.n3816 185
R2969 AVSS.n3818 AVSS.n3794 185
R2970 AVSS.n3818 AVSS.t107 185
R2971 AVSS.n3821 AVSS.n3820 185
R2972 AVSS.n3822 AVSS.n3793 185
R2973 AVSS.n3824 AVSS.n3823 185
R2974 AVSS.n3826 AVSS.n3792 185
R2975 AVSS.n3829 AVSS.n3828 185
R2976 AVSS.n3830 AVSS.n3791 185
R2977 AVSS.n3832 AVSS.n3831 185
R2978 AVSS.n3850 AVSS.n3849 185
R2979 AVSS.n3847 AVSS.n3786 185
R2980 AVSS.n3846 AVSS.n3845 185
R2981 AVSS.n3844 AVSS.n3843 185
R2982 AVSS.n3842 AVSS.n3788 185
R2983 AVSS.n3840 AVSS.n3839 185
R2984 AVSS.n3838 AVSS.n3789 185
R2985 AVSS.n3837 AVSS.n3836 185
R2986 AVSS.n3834 AVSS.n3790 185
R2987 AVSS.n3868 AVSS.n3867 185
R2988 AVSS.n3865 AVSS.n3780 185
R2989 AVSS.n3864 AVSS.n3782 185
R2990 AVSS.n3862 AVSS.n3861 185
R2991 AVSS.n3860 AVSS.n3783 185
R2992 AVSS.n3859 AVSS.n3858 185
R2993 AVSS.n3856 AVSS.n3784 185
R2994 AVSS.n3854 AVSS.n3853 185
R2995 AVSS.n3852 AVSS.n3785 185
R2996 AVSS.n3785 AVSS.t107 185
R2997 AVSS.n3456 AVSS.n3455 185
R2998 AVSS.n3454 AVSS.n3437 185
R2999 AVSS.n3452 AVSS.n3451 185
R3000 AVSS.n3450 AVSS.n3438 185
R3001 AVSS.n3449 AVSS.n3448 185
R3002 AVSS.n3446 AVSS.n3439 185
R3003 AVSS.n3444 AVSS.n3443 185
R3004 AVSS.n3442 AVSS.n3441 185
R3005 AVSS.n3422 AVSS.n3420 185
R3006 AVSS.n3458 AVSS.n3457 185
R3007 AVSS.n3459 AVSS.n3435 185
R3008 AVSS.n3459 AVSS.t109 185
R3009 AVSS.n3462 AVSS.n3461 185
R3010 AVSS.n3463 AVSS.n3434 185
R3011 AVSS.n3465 AVSS.n3464 185
R3012 AVSS.n3467 AVSS.n3433 185
R3013 AVSS.n3470 AVSS.n3469 185
R3014 AVSS.n3471 AVSS.n3432 185
R3015 AVSS.n3473 AVSS.n3472 185
R3016 AVSS.n3491 AVSS.n3490 185
R3017 AVSS.n3488 AVSS.n3427 185
R3018 AVSS.n3487 AVSS.n3486 185
R3019 AVSS.n3485 AVSS.n3484 185
R3020 AVSS.n3483 AVSS.n3429 185
R3021 AVSS.n3481 AVSS.n3480 185
R3022 AVSS.n3479 AVSS.n3430 185
R3023 AVSS.n3478 AVSS.n3477 185
R3024 AVSS.n3475 AVSS.n3431 185
R3025 AVSS.n3508 AVSS.n3507 185
R3026 AVSS.n3505 AVSS.n3421 185
R3027 AVSS.n3504 AVSS.n3423 185
R3028 AVSS.n3502 AVSS.n3501 185
R3029 AVSS.n3500 AVSS.n3424 185
R3030 AVSS.n3499 AVSS.n3498 185
R3031 AVSS.n3496 AVSS.n3425 185
R3032 AVSS.n3494 AVSS.n3493 185
R3033 AVSS.n3492 AVSS.n3426 185
R3034 AVSS.n3426 AVSS.t109 185
R3035 AVSS.n5797 AVSS.n5746 185
R3036 AVSS.n5811 AVSS.n5810 185
R3037 AVSS.n5809 AVSS.n5747 185
R3038 AVSS.n5808 AVSS.n5807 185
R3039 AVSS.n5806 AVSS.n5805 185
R3040 AVSS.n5804 AVSS.n5803 185
R3041 AVSS.n5802 AVSS.n5801 185
R3042 AVSS.n5800 AVSS.n5799 185
R3043 AVSS.n5798 AVSS.n5727 185
R3044 AVSS.n5780 AVSS.n5779 185
R3045 AVSS.n5782 AVSS.n5781 185
R3046 AVSS.n5784 AVSS.n5783 185
R3047 AVSS.n5786 AVSS.n5785 185
R3048 AVSS.n5788 AVSS.n5787 185
R3049 AVSS.n5790 AVSS.n5789 185
R3050 AVSS.n5792 AVSS.n5791 185
R3051 AVSS.n5794 AVSS.n5793 185
R3052 AVSS.n5796 AVSS.n5795 185
R3053 AVSS.n5762 AVSS.n5761 185
R3054 AVSS.n5764 AVSS.n5763 185
R3055 AVSS.n5766 AVSS.n5765 185
R3056 AVSS.n5768 AVSS.n5767 185
R3057 AVSS.n5770 AVSS.n5769 185
R3058 AVSS.n5772 AVSS.n5771 185
R3059 AVSS.n5774 AVSS.n5773 185
R3060 AVSS.n5776 AVSS.n5775 185
R3061 AVSS.n5778 AVSS.n5777 185
R3062 AVSS.n5760 AVSS.n5759 185
R3063 AVSS.n5758 AVSS.n5757 185
R3064 AVSS.n5756 AVSS.n5755 185
R3065 AVSS.n5754 AVSS.n5753 185
R3066 AVSS.n5752 AVSS.n5751 185
R3067 AVSS.n5750 AVSS.n5749 185
R3068 AVSS.n5748 AVSS.n5730 185
R3069 AVSS.n5814 AVSS.n5728 185
R3070 AVSS.n5816 AVSS.n5815 185
R3071 AVSS.n5525 AVSS.n5474 185
R3072 AVSS.n5539 AVSS.n5538 185
R3073 AVSS.n5537 AVSS.n5475 185
R3074 AVSS.n5536 AVSS.n5535 185
R3075 AVSS.n5534 AVSS.n5533 185
R3076 AVSS.n5532 AVSS.n5531 185
R3077 AVSS.n5530 AVSS.n5529 185
R3078 AVSS.n5528 AVSS.n5527 185
R3079 AVSS.n5526 AVSS.n5455 185
R3080 AVSS.n5508 AVSS.n5507 185
R3081 AVSS.n5510 AVSS.n5509 185
R3082 AVSS.n5512 AVSS.n5511 185
R3083 AVSS.n5514 AVSS.n5513 185
R3084 AVSS.n5516 AVSS.n5515 185
R3085 AVSS.n5518 AVSS.n5517 185
R3086 AVSS.n5520 AVSS.n5519 185
R3087 AVSS.n5522 AVSS.n5521 185
R3088 AVSS.n5524 AVSS.n5523 185
R3089 AVSS.n5490 AVSS.n5489 185
R3090 AVSS.n5492 AVSS.n5491 185
R3091 AVSS.n5494 AVSS.n5493 185
R3092 AVSS.n5496 AVSS.n5495 185
R3093 AVSS.n5498 AVSS.n5497 185
R3094 AVSS.n5500 AVSS.n5499 185
R3095 AVSS.n5502 AVSS.n5501 185
R3096 AVSS.n5504 AVSS.n5503 185
R3097 AVSS.n5506 AVSS.n5505 185
R3098 AVSS.n5488 AVSS.n5487 185
R3099 AVSS.n5486 AVSS.n5485 185
R3100 AVSS.n5484 AVSS.n5483 185
R3101 AVSS.n5482 AVSS.n5481 185
R3102 AVSS.n5480 AVSS.n5479 185
R3103 AVSS.n5478 AVSS.n5477 185
R3104 AVSS.n5476 AVSS.n5458 185
R3105 AVSS.n5542 AVSS.n5456 185
R3106 AVSS.n5544 AVSS.n5543 185
R3107 AVSS.n5357 AVSS.n5356 185
R3108 AVSS.n5358 AVSS.n5311 185
R3109 AVSS.n5360 AVSS.n5359 185
R3110 AVSS.n5362 AVSS.n5310 185
R3111 AVSS.n5365 AVSS.n5364 185
R3112 AVSS.n5366 AVSS.n5309 185
R3113 AVSS.n5368 AVSS.n5367 185
R3114 AVSS.n5370 AVSS.n5308 185
R3115 AVSS.n5373 AVSS.n5372 185
R3116 AVSS.n5338 AVSS.n5316 185
R3117 AVSS.n5341 AVSS.n5340 185
R3118 AVSS.n5342 AVSS.n5315 185
R3119 AVSS.n5344 AVSS.n5343 185
R3120 AVSS.n5346 AVSS.n5314 185
R3121 AVSS.n5349 AVSS.n5348 185
R3122 AVSS.n5350 AVSS.n5313 185
R3123 AVSS.n5352 AVSS.n5351 185
R3124 AVSS.n5354 AVSS.n5312 185
R3125 AVSS.n5303 AVSS.n5301 185
R3126 AVSS.n5324 AVSS.n5321 185
R3127 AVSS.n5326 AVSS.n5325 185
R3128 AVSS.n5327 AVSS.n5320 185
R3129 AVSS.n5329 AVSS.n5328 185
R3130 AVSS.n5331 AVSS.n5318 185
R3131 AVSS.n5333 AVSS.n5332 185
R3132 AVSS.n5334 AVSS.n5317 185
R3133 AVSS.n5336 AVSS.n5335 185
R3134 AVSS.n5391 AVSS.n5390 185
R3135 AVSS.n5388 AVSS.n5302 185
R3136 AVSS.n5387 AVSS.n5304 185
R3137 AVSS.n5385 AVSS.n5384 185
R3138 AVSS.n5383 AVSS.n5305 185
R3139 AVSS.n5382 AVSS.n5381 185
R3140 AVSS.n5379 AVSS.n5306 185
R3141 AVSS.n5377 AVSS.n5376 185
R3142 AVSS.n5375 AVSS.n5307 185
R3143 AVSS.n5158 AVSS.n5157 185
R3144 AVSS.n5159 AVSS.n5112 185
R3145 AVSS.n5161 AVSS.n5160 185
R3146 AVSS.n5163 AVSS.n5111 185
R3147 AVSS.n5166 AVSS.n5165 185
R3148 AVSS.n5167 AVSS.n5110 185
R3149 AVSS.n5169 AVSS.n5168 185
R3150 AVSS.n5171 AVSS.n5109 185
R3151 AVSS.n5174 AVSS.n5173 185
R3152 AVSS.n5139 AVSS.n5117 185
R3153 AVSS.n5142 AVSS.n5141 185
R3154 AVSS.n5143 AVSS.n5116 185
R3155 AVSS.n5145 AVSS.n5144 185
R3156 AVSS.n5147 AVSS.n5115 185
R3157 AVSS.n5150 AVSS.n5149 185
R3158 AVSS.n5151 AVSS.n5114 185
R3159 AVSS.n5153 AVSS.n5152 185
R3160 AVSS.n5155 AVSS.n5113 185
R3161 AVSS.n5104 AVSS.n5102 185
R3162 AVSS.n5125 AVSS.n5122 185
R3163 AVSS.n5127 AVSS.n5126 185
R3164 AVSS.n5128 AVSS.n5121 185
R3165 AVSS.n5130 AVSS.n5129 185
R3166 AVSS.n5132 AVSS.n5119 185
R3167 AVSS.n5134 AVSS.n5133 185
R3168 AVSS.n5135 AVSS.n5118 185
R3169 AVSS.n5137 AVSS.n5136 185
R3170 AVSS.n5192 AVSS.n5191 185
R3171 AVSS.n5189 AVSS.n5103 185
R3172 AVSS.n5188 AVSS.n5105 185
R3173 AVSS.n5186 AVSS.n5185 185
R3174 AVSS.n5184 AVSS.n5106 185
R3175 AVSS.n5183 AVSS.n5182 185
R3176 AVSS.n5180 AVSS.n5107 185
R3177 AVSS.n5178 AVSS.n5177 185
R3178 AVSS.n5176 AVSS.n5108 185
R3179 AVSS.n465 AVSS.n462 185
R3180 AVSS.n486 AVSS.n485 185
R3181 AVSS.n488 AVSS.n487 185
R3182 AVSS.n490 AVSS.n489 185
R3183 AVSS.n492 AVSS.n491 185
R3184 AVSS.n494 AVSS.n493 185
R3185 AVSS.n496 AVSS.n495 185
R3186 AVSS.n498 AVSS.n497 185
R3187 AVSS.n500 AVSS.n499 185
R3188 AVSS.n501 AVSS.n469 185
R3189 AVSS.t103 AVSS.n469 185
R3190 AVSS.n503 AVSS.n502 185
R3191 AVSS.n505 AVSS.n504 185
R3192 AVSS.n507 AVSS.n506 185
R3193 AVSS.n509 AVSS.n508 185
R3194 AVSS.n511 AVSS.n510 185
R3195 AVSS.n513 AVSS.n512 185
R3196 AVSS.n514 AVSS.n482 185
R3197 AVSS.t103 AVSS.n482 185
R3198 AVSS.n516 AVSS.n515 185
R3199 AVSS.n518 AVSS.n517 185
R3200 AVSS.n520 AVSS.n519 185
R3201 AVSS.n522 AVSS.n521 185
R3202 AVSS.n524 AVSS.n523 185
R3203 AVSS.n526 AVSS.n525 185
R3204 AVSS.n528 AVSS.n527 185
R3205 AVSS.n530 AVSS.n529 185
R3206 AVSS.n532 AVSS.n531 185
R3207 AVSS.n533 AVSS.n484 185
R3208 AVSS.n550 AVSS.n549 185
R3209 AVSS.n464 AVSS.n463 185
R3210 AVSS.n535 AVSS.n534 185
R3211 AVSS.n537 AVSS.n536 185
R3212 AVSS.n539 AVSS.n538 185
R3213 AVSS.n541 AVSS.n540 185
R3214 AVSS.n543 AVSS.n542 185
R3215 AVSS.n544 AVSS.n483 185
R3216 AVSS.n546 AVSS.n545 185
R3217 AVSS.n1458 AVSS.n1457 185
R3218 AVSS.n1456 AVSS.n1455 185
R3219 AVSS.n1454 AVSS.n1453 185
R3220 AVSS.n1452 AVSS.n1451 185
R3221 AVSS.n1450 AVSS.n1449 185
R3222 AVSS.n1448 AVSS.n1447 185
R3223 AVSS.n1446 AVSS.n1445 185
R3224 AVSS.n1444 AVSS.n1443 185
R3225 AVSS.n1393 AVSS.n1390 185
R3226 AVSS.n1479 AVSS.n1478 185
R3227 AVSS.n1478 AVSS.t86 185
R3228 AVSS.n1392 AVSS.n1391 185
R3229 AVSS.n1414 AVSS.n1413 185
R3230 AVSS.n1416 AVSS.n1415 185
R3231 AVSS.n1418 AVSS.n1417 185
R3232 AVSS.n1420 AVSS.n1419 185
R3233 AVSS.n1422 AVSS.n1421 185
R3234 AVSS.n1423 AVSS.n1410 185
R3235 AVSS.t86 AVSS.n1410 185
R3236 AVSS.n1425 AVSS.n1424 185
R3237 AVSS.n1427 AVSS.n1426 185
R3238 AVSS.n1429 AVSS.n1428 185
R3239 AVSS.n1431 AVSS.n1430 185
R3240 AVSS.n1433 AVSS.n1432 185
R3241 AVSS.n1435 AVSS.n1434 185
R3242 AVSS.n1437 AVSS.n1436 185
R3243 AVSS.n1439 AVSS.n1438 185
R3244 AVSS.n1441 AVSS.n1440 185
R3245 AVSS.n1442 AVSS.n1412 185
R3246 AVSS.n1461 AVSS.n1460 185
R3247 AVSS.n1463 AVSS.n1462 185
R3248 AVSS.n1465 AVSS.n1464 185
R3249 AVSS.n1467 AVSS.n1466 185
R3250 AVSS.n1469 AVSS.n1468 185
R3251 AVSS.n1471 AVSS.n1470 185
R3252 AVSS.n1473 AVSS.n1472 185
R3253 AVSS.n1474 AVSS.n1411 185
R3254 AVSS.n1476 AVSS.n1475 185
R3255 AVSS.n4878 AVSS.n4877 185
R3256 AVSS.n4876 AVSS.n4875 185
R3257 AVSS.n4874 AVSS.n4873 185
R3258 AVSS.n4872 AVSS.n4871 185
R3259 AVSS.n4870 AVSS.n4869 185
R3260 AVSS.n4868 AVSS.n4867 185
R3261 AVSS.n4866 AVSS.n4865 185
R3262 AVSS.n4864 AVSS.n4863 185
R3263 AVSS.n4813 AVSS.n4810 185
R3264 AVSS.n4899 AVSS.n4898 185
R3265 AVSS.n4898 AVSS.t93 185
R3266 AVSS.n4812 AVSS.n4811 185
R3267 AVSS.n4834 AVSS.n4833 185
R3268 AVSS.n4836 AVSS.n4835 185
R3269 AVSS.n4838 AVSS.n4837 185
R3270 AVSS.n4840 AVSS.n4839 185
R3271 AVSS.n4842 AVSS.n4841 185
R3272 AVSS.n4843 AVSS.n4830 185
R3273 AVSS.t93 AVSS.n4830 185
R3274 AVSS.n4845 AVSS.n4844 185
R3275 AVSS.n4847 AVSS.n4846 185
R3276 AVSS.n4849 AVSS.n4848 185
R3277 AVSS.n4851 AVSS.n4850 185
R3278 AVSS.n4853 AVSS.n4852 185
R3279 AVSS.n4855 AVSS.n4854 185
R3280 AVSS.n4857 AVSS.n4856 185
R3281 AVSS.n4859 AVSS.n4858 185
R3282 AVSS.n4861 AVSS.n4860 185
R3283 AVSS.n4862 AVSS.n4832 185
R3284 AVSS.n4881 AVSS.n4880 185
R3285 AVSS.n4883 AVSS.n4882 185
R3286 AVSS.n4885 AVSS.n4884 185
R3287 AVSS.n4887 AVSS.n4886 185
R3288 AVSS.n4889 AVSS.n4888 185
R3289 AVSS.n4891 AVSS.n4890 185
R3290 AVSS.n4893 AVSS.n4892 185
R3291 AVSS.n4894 AVSS.n4831 185
R3292 AVSS.n4896 AVSS.n4895 185
R3293 AVSS.n3125 AVSS.n3123 185
R3294 AVSS.n3146 AVSS.n3145 185
R3295 AVSS.n3148 AVSS.n3147 185
R3296 AVSS.n3150 AVSS.n3149 185
R3297 AVSS.n3152 AVSS.n3151 185
R3298 AVSS.n3154 AVSS.n3153 185
R3299 AVSS.n3156 AVSS.n3155 185
R3300 AVSS.n3158 AVSS.n3157 185
R3301 AVSS.n3159 AVSS.n3143 185
R3302 AVSS.n3174 AVSS.n3173 185
R3303 AVSS.n3172 AVSS.n3171 185
R3304 AVSS.n3170 AVSS.n3169 185
R3305 AVSS.n3168 AVSS.n3167 185
R3306 AVSS.n3166 AVSS.n3165 185
R3307 AVSS.n3164 AVSS.n3163 185
R3308 AVSS.n3162 AVSS.n3161 185
R3309 AVSS.n3126 AVSS.n3124 185
R3310 AVSS.n3213 AVSS.n3212 185
R3311 AVSS.n3192 AVSS.n3191 185
R3312 AVSS.n3190 AVSS.n3189 185
R3313 AVSS.n3188 AVSS.n3187 185
R3314 AVSS.n3186 AVSS.n3185 185
R3315 AVSS.n3184 AVSS.n3183 185
R3316 AVSS.n3182 AVSS.n3181 185
R3317 AVSS.n3180 AVSS.n3179 185
R3318 AVSS.n3178 AVSS.n3177 185
R3319 AVSS.n3176 AVSS.n3175 185
R3320 AVSS.n3194 AVSS.n3193 185
R3321 AVSS.n3196 AVSS.n3195 185
R3322 AVSS.n3198 AVSS.n3197 185
R3323 AVSS.n3200 AVSS.n3199 185
R3324 AVSS.n3202 AVSS.n3201 185
R3325 AVSS.n3204 AVSS.n3203 185
R3326 AVSS.n3206 AVSS.n3205 185
R3327 AVSS.n3207 AVSS.n3144 185
R3328 AVSS.n3209 AVSS.n3208 185
R3329 AVSS.n1201 AVSS.n1199 185
R3330 AVSS.n1222 AVSS.n1221 185
R3331 AVSS.n1224 AVSS.n1223 185
R3332 AVSS.n1226 AVSS.n1225 185
R3333 AVSS.n1228 AVSS.n1227 185
R3334 AVSS.n1230 AVSS.n1229 185
R3335 AVSS.n1232 AVSS.n1231 185
R3336 AVSS.n1234 AVSS.n1233 185
R3337 AVSS.n1235 AVSS.n1219 185
R3338 AVSS.n1250 AVSS.n1249 185
R3339 AVSS.n1248 AVSS.n1247 185
R3340 AVSS.n1246 AVSS.n1245 185
R3341 AVSS.n1244 AVSS.n1243 185
R3342 AVSS.n1242 AVSS.n1241 185
R3343 AVSS.n1240 AVSS.n1239 185
R3344 AVSS.n1238 AVSS.n1237 185
R3345 AVSS.n1202 AVSS.n1200 185
R3346 AVSS.n1289 AVSS.n1288 185
R3347 AVSS.n1268 AVSS.n1267 185
R3348 AVSS.n1266 AVSS.n1265 185
R3349 AVSS.n1264 AVSS.n1263 185
R3350 AVSS.n1262 AVSS.n1261 185
R3351 AVSS.n1260 AVSS.n1259 185
R3352 AVSS.n1258 AVSS.n1257 185
R3353 AVSS.n1256 AVSS.n1255 185
R3354 AVSS.n1254 AVSS.n1253 185
R3355 AVSS.n1252 AVSS.n1251 185
R3356 AVSS.n1270 AVSS.n1269 185
R3357 AVSS.n1272 AVSS.n1271 185
R3358 AVSS.n1274 AVSS.n1273 185
R3359 AVSS.n1276 AVSS.n1275 185
R3360 AVSS.n1278 AVSS.n1277 185
R3361 AVSS.n1280 AVSS.n1279 185
R3362 AVSS.n1282 AVSS.n1281 185
R3363 AVSS.n1283 AVSS.n1220 185
R3364 AVSS.n1285 AVSS.n1284 185
R3365 AVSS.n4595 AVSS.n4543 185
R3366 AVSS.n4609 AVSS.n4608 185
R3367 AVSS.n4607 AVSS.n4544 185
R3368 AVSS.n4606 AVSS.n4605 185
R3369 AVSS.n4604 AVSS.n4603 185
R3370 AVSS.n4602 AVSS.n4601 185
R3371 AVSS.n4600 AVSS.n4599 185
R3372 AVSS.n4598 AVSS.n4597 185
R3373 AVSS.n4596 AVSS.n4524 185
R3374 AVSS.n4577 AVSS.n4576 185
R3375 AVSS.n4579 AVSS.n4578 185
R3376 AVSS.n4581 AVSS.n4580 185
R3377 AVSS.n4583 AVSS.n4582 185
R3378 AVSS.n4585 AVSS.n4584 185
R3379 AVSS.n4587 AVSS.n4586 185
R3380 AVSS.n4589 AVSS.n4588 185
R3381 AVSS.n4591 AVSS.n4590 185
R3382 AVSS.n4593 AVSS.n4592 185
R3383 AVSS.n4559 AVSS.n4558 185
R3384 AVSS.n4561 AVSS.n4560 185
R3385 AVSS.n4563 AVSS.n4562 185
R3386 AVSS.n4565 AVSS.n4564 185
R3387 AVSS.n4567 AVSS.n4566 185
R3388 AVSS.n4569 AVSS.n4568 185
R3389 AVSS.n4571 AVSS.n4570 185
R3390 AVSS.n4573 AVSS.n4572 185
R3391 AVSS.n4575 AVSS.n4574 185
R3392 AVSS.n4557 AVSS.n4556 185
R3393 AVSS.n4555 AVSS.n4554 185
R3394 AVSS.n4553 AVSS.n4552 185
R3395 AVSS.n4551 AVSS.n4550 185
R3396 AVSS.n4549 AVSS.n4548 185
R3397 AVSS.n4547 AVSS.n4546 185
R3398 AVSS.n4545 AVSS.n4527 185
R3399 AVSS.n4612 AVSS.n4525 185
R3400 AVSS.n4614 AVSS.n4613 185
R3401 AVSS.n2686 AVSS.n2684 185
R3402 AVSS.n2707 AVSS.n2706 185
R3403 AVSS.n2709 AVSS.n2708 185
R3404 AVSS.n2711 AVSS.n2710 185
R3405 AVSS.n2713 AVSS.n2712 185
R3406 AVSS.n2714 AVSS.n2705 185
R3407 AVSS.n2769 AVSS.n2768 185
R3408 AVSS.n2767 AVSS.n2704 185
R3409 AVSS.n2766 AVSS.n2765 185
R3410 AVSS.n2748 AVSS.n2747 185
R3411 AVSS.n2750 AVSS.n2749 185
R3412 AVSS.n2752 AVSS.n2751 185
R3413 AVSS.n2754 AVSS.n2753 185
R3414 AVSS.n2756 AVSS.n2755 185
R3415 AVSS.n2758 AVSS.n2757 185
R3416 AVSS.n2760 AVSS.n2759 185
R3417 AVSS.n2762 AVSS.n2761 185
R3418 AVSS.n2764 AVSS.n2763 185
R3419 AVSS.n2746 AVSS.n2745 185
R3420 AVSS.n2744 AVSS.n2743 185
R3421 AVSS.n2742 AVSS.n2741 185
R3422 AVSS.n2740 AVSS.n2739 185
R3423 AVSS.n2738 AVSS.n2737 185
R3424 AVSS.n2736 AVSS.n2735 185
R3425 AVSS.n2734 AVSS.n2733 185
R3426 AVSS.n2732 AVSS.n2731 185
R3427 AVSS.n2730 AVSS.n2729 185
R3428 AVSS.n2728 AVSS.n2727 185
R3429 AVSS.n2726 AVSS.n2725 185
R3430 AVSS.n2724 AVSS.n2723 185
R3431 AVSS.n2722 AVSS.n2721 185
R3432 AVSS.n2720 AVSS.n2719 185
R3433 AVSS.n2718 AVSS.n2717 185
R3434 AVSS.n2716 AVSS.n2715 185
R3435 AVSS.n2687 AVSS.n2685 185
R3436 AVSS.n2773 AVSS.n2772 185
R3437 AVSS.n2628 AVSS.n2627 185
R3438 AVSS.n2626 AVSS.n2609 185
R3439 AVSS.n2624 AVSS.n2623 185
R3440 AVSS.n2622 AVSS.n2610 185
R3441 AVSS.n2621 AVSS.n2620 185
R3442 AVSS.n2618 AVSS.n2611 185
R3443 AVSS.n2616 AVSS.n2615 185
R3444 AVSS.n2614 AVSS.n2613 185
R3445 AVSS.n2594 AVSS.n2592 185
R3446 AVSS.n2630 AVSS.n2629 185
R3447 AVSS.n2631 AVSS.n2607 185
R3448 AVSS.n2631 AVSS.t111 185
R3449 AVSS.n2634 AVSS.n2633 185
R3450 AVSS.n2635 AVSS.n2606 185
R3451 AVSS.n2637 AVSS.n2636 185
R3452 AVSS.n2639 AVSS.n2605 185
R3453 AVSS.n2642 AVSS.n2641 185
R3454 AVSS.n2643 AVSS.n2604 185
R3455 AVSS.n2645 AVSS.n2644 185
R3456 AVSS.n2663 AVSS.n2662 185
R3457 AVSS.n2660 AVSS.n2599 185
R3458 AVSS.n2659 AVSS.n2658 185
R3459 AVSS.n2657 AVSS.n2656 185
R3460 AVSS.n2655 AVSS.n2601 185
R3461 AVSS.n2653 AVSS.n2652 185
R3462 AVSS.n2651 AVSS.n2602 185
R3463 AVSS.n2650 AVSS.n2649 185
R3464 AVSS.n2647 AVSS.n2603 185
R3465 AVSS.n2681 AVSS.n2680 185
R3466 AVSS.n2678 AVSS.n2593 185
R3467 AVSS.n2677 AVSS.n2595 185
R3468 AVSS.n2675 AVSS.n2674 185
R3469 AVSS.n2673 AVSS.n2596 185
R3470 AVSS.n2672 AVSS.n2671 185
R3471 AVSS.n2669 AVSS.n2597 185
R3472 AVSS.n2667 AVSS.n2666 185
R3473 AVSS.n2665 AVSS.n2598 185
R3474 AVSS.n2598 AVSS.t111 185
R3475 AVSS.n1661 AVSS.n1660 185
R3476 AVSS.n1659 AVSS.n1642 185
R3477 AVSS.n1657 AVSS.n1656 185
R3478 AVSS.n1655 AVSS.n1643 185
R3479 AVSS.n1654 AVSS.n1653 185
R3480 AVSS.n1651 AVSS.n1644 185
R3481 AVSS.n1649 AVSS.n1648 185
R3482 AVSS.n1647 AVSS.n1646 185
R3483 AVSS.n1627 AVSS.n1625 185
R3484 AVSS.n1663 AVSS.n1662 185
R3485 AVSS.n1664 AVSS.n1640 185
R3486 AVSS.n1664 AVSS.t113 185
R3487 AVSS.n1667 AVSS.n1666 185
R3488 AVSS.n1668 AVSS.n1639 185
R3489 AVSS.n1670 AVSS.n1669 185
R3490 AVSS.n1672 AVSS.n1638 185
R3491 AVSS.n1675 AVSS.n1674 185
R3492 AVSS.n1676 AVSS.n1637 185
R3493 AVSS.n1678 AVSS.n1677 185
R3494 AVSS.n1696 AVSS.n1695 185
R3495 AVSS.n1693 AVSS.n1632 185
R3496 AVSS.n1692 AVSS.n1691 185
R3497 AVSS.n1690 AVSS.n1689 185
R3498 AVSS.n1688 AVSS.n1634 185
R3499 AVSS.n1686 AVSS.n1685 185
R3500 AVSS.n1684 AVSS.n1635 185
R3501 AVSS.n1683 AVSS.n1682 185
R3502 AVSS.n1680 AVSS.n1636 185
R3503 AVSS.n1713 AVSS.n1712 185
R3504 AVSS.n1710 AVSS.n1626 185
R3505 AVSS.n1709 AVSS.n1628 185
R3506 AVSS.n1707 AVSS.n1706 185
R3507 AVSS.n1705 AVSS.n1629 185
R3508 AVSS.n1704 AVSS.n1703 185
R3509 AVSS.n1701 AVSS.n1630 185
R3510 AVSS.n1699 AVSS.n1698 185
R3511 AVSS.n1697 AVSS.n1631 185
R3512 AVSS.n1631 AVSS.t113 185
R3513 AVSS.n2045 AVSS.n2044 185
R3514 AVSS.n2043 AVSS.n2042 185
R3515 AVSS.n2041 AVSS.n2040 185
R3516 AVSS.n2039 AVSS.n2038 185
R3517 AVSS.n2037 AVSS.n2036 185
R3518 AVSS.n2035 AVSS.n2034 185
R3519 AVSS.n2033 AVSS.n2032 185
R3520 AVSS.n2031 AVSS.n2030 185
R3521 AVSS.n1980 AVSS.n1977 185
R3522 AVSS.n2066 AVSS.n2065 185
R3523 AVSS.n2065 AVSS.t77 185
R3524 AVSS.n1979 AVSS.n1978 185
R3525 AVSS.n2001 AVSS.n2000 185
R3526 AVSS.n2003 AVSS.n2002 185
R3527 AVSS.n2005 AVSS.n2004 185
R3528 AVSS.n2007 AVSS.n2006 185
R3529 AVSS.n2009 AVSS.n2008 185
R3530 AVSS.n2010 AVSS.n1997 185
R3531 AVSS.t77 AVSS.n1997 185
R3532 AVSS.n2012 AVSS.n2011 185
R3533 AVSS.n2014 AVSS.n2013 185
R3534 AVSS.n2016 AVSS.n2015 185
R3535 AVSS.n2018 AVSS.n2017 185
R3536 AVSS.n2020 AVSS.n2019 185
R3537 AVSS.n2022 AVSS.n2021 185
R3538 AVSS.n2024 AVSS.n2023 185
R3539 AVSS.n2026 AVSS.n2025 185
R3540 AVSS.n2028 AVSS.n2027 185
R3541 AVSS.n2029 AVSS.n1999 185
R3542 AVSS.n2048 AVSS.n2047 185
R3543 AVSS.n2050 AVSS.n2049 185
R3544 AVSS.n2052 AVSS.n2051 185
R3545 AVSS.n2054 AVSS.n2053 185
R3546 AVSS.n2056 AVSS.n2055 185
R3547 AVSS.n2058 AVSS.n2057 185
R3548 AVSS.n2060 AVSS.n2059 185
R3549 AVSS.n2061 AVSS.n1998 185
R3550 AVSS.n2063 AVSS.n2062 185
R3551 AVSS.n742 AVSS.n740 185
R3552 AVSS.n763 AVSS.n762 185
R3553 AVSS.n765 AVSS.n764 185
R3554 AVSS.n767 AVSS.n766 185
R3555 AVSS.n769 AVSS.n768 185
R3556 AVSS.n771 AVSS.n770 185
R3557 AVSS.n773 AVSS.n772 185
R3558 AVSS.n775 AVSS.n774 185
R3559 AVSS.n776 AVSS.n760 185
R3560 AVSS.n791 AVSS.n790 185
R3561 AVSS.n789 AVSS.n788 185
R3562 AVSS.n787 AVSS.n786 185
R3563 AVSS.n785 AVSS.n784 185
R3564 AVSS.n783 AVSS.n782 185
R3565 AVSS.n781 AVSS.n780 185
R3566 AVSS.n779 AVSS.n778 185
R3567 AVSS.n743 AVSS.n741 185
R3568 AVSS.n830 AVSS.n829 185
R3569 AVSS.n809 AVSS.n808 185
R3570 AVSS.n807 AVSS.n806 185
R3571 AVSS.n805 AVSS.n804 185
R3572 AVSS.n803 AVSS.n802 185
R3573 AVSS.n801 AVSS.n800 185
R3574 AVSS.n799 AVSS.n798 185
R3575 AVSS.n797 AVSS.n796 185
R3576 AVSS.n795 AVSS.n794 185
R3577 AVSS.n793 AVSS.n792 185
R3578 AVSS.n811 AVSS.n810 185
R3579 AVSS.n813 AVSS.n812 185
R3580 AVSS.n815 AVSS.n814 185
R3581 AVSS.n817 AVSS.n816 185
R3582 AVSS.n819 AVSS.n818 185
R3583 AVSS.n821 AVSS.n820 185
R3584 AVSS.n823 AVSS.n822 185
R3585 AVSS.n824 AVSS.n761 185
R3586 AVSS.n826 AVSS.n825 185
R3587 AVSS.n1045 AVSS.n994 185
R3588 AVSS.n1059 AVSS.n1058 185
R3589 AVSS.n1057 AVSS.n995 185
R3590 AVSS.n1056 AVSS.n1055 185
R3591 AVSS.n1054 AVSS.n1053 185
R3592 AVSS.n1052 AVSS.n1051 185
R3593 AVSS.n1050 AVSS.n1049 185
R3594 AVSS.n1048 AVSS.n1047 185
R3595 AVSS.n1046 AVSS.n975 185
R3596 AVSS.n1028 AVSS.n1027 185
R3597 AVSS.n1030 AVSS.n1029 185
R3598 AVSS.n1032 AVSS.n1031 185
R3599 AVSS.n1034 AVSS.n1033 185
R3600 AVSS.n1036 AVSS.n1035 185
R3601 AVSS.n1038 AVSS.n1037 185
R3602 AVSS.n1040 AVSS.n1039 185
R3603 AVSS.n1042 AVSS.n1041 185
R3604 AVSS.n1044 AVSS.n1043 185
R3605 AVSS.n1010 AVSS.n1009 185
R3606 AVSS.n1012 AVSS.n1011 185
R3607 AVSS.n1014 AVSS.n1013 185
R3608 AVSS.n1016 AVSS.n1015 185
R3609 AVSS.n1018 AVSS.n1017 185
R3610 AVSS.n1020 AVSS.n1019 185
R3611 AVSS.n1022 AVSS.n1021 185
R3612 AVSS.n1024 AVSS.n1023 185
R3613 AVSS.n1026 AVSS.n1025 185
R3614 AVSS.n1008 AVSS.n1007 185
R3615 AVSS.n1006 AVSS.n1005 185
R3616 AVSS.n1004 AVSS.n1003 185
R3617 AVSS.n1002 AVSS.n1001 185
R3618 AVSS.n1000 AVSS.n999 185
R3619 AVSS.n998 AVSS.n997 185
R3620 AVSS.n996 AVSS.n978 185
R3621 AVSS.n1062 AVSS.n976 185
R3622 AVSS.n1064 AVSS.n1063 185
R3623 AVSS.n2490 AVSS.n2489 185
R3624 AVSS.n2491 AVSS.n2423 185
R3625 AVSS.n2493 AVSS.n2492 185
R3626 AVSS.n2495 AVSS.n2422 185
R3627 AVSS.n2498 AVSS.n2497 185
R3628 AVSS.n2499 AVSS.n2421 185
R3629 AVSS.n2501 AVSS.n2500 185
R3630 AVSS.n2503 AVSS.n2420 185
R3631 AVSS.n2504 AVSS.n2417 185
R3632 AVSS.n2471 AVSS.n2428 185
R3633 AVSS.n2474 AVSS.n2473 185
R3634 AVSS.n2475 AVSS.n2427 185
R3635 AVSS.n2477 AVSS.n2476 185
R3636 AVSS.n2479 AVSS.n2426 185
R3637 AVSS.n2482 AVSS.n2481 185
R3638 AVSS.n2483 AVSS.n2425 185
R3639 AVSS.n2485 AVSS.n2484 185
R3640 AVSS.n2487 AVSS.n2424 185
R3641 AVSS.n2455 AVSS.n2454 185
R3642 AVSS.n2457 AVSS.n2433 185
R3643 AVSS.n2459 AVSS.n2458 185
R3644 AVSS.n2460 AVSS.n2432 185
R3645 AVSS.n2462 AVSS.n2461 185
R3646 AVSS.n2464 AVSS.n2430 185
R3647 AVSS.n2466 AVSS.n2465 185
R3648 AVSS.n2467 AVSS.n2429 185
R3649 AVSS.n2469 AVSS.n2468 185
R3650 AVSS.n2452 AVSS.n2435 185
R3651 AVSS.n2451 AVSS.n2450 185
R3652 AVSS.n2448 AVSS.n2436 185
R3653 AVSS.n2446 AVSS.n2445 185
R3654 AVSS.n2444 AVSS.n2437 185
R3655 AVSS.n2443 AVSS.n2442 185
R3656 AVSS.n2440 AVSS.n2438 185
R3657 AVSS.n2419 AVSS.n2418 185
R3658 AVSS.n2507 AVSS.n2506 185
R3659 AVSS.n1889 AVSS.n1886 185
R3660 AVSS.n1910 AVSS.n1909 185
R3661 AVSS.n1912 AVSS.n1911 185
R3662 AVSS.n1914 AVSS.n1913 185
R3663 AVSS.n1916 AVSS.n1915 185
R3664 AVSS.n1918 AVSS.n1917 185
R3665 AVSS.n1920 AVSS.n1919 185
R3666 AVSS.n1922 AVSS.n1921 185
R3667 AVSS.n1924 AVSS.n1923 185
R3668 AVSS.n1925 AVSS.n1893 185
R3669 AVSS.t81 AVSS.n1893 185
R3670 AVSS.n1927 AVSS.n1926 185
R3671 AVSS.n1929 AVSS.n1928 185
R3672 AVSS.n1931 AVSS.n1930 185
R3673 AVSS.n1933 AVSS.n1932 185
R3674 AVSS.n1935 AVSS.n1934 185
R3675 AVSS.n1937 AVSS.n1936 185
R3676 AVSS.n1938 AVSS.n1906 185
R3677 AVSS.t81 AVSS.n1906 185
R3678 AVSS.n1940 AVSS.n1939 185
R3679 AVSS.n1942 AVSS.n1941 185
R3680 AVSS.n1944 AVSS.n1943 185
R3681 AVSS.n1946 AVSS.n1945 185
R3682 AVSS.n1948 AVSS.n1947 185
R3683 AVSS.n1950 AVSS.n1949 185
R3684 AVSS.n1952 AVSS.n1951 185
R3685 AVSS.n1954 AVSS.n1953 185
R3686 AVSS.n1956 AVSS.n1955 185
R3687 AVSS.n1957 AVSS.n1908 185
R3688 AVSS.n1974 AVSS.n1973 185
R3689 AVSS.n1888 AVSS.n1887 185
R3690 AVSS.n1959 AVSS.n1958 185
R3691 AVSS.n1961 AVSS.n1960 185
R3692 AVSS.n1963 AVSS.n1962 185
R3693 AVSS.n1965 AVSS.n1964 185
R3694 AVSS.n1967 AVSS.n1966 185
R3695 AVSS.n1968 AVSS.n1907 185
R3696 AVSS.n1970 AVSS.n1969 185
R3697 AVSS.n1787 AVSS.n1770 185
R3698 AVSS.n2555 AVSS.n2554 185
R3699 AVSS.n2553 AVSS.n1771 185
R3700 AVSS.n2552 AVSS.n2551 185
R3701 AVSS.n2550 AVSS.n2549 185
R3702 AVSS.n2548 AVSS.n2547 185
R3703 AVSS.n2546 AVSS.n2545 185
R3704 AVSS.n2544 AVSS.n2543 185
R3705 AVSS.n2542 AVSS.n2541 185
R3706 AVSS.n2559 AVSS.n2558 185
R3707 AVSS.n1752 AVSS.n1751 185
R3708 AVSS.n1773 AVSS.n1772 185
R3709 AVSS.n1775 AVSS.n1774 185
R3710 AVSS.n1777 AVSS.n1776 185
R3711 AVSS.n1779 AVSS.n1778 185
R3712 AVSS.n1781 AVSS.n1780 185
R3713 AVSS.n1783 AVSS.n1782 185
R3714 AVSS.n1785 AVSS.n1784 185
R3715 AVSS.n1804 AVSS.n1803 185
R3716 AVSS.n1802 AVSS.n1801 185
R3717 AVSS.n1800 AVSS.n1799 185
R3718 AVSS.n1798 AVSS.n1797 185
R3719 AVSS.n1796 AVSS.n1795 185
R3720 AVSS.n1794 AVSS.n1793 185
R3721 AVSS.n1792 AVSS.n1791 185
R3722 AVSS.n1790 AVSS.n1789 185
R3723 AVSS.n1753 AVSS.n1750 185
R3724 AVSS.n1806 AVSS.n1805 185
R3725 AVSS.n1808 AVSS.n1807 185
R3726 AVSS.n1810 AVSS.n1809 185
R3727 AVSS.n1812 AVSS.n1811 185
R3728 AVSS.n1814 AVSS.n1813 185
R3729 AVSS.n1816 AVSS.n1815 185
R3730 AVSS.n1818 AVSS.n1817 185
R3731 AVSS.n1820 AVSS.n1819 185
R3732 AVSS.n1822 AVSS.n1821 185
R3733 AVSS.n3307 AVSS.n3304 185
R3734 AVSS.n3328 AVSS.n3327 185
R3735 AVSS.n3330 AVSS.n3329 185
R3736 AVSS.n3332 AVSS.n3331 185
R3737 AVSS.n3334 AVSS.n3333 185
R3738 AVSS.n3336 AVSS.n3335 185
R3739 AVSS.n3338 AVSS.n3337 185
R3740 AVSS.n3340 AVSS.n3339 185
R3741 AVSS.n3342 AVSS.n3341 185
R3742 AVSS.n3344 AVSS.n3311 185
R3743 AVSS.t97 AVSS.n3311 185
R3744 AVSS.n3346 AVSS.n3345 185
R3745 AVSS.n3348 AVSS.n3347 185
R3746 AVSS.n3350 AVSS.n3349 185
R3747 AVSS.n3352 AVSS.n3351 185
R3748 AVSS.n3354 AVSS.n3353 185
R3749 AVSS.n3356 AVSS.n3355 185
R3750 AVSS.n3357 AVSS.n3324 185
R3751 AVSS.t97 AVSS.n3324 185
R3752 AVSS.n3359 AVSS.n3358 185
R3753 AVSS.n3361 AVSS.n3360 185
R3754 AVSS.n3363 AVSS.n3362 185
R3755 AVSS.n3365 AVSS.n3364 185
R3756 AVSS.n3367 AVSS.n3366 185
R3757 AVSS.n3369 AVSS.n3368 185
R3758 AVSS.n3371 AVSS.n3370 185
R3759 AVSS.n3373 AVSS.n3372 185
R3760 AVSS.n3375 AVSS.n3374 185
R3761 AVSS.n3376 AVSS.n3326 185
R3762 AVSS.n3393 AVSS.n3392 185
R3763 AVSS.n3306 AVSS.n3305 185
R3764 AVSS.n3378 AVSS.n3377 185
R3765 AVSS.n3380 AVSS.n3379 185
R3766 AVSS.n3382 AVSS.n3381 185
R3767 AVSS.n3384 AVSS.n3383 185
R3768 AVSS.n3386 AVSS.n3385 185
R3769 AVSS.n3387 AVSS.n3325 185
R3770 AVSS.n3389 AVSS.n3388 185
R3771 AVSS.n4926 AVSS.t78 183.917
R3772 AVSS.n2073 AVSS.t78 183.917
R3773 AVSS.n2582 AVSS.t78 183.917
R3774 AVSS.t78 AVSS.n1082 183.917
R3775 AVSS.n6187 AVSS.n160 175.546
R3776 AVSS.n6183 AVSS.n160 175.546
R3777 AVSS.n6183 AVSS.n163 175.546
R3778 AVSS.n6179 AVSS.n163 175.546
R3779 AVSS.n6179 AVSS.n165 175.546
R3780 AVSS.n6175 AVSS.n165 175.546
R3781 AVSS.n6175 AVSS.n170 175.546
R3782 AVSS.n6171 AVSS.n170 175.546
R3783 AVSS.n6171 AVSS.n172 175.546
R3784 AVSS.n6167 AVSS.n172 175.546
R3785 AVSS.n6167 AVSS.n174 175.546
R3786 AVSS.n6139 AVSS.n184 175.546
R3787 AVSS.n6143 AVSS.n184 175.546
R3788 AVSS.n6143 AVSS.n182 175.546
R3789 AVSS.n6147 AVSS.n182 175.546
R3790 AVSS.n6147 AVSS.n180 175.546
R3791 AVSS.n6151 AVSS.n180 175.546
R3792 AVSS.n6152 AVSS.n6151 175.546
R3793 AVSS.n6155 AVSS.n6152 175.546
R3794 AVSS.n6155 AVSS.n178 175.546
R3795 AVSS.n6159 AVSS.n178 175.546
R3796 AVSS.n6159 AVSS.n176 175.546
R3797 AVSS.n6163 AVSS.n176 175.546
R3798 AVSS.n259 AVSS.n255 175.546
R3799 AVSS.n253 AVSS.n234 175.546
R3800 AVSS.n249 AVSS.n247 175.546
R3801 AVSS.n245 AVSS.n236 175.546
R3802 AVSS.n241 AVSS.n239 175.546
R3803 AVSS.n6208 AVSS.n6207 175.546
R3804 AVSS.n6205 AVSS.n152 175.546
R3805 AVSS.n6201 AVSS.n6200 175.546
R3806 AVSS.n6198 AVSS.n155 175.546
R3807 AVSS.n6194 AVSS.n6193 175.546
R3808 AVSS.n6191 AVSS.n158 175.546
R3809 AVSS.n1194 AVSS.n1167 175.546
R3810 AVSS.n1190 AVSS.n1172 175.546
R3811 AVSS.n1186 AVSS.n1185 175.546
R3812 AVSS.n1182 AVSS.n1181 175.546
R3813 AVSS.n1178 AVSS.n1177 175.546
R3814 AVSS.n1299 AVSS.n1297 175.546
R3815 AVSS.n1303 AVSS.n1163 175.546
R3816 AVSS.n1307 AVSS.n1305 175.546
R3817 AVSS.n1311 AVSS.n1161 175.546
R3818 AVSS.n1314 AVSS.n1313 175.546
R3819 AVSS.n1318 AVSS.n1317 175.546
R3820 AVSS.n1321 AVSS.n1157 175.546
R3821 AVSS.n1325 AVSS.n1157 175.546
R3822 AVSS.n1325 AVSS.n1155 175.546
R3823 AVSS.n1330 AVSS.n1155 175.546
R3824 AVSS.n1330 AVSS.n1153 175.546
R3825 AVSS.n1334 AVSS.n1153 175.546
R3826 AVSS.n1335 AVSS.n1334 175.546
R3827 AVSS.n1337 AVSS.n1335 175.546
R3828 AVSS.n1337 AVSS.n1151 175.546
R3829 AVSS.n1342 AVSS.n1151 175.546
R3830 AVSS.n1342 AVSS.n1149 175.546
R3831 AVSS.n1367 AVSS.n1146 175.546
R3832 AVSS.n1363 AVSS.n1362 175.546
R3833 AVSS.n1359 AVSS.n1358 175.546
R3834 AVSS.n1355 AVSS.n1354 175.546
R3835 AVSS.n1351 AVSS.n1350 175.546
R3836 AVSS.n1347 AVSS.n1346 175.546
R3837 AVSS.n4629 AVSS.n4627 175.546
R3838 AVSS.n4633 AVSS.n4622 175.546
R3839 AVSS.n4637 AVSS.n4635 175.546
R3840 AVSS.n4641 AVSS.n4620 175.546
R3841 AVSS.n4644 AVSS.n4643 175.546
R3842 AVSS.n4979 AVSS.n1070 175.546
R3843 AVSS.n4977 AVSS.n4976 175.546
R3844 AVSS.n4974 AVSS.n1073 175.546
R3845 AVSS.n4970 AVSS.n4969 175.546
R3846 AVSS.n4967 AVSS.n1076 175.546
R3847 AVSS.n4963 AVSS.n4962 175.546
R3848 AVSS.n4956 AVSS.n4955 175.546
R3849 AVSS.n4953 AVSS.n1083 175.546
R3850 AVSS.n4949 AVSS.n4948 175.546
R3851 AVSS.n4946 AVSS.n1086 175.546
R3852 AVSS.n4942 AVSS.n4941 175.546
R3853 AVSS.n4665 AVSS.n1126 175.546
R3854 AVSS.n4663 AVSS.n4662 175.546
R3855 AVSS.n4659 AVSS.n4658 175.546
R3856 AVSS.n4655 AVSS.n4654 175.546
R3857 AVSS.n4651 AVSS.n4650 175.546
R3858 AVSS.n4935 AVSS.n1091 175.546
R3859 AVSS.n2119 AVSS.n2117 175.546
R3860 AVSS.n2123 AVSS.n2087 175.546
R3861 AVSS.n2127 AVSS.n2125 175.546
R3862 AVSS.n2131 AVSS.n2085 175.546
R3863 AVSS.n2134 AVSS.n2133 175.546
R3864 AVSS.n2111 AVSS.n2089 175.546
R3865 AVSS.n2109 AVSS.n2108 175.546
R3866 AVSS.n2106 AVSS.n2092 175.546
R3867 AVSS.n2102 AVSS.n2101 175.546
R3868 AVSS.n2099 AVSS.n2096 175.546
R3869 AVSS.n2187 AVSS.n2071 175.546
R3870 AVSS.n2182 AVSS.n2074 175.546
R3871 AVSS.n2178 AVSS.n2177 175.546
R3872 AVSS.n2175 AVSS.n2077 175.546
R3873 AVSS.n2171 AVSS.n2170 175.546
R3874 AVSS.n2168 AVSS.n2080 175.546
R3875 AVSS.n2139 AVSS.n1139 175.546
R3876 AVSS.n2143 AVSS.n2142 175.546
R3877 AVSS.n2147 AVSS.n2146 175.546
R3878 AVSS.n2151 AVSS.n2150 175.546
R3879 AVSS.n2155 AVSS.n2154 175.546
R3880 AVSS.n2159 AVSS.n2158 175.546
R3881 AVSS.n837 AVSS.n836 175.546
R3882 AVSS.n841 AVSS.n840 175.546
R3883 AVSS.n845 AVSS.n844 175.546
R3884 AVSS.n849 AVSS.n848 175.546
R3885 AVSS.n853 AVSS.n852 175.546
R3886 AVSS.n857 AVSS.n682 175.546
R3887 AVSS.n861 AVSS.n681 175.546
R3888 AVSS.n861 AVSS.n679 175.546
R3889 AVSS.n866 AVSS.n679 175.546
R3890 AVSS.n866 AVSS.n677 175.546
R3891 AVSS.n870 AVSS.n677 175.546
R3892 AVSS.n872 AVSS.n870 175.546
R3893 AVSS.n872 AVSS.n675 175.546
R3894 AVSS.n876 AVSS.n675 175.546
R3895 AVSS.n876 AVSS.n673 175.546
R3896 AVSS.n880 AVSS.n673 175.546
R3897 AVSS.n880 AVSS.n670 175.546
R3898 AVSS.n735 AVSS.n734 175.546
R3899 AVSS.n731 AVSS.n730 175.546
R3900 AVSS.n727 AVSS.n726 175.546
R3901 AVSS.n723 AVSS.n722 175.546
R3902 AVSS.n719 AVSS.n718 175.546
R3903 AVSS.n884 AVSS.n669 175.546
R3904 AVSS.n696 AVSS.n689 175.546
R3905 AVSS.n700 AVSS.n698 175.546
R3906 AVSS.n704 AVSS.n687 175.546
R3907 AVSS.n708 AVSS.n706 175.546
R3908 AVSS.n712 AVSS.n685 175.546
R3909 AVSS.n5571 AVSS.n5277 175.546
R3910 AVSS.n5575 AVSS.n5277 175.546
R3911 AVSS.n5575 AVSS.n5275 175.546
R3912 AVSS.n5579 AVSS.n5275 175.546
R3913 AVSS.n5579 AVSS.n5273 175.546
R3914 AVSS.n5583 AVSS.n5273 175.546
R3915 AVSS.n5583 AVSS.n5271 175.546
R3916 AVSS.n5587 AVSS.n5271 175.546
R3917 AVSS.n5587 AVSS.n5269 175.546
R3918 AVSS.n5591 AVSS.n5269 175.546
R3919 AVSS.n5591 AVSS.n5266 175.546
R3920 AVSS.n5615 AVSS.n5266 175.546
R3921 AVSS.n5611 AVSS.n5610 175.546
R3922 AVSS.n5607 AVSS.n5606 175.546
R3923 AVSS.n5603 AVSS.n5602 175.546
R3924 AVSS.n5599 AVSS.n5598 175.546
R3925 AVSS.n5595 AVSS.n5259 175.546
R3926 AVSS.n5872 AVSS.n5256 175.546
R3927 AVSS.n5868 AVSS.n5867 175.546
R3928 AVSS.n5864 AVSS.n5863 175.546
R3929 AVSS.n5860 AVSS.n5859 175.546
R3930 AVSS.n5856 AVSS.n5855 175.546
R3931 AVSS.n5852 AVSS.n5851 175.546
R3932 AVSS.n5567 AVSS.n5449 175.546
R3933 AVSS.n5563 AVSS.n5454 175.546
R3934 AVSS.n5559 AVSS.n5558 175.546
R3935 AVSS.n5555 AVSS.n5554 175.546
R3936 AVSS.n5551 AVSS.n5550 175.546
R3937 AVSS.n6275 AVSS.n11 175.546
R3938 AVSS.n6275 AVSS.n13 175.546
R3939 AVSS.n6271 AVSS.n13 175.546
R3940 AVSS.n6271 AVSS.n16 175.546
R3941 AVSS.n6267 AVSS.n16 175.546
R3942 AVSS.n6267 AVSS.n18 175.546
R3943 AVSS.n5285 AVSS.n18 175.546
R3944 AVSS.n5288 AVSS.n5285 175.546
R3945 AVSS.n5288 AVSS.n5283 175.546
R3946 AVSS.n5292 AVSS.n5283 175.546
R3947 AVSS.n5292 AVSS.n5280 175.546
R3948 AVSS.n5444 AVSS.n5280 175.546
R3949 AVSS.n6283 AVSS.n6281 175.546
R3950 AVSS.n6287 AVSS.n9 175.546
R3951 AVSS.n6291 AVSS.n6289 175.546
R3952 AVSS.n6295 AVSS.n7 175.546
R3953 AVSS.n6298 AVSS.n6297 175.546
R3954 AVSS.n5396 AVSS.n4 175.546
R3955 AVSS.n5400 AVSS.n5399 175.546
R3956 AVSS.n5404 AVSS.n5403 175.546
R3957 AVSS.n5408 AVSS.n5407 175.546
R3958 AVSS.n5412 AVSS.n5411 175.546
R3959 AVSS.n5416 AVSS.n5415 175.546
R3960 AVSS.n5440 AVSS.n5438 175.546
R3961 AVSS.n5436 AVSS.n5296 175.546
R3962 AVSS.n5432 AVSS.n5430 175.546
R3963 AVSS.n5428 AVSS.n5298 175.546
R3964 AVSS.n5424 AVSS.n5422 175.546
R3965 AVSS.n5074 AVSS.n428 175.546
R3966 AVSS.n5074 AVSS.n430 175.546
R3967 AVSS.n5070 AVSS.n430 175.546
R3968 AVSS.n5070 AVSS.n433 175.546
R3969 AVSS.n5066 AVSS.n433 175.546
R3970 AVSS.n5066 AVSS.n435 175.546
R3971 AVSS.n446 AVSS.n435 175.546
R3972 AVSS.n446 AVSS.n437 175.546
R3973 AVSS.n442 AVSS.n437 175.546
R3974 AVSS.n442 AVSS.n439 175.546
R3975 AVSS.n439 AVSS.n417 175.546
R3976 AVSS.n5218 AVSS.n417 175.546
R3977 AVSS.n5089 AVSS.n427 175.546
R3978 AVSS.n5087 AVSS.n5086 175.546
R3979 AVSS.n5083 AVSS.n5082 175.546
R3980 AVSS.n5079 AVSS.n5078 175.546
R3981 AVSS.n5097 AVSS.n422 175.546
R3982 AVSS.n5248 AVSS.n407 175.546
R3983 AVSS.n5244 AVSS.n5243 175.546
R3984 AVSS.n5240 AVSS.n5239 175.546
R3985 AVSS.n5236 AVSS.n5235 175.546
R3986 AVSS.n5232 AVSS.n5231 175.546
R3987 AVSS.n5228 AVSS.n5227 175.546
R3988 AVSS.n5214 AVSS.n5213 175.546
R3989 AVSS.n5210 AVSS.n5209 175.546
R3990 AVSS.n5206 AVSS.n5205 175.546
R3991 AVSS.n5202 AVSS.n5201 175.546
R3992 AVSS.n5198 AVSS.n410 175.546
R3993 AVSS.n5924 AVSS.n301 175.546
R3994 AVSS.n5920 AVSS.n301 175.546
R3995 AVSS.n5920 AVSS.n304 175.546
R3996 AVSS.n5916 AVSS.n304 175.546
R3997 AVSS.n5916 AVSS.n306 175.546
R3998 AVSS.n5912 AVSS.n306 175.546
R3999 AVSS.n5912 AVSS.n308 175.546
R4000 AVSS.n5908 AVSS.n308 175.546
R4001 AVSS.n5908 AVSS.n310 175.546
R4002 AVSS.n5904 AVSS.n310 175.546
R4003 AVSS.n5904 AVSS.n312 175.546
R4004 AVSS.n5900 AVSS.n312 175.546
R4005 AVSS.n357 AVSS.n300 175.546
R4006 AVSS.n357 AVSS.n355 175.546
R4007 AVSS.n361 AVSS.n355 175.546
R4008 AVSS.n361 AVSS.n353 175.546
R4009 AVSS.n365 AVSS.n353 175.546
R4010 AVSS.n365 AVSS.n351 175.546
R4011 AVSS.n369 AVSS.n351 175.546
R4012 AVSS.n369 AVSS.n349 175.546
R4013 AVSS.n373 AVSS.n349 175.546
R4014 AVSS.n373 AVSS.n347 175.546
R4015 AVSS.n397 AVSS.n347 175.546
R4016 AVSS.n393 AVSS.n340 175.546
R4017 AVSS.n391 AVSS.n390 175.546
R4018 AVSS.n387 AVSS.n386 175.546
R4019 AVSS.n383 AVSS.n382 175.546
R4020 AVSS.n379 AVSS.n378 175.546
R4021 AVSS.n5875 AVSS.n327 175.546
R4022 AVSS.n5896 AVSS.n5895 175.546
R4023 AVSS.n5893 AVSS.n318 175.546
R4024 AVSS.n5889 AVSS.n5888 175.546
R4025 AVSS.n5886 AVSS.n321 175.546
R4026 AVSS.n5882 AVSS.n5881 175.546
R4027 AVSS.n5651 AVSS.n5624 175.546
R4028 AVSS.n5655 AVSS.n5651 175.546
R4029 AVSS.n5655 AVSS.n5649 175.546
R4030 AVSS.n5659 AVSS.n5649 175.546
R4031 AVSS.n5660 AVSS.n5659 175.546
R4032 AVSS.n5660 AVSS.n5647 175.546
R4033 AVSS.n5664 AVSS.n5647 175.546
R4034 AVSS.n5664 AVSS.n5646 175.546
R4035 AVSS.n5668 AVSS.n5646 175.546
R4036 AVSS.n5668 AVSS.n5644 175.546
R4037 AVSS.n5672 AVSS.n5644 175.546
R4038 AVSS.n5672 AVSS.n5642 175.546
R4039 AVSS.n5676 AVSS.n5640 175.546
R4040 AVSS.n5680 AVSS.n5640 175.546
R4041 AVSS.n5680 AVSS.n5638 175.546
R4042 AVSS.n5685 AVSS.n5638 175.546
R4043 AVSS.n5685 AVSS.n5636 175.546
R4044 AVSS.n5689 AVSS.n5636 175.546
R4045 AVSS.n5689 AVSS.n5635 175.546
R4046 AVSS.n5693 AVSS.n5635 175.546
R4047 AVSS.n5693 AVSS.n5633 175.546
R4048 AVSS.n5698 AVSS.n5633 175.546
R4049 AVSS.n5698 AVSS.n5631 175.546
R4050 AVSS.n5723 AVSS.n5722 175.546
R4051 AVSS.n5719 AVSS.n5718 175.546
R4052 AVSS.n5715 AVSS.n5714 175.546
R4053 AVSS.n5711 AVSS.n5710 175.546
R4054 AVSS.n5707 AVSS.n5706 175.546
R4055 AVSS.n5703 AVSS.n5702 175.546
R4056 AVSS.n5837 AVSS.n5623 175.546
R4057 AVSS.n5835 AVSS.n5834 175.546
R4058 AVSS.n5831 AVSS.n5830 175.546
R4059 AVSS.n5827 AVSS.n5826 175.546
R4060 AVSS.n5823 AVSS.n5822 175.546
R4061 AVSS.n2275 AVSS.n606 175.546
R4062 AVSS.n2273 AVSS.n2272 175.546
R4063 AVSS.n2269 AVSS.n2268 175.546
R4064 AVSS.n2265 AVSS.n2264 175.546
R4065 AVSS.n2261 AVSS.n2260 175.546
R4066 AVSS.n2257 AVSS.n2256 175.546
R4067 AVSS.n2250 AVSS.n2202 175.546
R4068 AVSS.n2246 AVSS.n2245 175.546
R4069 AVSS.n2243 AVSS.n2205 175.546
R4070 AVSS.n2239 AVSS.n2238 175.546
R4071 AVSS.n2236 AVSS.n2208 175.546
R4072 AVSS.n4987 AVSS.n972 175.546
R4073 AVSS.n2211 AVSS.n2210 175.546
R4074 AVSS.n2215 AVSS.n2214 175.546
R4075 AVSS.n2219 AVSS.n2218 175.546
R4076 AVSS.n2223 AVSS.n2222 175.546
R4077 AVSS.n2227 AVSS.n2226 175.546
R4078 AVSS.n2283 AVSS.n2281 175.546
R4079 AVSS.n2287 AVSS.n2199 175.546
R4080 AVSS.n2291 AVSS.n2289 175.546
R4081 AVSS.n2295 AVSS.n2197 175.546
R4082 AVSS.n2299 AVSS.n2297 175.546
R4083 AVSS.n2365 AVSS.n626 175.546
R4084 AVSS.n2369 AVSS.n2368 175.546
R4085 AVSS.n2373 AVSS.n2372 175.546
R4086 AVSS.n2377 AVSS.n2376 175.546
R4087 AVSS.n2381 AVSS.n2380 175.546
R4088 AVSS.n2385 AVSS.n2384 175.546
R4089 AVSS.n2394 AVSS.n2309 175.546
R4090 AVSS.n2398 AVSS.n2396 175.546
R4091 AVSS.n2402 AVSS.n2307 175.546
R4092 AVSS.n2405 AVSS.n2404 175.546
R4093 AVSS.n2409 AVSS.n2408 175.546
R4094 AVSS.n2336 AVSS.n654 175.546
R4095 AVSS.n2334 AVSS.n2333 175.546
R4096 AVSS.n2330 AVSS.n2329 175.546
R4097 AVSS.n2326 AVSS.n2325 175.546
R4098 AVSS.n2322 AVSS.n2321 175.546
R4099 AVSS.n2318 AVSS.n2317 175.546
R4100 AVSS.n2360 AVSS.n2359 175.546
R4101 AVSS.n2356 AVSS.n2355 175.546
R4102 AVSS.n2353 AVSS.n2313 175.546
R4103 AVSS.n2349 AVSS.n2347 175.546
R4104 AVSS.n2345 AVSS.n2315 175.546
R4105 AVSS.n1540 AVSS.n613 175.546
R4106 AVSS.n1544 AVSS.n1543 175.546
R4107 AVSS.n1548 AVSS.n1547 175.546
R4108 AVSS.n1552 AVSS.n1551 175.546
R4109 AVSS.n1556 AVSS.n1555 175.546
R4110 AVSS.n1560 AVSS.n1559 175.546
R4111 AVSS.n1537 AVSS.n1485 175.546
R4112 AVSS.n1533 AVSS.n1485 175.546
R4113 AVSS.n1533 AVSS.n1487 175.546
R4114 AVSS.n1529 AVSS.n1487 175.546
R4115 AVSS.n1529 AVSS.n1526 175.546
R4116 AVSS.n1526 AVSS.n1525 175.546
R4117 AVSS.n1525 AVSS.n1489 175.546
R4118 AVSS.n1521 AVSS.n1489 175.546
R4119 AVSS.n1521 AVSS.n1492 175.546
R4120 AVSS.n1517 AVSS.n1492 175.546
R4121 AVSS.n1517 AVSS.n1514 175.546
R4122 AVSS.n1510 AVSS.n661 175.546
R4123 AVSS.n1508 AVSS.n1507 175.546
R4124 AVSS.n1504 AVSS.n1503 175.546
R4125 AVSS.n1500 AVSS.n1499 175.546
R4126 AVSS.n1496 AVSS.n1495 175.546
R4127 AVSS.n1591 AVSS.n1590 175.546
R4128 AVSS.n1569 AVSS.n1389 175.546
R4129 AVSS.n1573 AVSS.n1571 175.546
R4130 AVSS.n1577 AVSS.n1387 175.546
R4131 AVSS.n1581 AVSS.n1579 175.546
R4132 AVSS.n1585 AVSS.n1385 175.546
R4133 AVSS.n5011 AVSS.n5010 175.546
R4134 AVSS.n5008 AVSS.n638 175.546
R4135 AVSS.n5004 AVSS.n5003 175.546
R4136 AVSS.n5001 AVSS.n641 175.546
R4137 AVSS.n4997 AVSS.n4996 175.546
R4138 AVSS.n964 AVSS.n893 175.546
R4139 AVSS.n960 AVSS.n959 175.546
R4140 AVSS.n956 AVSS.n955 175.546
R4141 AVSS.n952 AVSS.n951 175.546
R4142 AVSS.n948 AVSS.n947 175.546
R4143 AVSS.n4990 AVSS.n647 175.546
R4144 AVSS.n926 AVSS.n924 175.546
R4145 AVSS.n930 AVSS.n897 175.546
R4146 AVSS.n934 AVSS.n932 175.546
R4147 AVSS.n938 AVSS.n895 175.546
R4148 AVSS.n942 AVSS.n940 175.546
R4149 AVSS.n918 AVSS.n917 175.546
R4150 AVSS.n914 AVSS.n913 175.546
R4151 AVSS.n910 AVSS.n909 175.546
R4152 AVSS.n906 AVSS.n905 175.546
R4153 AVSS.n902 AVSS.n901 175.546
R4154 AVSS.n5015 AVSS.n633 175.546
R4155 AVSS.n3223 AVSS.n3221 175.546
R4156 AVSS.n3227 AVSS.n3089 175.546
R4157 AVSS.n3231 AVSS.n3229 175.546
R4158 AVSS.n3235 AVSS.n3087 175.546
R4159 AVSS.n3238 AVSS.n3237 175.546
R4160 AVSS.n3242 AVSS.n3241 175.546
R4161 AVSS.n3245 AVSS.n3083 175.546
R4162 AVSS.n3249 AVSS.n3083 175.546
R4163 AVSS.n3249 AVSS.n3081 175.546
R4164 AVSS.n3254 AVSS.n3081 175.546
R4165 AVSS.n3254 AVSS.n3079 175.546
R4166 AVSS.n3258 AVSS.n3079 175.546
R4167 AVSS.n3258 AVSS.n3078 175.546
R4168 AVSS.n3262 AVSS.n3078 175.546
R4169 AVSS.n3262 AVSS.n3076 175.546
R4170 AVSS.n3267 AVSS.n3076 175.546
R4171 AVSS.n3267 AVSS.n3074 175.546
R4172 AVSS.n3292 AVSS.n3071 175.546
R4173 AVSS.n3288 AVSS.n3287 175.546
R4174 AVSS.n3284 AVSS.n3283 175.546
R4175 AVSS.n3280 AVSS.n3279 175.546
R4176 AVSS.n3276 AVSS.n3275 175.546
R4177 AVSS.n3272 AVSS.n3271 175.546
R4178 AVSS.n3119 AVSS.n3117 175.546
R4179 AVSS.n3115 AVSS.n3093 175.546
R4180 AVSS.n3111 AVSS.n3109 175.546
R4181 AVSS.n3107 AVSS.n3095 175.546
R4182 AVSS.n3103 AVSS.n3101 175.546
R4183 AVSS.n4673 AVSS.n2780 175.546
R4184 AVSS.n4521 AVSS.n4520 175.546
R4185 AVSS.n4518 AVSS.n2783 175.546
R4186 AVSS.n4514 AVSS.n4513 175.546
R4187 AVSS.n4511 AVSS.n2786 175.546
R4188 AVSS.n4507 AVSS.n4506 175.546
R4189 AVSS.n4676 AVSS.n2778 175.546
R4190 AVSS.n2845 AVSS.n2842 175.546
R4191 AVSS.n2849 AVSS.n2847 175.546
R4192 AVSS.n2853 AVSS.n2839 175.546
R4193 AVSS.n2856 AVSS.n2855 175.546
R4194 AVSS.n2861 AVSS.n2829 175.546
R4195 AVSS.n2865 AVSS.n2864 175.546
R4196 AVSS.n2869 AVSS.n2868 175.546
R4197 AVSS.n2873 AVSS.n2872 175.546
R4198 AVSS.n2877 AVSS.n2876 175.546
R4199 AVSS.n2879 AVSS.n2835 175.546
R4200 AVSS.n4500 AVSS.n2791 175.546
R4201 AVSS.n2884 AVSS.n2883 175.546
R4202 AVSS.n2888 AVSS.n2887 175.546
R4203 AVSS.n2892 AVSS.n2891 175.546
R4204 AVSS.n2896 AVSS.n2895 175.546
R4205 AVSS.n4705 AVSS.n1727 175.546
R4206 AVSS.n4701 AVSS.n4700 175.546
R4207 AVSS.n4698 AVSS.n1730 175.546
R4208 AVSS.n4694 AVSS.n4693 175.546
R4209 AVSS.n4691 AVSS.n1733 175.546
R4210 AVSS.n4687 AVSS.n4686 175.546
R4211 AVSS.n4708 AVSS.n1725 175.546
R4212 AVSS.n2998 AVSS.n2995 175.546
R4213 AVSS.n3002 AVSS.n3000 175.546
R4214 AVSS.n3006 AVSS.n2992 175.546
R4215 AVSS.n3010 AVSS.n3008 175.546
R4216 AVSS.n3064 AVSS.n2990 175.546
R4217 AVSS.n3060 AVSS.n3059 175.546
R4218 AVSS.n3056 AVSS.n3055 175.546
R4219 AVSS.n3052 AVSS.n3051 175.546
R4220 AVSS.n3048 AVSS.n3047 175.546
R4221 AVSS.n3044 AVSS.n3043 175.546
R4222 AVSS.n3021 AVSS.n3019 175.546
R4223 AVSS.n3025 AVSS.n3023 175.546
R4224 AVSS.n3029 AVSS.n3016 175.546
R4225 AVSS.n3033 AVSS.n3031 175.546
R4226 AVSS.n3037 AVSS.n3014 175.546
R4227 AVSS.n2938 AVSS.n2937 175.546
R4228 AVSS.n2935 AVSS.n2916 175.546
R4229 AVSS.n2931 AVSS.n2930 175.546
R4230 AVSS.n2928 AVSS.n2919 175.546
R4231 AVSS.n2924 AVSS.n2923 175.546
R4232 AVSS.n4718 AVSS.n1718 175.546
R4233 AVSS.n2944 AVSS.n2913 175.546
R4234 AVSS.n2948 AVSS.n2946 175.546
R4235 AVSS.n2952 AVSS.n2911 175.546
R4236 AVSS.n2955 AVSS.n2954 175.546
R4237 AVSS.n2959 AVSS.n2958 175.546
R4238 AVSS.n2964 AVSS.n2902 175.546
R4239 AVSS.n2968 AVSS.n2967 175.546
R4240 AVSS.n2972 AVSS.n2971 175.546
R4241 AVSS.n2976 AVSS.n2975 175.546
R4242 AVSS.n2980 AVSS.n2907 175.546
R4243 AVSS.n4470 AVSS.n2828 175.546
R4244 AVSS.n2810 AVSS.n2809 175.546
R4245 AVSS.n2814 AVSS.n2813 175.546
R4246 AVSS.n2818 AVSS.n2817 175.546
R4247 AVSS.n2822 AVSS.n2821 175.546
R4248 AVSS.n2824 AVSS.n2807 175.546
R4249 AVSS.n4762 AVSS.n4759 175.546
R4250 AVSS.n4762 AVSS.n4732 175.546
R4251 AVSS.n4767 AVSS.n4732 175.546
R4252 AVSS.n4767 AVSS.n4729 175.546
R4253 AVSS.n4771 AVSS.n4729 175.546
R4254 AVSS.n4772 AVSS.n4771 175.546
R4255 AVSS.n4775 AVSS.n4772 175.546
R4256 AVSS.n4775 AVSS.n4727 175.546
R4257 AVSS.n4780 AVSS.n4727 175.546
R4258 AVSS.n4780 AVSS.n4725 175.546
R4259 AVSS.n4784 AVSS.n4725 175.546
R4260 AVSS.n4758 AVSS.n4734 175.546
R4261 AVSS.n4754 AVSS.n4753 175.546
R4262 AVSS.n4751 AVSS.n4737 175.546
R4263 AVSS.n4747 AVSS.n4746 175.546
R4264 AVSS.n4744 AVSS.n4741 175.546
R4265 AVSS.n4905 AVSS.n1380 175.546
R4266 AVSS.n4912 AVSS.n4911 175.546
R4267 AVSS.n4916 AVSS.n4915 175.546
R4268 AVSS.n4920 AVSS.n4919 175.546
R4269 AVSS.n4924 AVSS.n1378 175.546
R4270 AVSS.n4928 AVSS.n1373 175.546
R4271 AVSS.n4789 AVSS.n4788 175.546
R4272 AVSS.n4793 AVSS.n4792 175.546
R4273 AVSS.n4797 AVSS.n4796 175.546
R4274 AVSS.n4801 AVSS.n4800 175.546
R4275 AVSS.n4805 AVSS.n4804 175.546
R4276 AVSS.n4932 AVSS.n1369 175.546
R4277 AVSS.n2565 AVSS.n2564 175.546
R4278 AVSS.n2569 AVSS.n2568 175.546
R4279 AVSS.n2573 AVSS.n2572 175.546
R4280 AVSS.n2575 AVSS.n1746 175.546
R4281 AVSS.n2580 AVSS.n1741 175.546
R4282 AVSS.n1842 AVSS.n1841 175.546
R4283 AVSS.n1838 AVSS.n1837 175.546
R4284 AVSS.n1834 AVSS.n1833 175.546
R4285 AVSS.n1830 AVSS.n1829 175.546
R4286 AVSS.n1826 AVSS.n1825 175.546
R4287 AVSS.n2587 AVSS.n1119 175.546
R4288 AVSS.n2519 AVSS.n2517 175.546
R4289 AVSS.n2523 AVSS.n1851 175.546
R4290 AVSS.n2527 AVSS.n2525 175.546
R4291 AVSS.n2531 AVSS.n1849 175.546
R4292 AVSS.n2534 AVSS.n2533 175.546
R4293 AVSS.n1884 AVSS.n1882 175.546
R4294 AVSS.n1880 AVSS.n1855 175.546
R4295 AVSS.n1876 AVSS.n1874 175.546
R4296 AVSS.n1872 AVSS.n1857 175.546
R4297 AVSS.n1868 AVSS.n1866 175.546
R4298 AVSS.n1864 AVSS.n1860 175.546
R4299 AVSS.n4292 AVSS.n3892 175.546
R4300 AVSS.n4288 AVSS.n4287 175.546
R4301 AVSS.n4285 AVSS.n3895 175.546
R4302 AVSS.n4281 AVSS.n4280 175.546
R4303 AVSS.n4278 AVSS.n3898 175.546
R4304 AVSS.n4274 AVSS.n4273 175.546
R4305 AVSS.n4295 AVSS.n3891 175.546
R4306 AVSS.n3927 AVSS.n3924 175.546
R4307 AVSS.n3931 AVSS.n3929 175.546
R4308 AVSS.n3935 AVSS.n3921 175.546
R4309 AVSS.n3938 AVSS.n3937 175.546
R4310 AVSS.n3944 AVSS.n3918 175.546
R4311 AVSS.n3944 AVSS.n3917 175.546
R4312 AVSS.n3948 AVSS.n3917 175.546
R4313 AVSS.n3948 AVSS.n3915 175.546
R4314 AVSS.n3952 AVSS.n3915 175.546
R4315 AVSS.n3952 AVSS.n3913 175.546
R4316 AVSS.n3956 AVSS.n3913 175.546
R4317 AVSS.n3956 AVSS.n3911 175.546
R4318 AVSS.n3960 AVSS.n3911 175.546
R4319 AVSS.n3960 AVSS.n3909 175.546
R4320 AVSS.n3964 AVSS.n3909 175.546
R4321 AVSS.n3964 AVSS.n3907 175.546
R4322 AVSS.n3988 AVSS.n3986 175.546
R4323 AVSS.n3984 AVSS.n3903 175.546
R4324 AVSS.n3980 AVSS.n3978 175.546
R4325 AVSS.n3976 AVSS.n3905 175.546
R4326 AVSS.n3972 AVSS.n3970 175.546
R4327 AVSS.n4325 AVSS.n3681 175.546
R4328 AVSS.n4321 AVSS.n4320 175.546
R4329 AVSS.n4318 AVSS.n3684 175.546
R4330 AVSS.n4314 AVSS.n4313 175.546
R4331 AVSS.n4311 AVSS.n3687 175.546
R4332 AVSS.n4307 AVSS.n4306 175.546
R4333 AVSS.n4328 AVSS.n3680 175.546
R4334 AVSS.n3716 AVSS.n3713 175.546
R4335 AVSS.n3720 AVSS.n3718 175.546
R4336 AVSS.n3724 AVSS.n3710 175.546
R4337 AVSS.n3727 AVSS.n3726 175.546
R4338 AVSS.n3733 AVSS.n3707 175.546
R4339 AVSS.n3733 AVSS.n3706 175.546
R4340 AVSS.n3737 AVSS.n3706 175.546
R4341 AVSS.n3737 AVSS.n3704 175.546
R4342 AVSS.n3741 AVSS.n3704 175.546
R4343 AVSS.n3741 AVSS.n3702 175.546
R4344 AVSS.n3745 AVSS.n3702 175.546
R4345 AVSS.n3745 AVSS.n3700 175.546
R4346 AVSS.n3749 AVSS.n3700 175.546
R4347 AVSS.n3749 AVSS.n3698 175.546
R4348 AVSS.n3753 AVSS.n3698 175.546
R4349 AVSS.n3753 AVSS.n3696 175.546
R4350 AVSS.n3777 AVSS.n3775 175.546
R4351 AVSS.n3773 AVSS.n3692 175.546
R4352 AVSS.n3769 AVSS.n3767 175.546
R4353 AVSS.n3765 AVSS.n3694 175.546
R4354 AVSS.n3761 AVSS.n3759 175.546
R4355 AVSS.n3560 AVSS.n3559 175.546
R4356 AVSS.n3557 AVSS.n3538 175.546
R4357 AVSS.n3553 AVSS.n3552 175.546
R4358 AVSS.n3550 AVSS.n3541 175.546
R4359 AVSS.n3546 AVSS.n3545 175.546
R4360 AVSS.n4339 AVSS.n3513 175.546
R4361 AVSS.n3562 AVSS.n3535 175.546
R4362 AVSS.n3566 AVSS.n3535 175.546
R4363 AVSS.n3566 AVSS.n3533 175.546
R4364 AVSS.n3570 AVSS.n3533 175.546
R4365 AVSS.n3570 AVSS.n3530 175.546
R4366 AVSS.n3604 AVSS.n3530 175.546
R4367 AVSS.n3604 AVSS.n3531 175.546
R4368 AVSS.n3600 AVSS.n3531 175.546
R4369 AVSS.n3600 AVSS.n3574 175.546
R4370 AVSS.n3596 AVSS.n3574 175.546
R4371 AVSS.n3596 AVSS.n3576 175.546
R4372 AVSS.n3592 AVSS.n3578 175.546
R4373 AVSS.n3588 AVSS.n3578 175.546
R4374 AVSS.n3588 AVSS.n3580 175.546
R4375 AVSS.n3584 AVSS.n3580 175.546
R4376 AVSS.n3584 AVSS.n3582 175.546
R4377 AVSS.n3582 AVSS.n3526 175.546
R4378 AVSS.n3608 AVSS.n3526 175.546
R4379 AVSS.n3608 AVSS.n3524 175.546
R4380 AVSS.n3612 AVSS.n3524 175.546
R4381 AVSS.n3612 AVSS.n3522 175.546
R4382 AVSS.n3616 AVSS.n3522 175.546
R4383 AVSS.n3616 AVSS.n3520 175.546
R4384 AVSS.n3639 AVSS.n3638 175.546
R4385 AVSS.n3636 AVSS.n3516 175.546
R4386 AVSS.n3632 AVSS.n3630 175.546
R4387 AVSS.n3628 AVSS.n3518 175.546
R4388 AVSS.n3624 AVSS.n3622 175.546
R4389 AVSS.n6092 AVSS.n6090 175.546
R4390 AVSS.n6096 AVSS.n227 175.546
R4391 AVSS.n6100 AVSS.n6098 175.546
R4392 AVSS.n6104 AVSS.n225 175.546
R4393 AVSS.n6108 AVSS.n6106 175.546
R4394 AVSS.n6136 AVSS.n212 175.546
R4395 AVSS.n6132 AVSS.n212 175.546
R4396 AVSS.n6132 AVSS.n215 175.546
R4397 AVSS.n6128 AVSS.n215 175.546
R4398 AVSS.n6128 AVSS.n217 175.546
R4399 AVSS.n6124 AVSS.n217 175.546
R4400 AVSS.n6124 AVSS.n219 175.546
R4401 AVSS.n6120 AVSS.n219 175.546
R4402 AVSS.n6120 AVSS.n221 175.546
R4403 AVSS.n6116 AVSS.n221 175.546
R4404 AVSS.n6116 AVSS.n6113 175.546
R4405 AVSS.n6113 AVSS.n6112 175.546
R4406 AVSS.n4262 AVSS.n4229 175.546
R4407 AVSS.n4227 AVSS.n4208 175.546
R4408 AVSS.n4223 AVSS.n4221 175.546
R4409 AVSS.n4219 AVSS.n4210 175.546
R4410 AVSS.n4215 AVSS.n4213 175.546
R4411 AVSS.n4256 AVSS.n4255 175.546
R4412 AVSS.n4253 AVSS.n4232 175.546
R4413 AVSS.n4249 AVSS.n4247 175.546
R4414 AVSS.n4245 AVSS.n4234 175.546
R4415 AVSS.n4241 AVSS.n4239 175.546
R4416 AVSS.n4237 AVSS.n229 175.546
R4417 AVSS.n4395 AVSS.n4393 175.546
R4418 AVSS.n4399 AVSS.n4357 175.546
R4419 AVSS.n4403 AVSS.n4401 175.546
R4420 AVSS.n4407 AVSS.n4355 175.546
R4421 AVSS.n4411 AVSS.n4409 175.546
R4422 AVSS.n4416 AVSS.n4353 175.546
R4423 AVSS.n4424 AVSS.n4351 175.546
R4424 AVSS.n4428 AVSS.n4426 175.546
R4425 AVSS.n4432 AVSS.n4349 175.546
R4426 AVSS.n4436 AVSS.n4434 175.546
R4427 AVSS.n4440 AVSS.n4347 175.546
R4428 AVSS.n4467 AVSS.n3301 175.546
R4429 AVSS.n4463 AVSS.n4462 175.546
R4430 AVSS.n4459 AVSS.n4458 175.546
R4431 AVSS.n4455 AVSS.n4454 175.546
R4432 AVSS.n4451 AVSS.n4450 175.546
R4433 AVSS.n4447 AVSS.n4446 175.546
R4434 AVSS.n4392 AVSS.n4359 175.546
R4435 AVSS.n4388 AVSS.n4359 175.546
R4436 AVSS.n4388 AVSS.n4362 175.546
R4437 AVSS.n4384 AVSS.n4362 175.546
R4438 AVSS.n4384 AVSS.n4381 175.546
R4439 AVSS.n4381 AVSS.n4380 175.546
R4440 AVSS.n4380 AVSS.n4365 175.546
R4441 AVSS.n4376 AVSS.n4365 175.546
R4442 AVSS.n4376 AVSS.n4368 175.546
R4443 AVSS.n4372 AVSS.n4368 175.546
R4444 AVSS.n4372 AVSS.n3300 175.546
R4445 AVSS.n5911 AVSS.n5910 167.617
R4446 AVSS.n5065 AVSS.t99 163.958
R4447 AVSS.n6266 AVSS.t89 163.958
R4448 AVSS.t92 AVSS.n5581 163.958
R4449 AVSS.t106 AVSS.n36 163.958
R4450 AVSS.n4151 AVSS.n4150 163.333
R4451 AVSS.n4078 AVSS.n3992 163.333
R4452 AVSS.n3867 AVSS.n3781 163.333
R4453 AVSS.n3507 AVSS.n3422 163.333
R4454 AVSS.n499 AVSS.n469 163.333
R4455 AVSS.n1478 AVSS.n1393 163.333
R4456 AVSS.n4898 AVSS.n4813 163.333
R4457 AVSS.n2680 AVSS.n2594 163.333
R4458 AVSS.n1712 AVSS.n1627 163.333
R4459 AVSS.n2065 AVSS.n1980 163.333
R4460 AVSS.n1923 AVSS.n1893 163.333
R4461 AVSS.n3341 AVSS.n3311 163.333
R4462 AVSS.n87 AVSS.n59 150
R4463 AVSS.n91 AVSS.n90 150
R4464 AVSS.n95 AVSS.n94 150
R4465 AVSS.n99 AVSS.n98 150
R4466 AVSS.n103 AVSS.n102 150
R4467 AVSS.n107 AVSS.n106 150
R4468 AVSS.n111 AVSS.n110 150
R4469 AVSS.n115 AVSS.n114 150
R4470 AVSS.n135 AVSS.n134 150
R4471 AVSS.n131 AVSS.n130 150
R4472 AVSS.n127 AVSS.n126 150
R4473 AVSS.n123 AVSS.n122 150
R4474 AVSS.n80 AVSS.n79 150
R4475 AVSS.n84 AVSS.n83 150
R4476 AVSS.n141 AVSS.n77 150
R4477 AVSS.n137 AVSS.n76 150
R4478 AVSS.n4155 AVSS.n4154 150
R4479 AVSS.n4159 AVSS.n4158 150
R4480 AVSS.n4163 AVSS.n4162 150
R4481 AVSS.n4167 AVSS.n4166 150
R4482 AVSS.n4184 AVSS.n4183 150
R4483 AVSS.n4180 AVSS.n4179 150
R4484 AVSS.n4176 AVSS.n4175 150
R4485 AVSS.n4172 AVSS.n4124 150
R4486 AVSS.n4169 AVSS.n4124 150
R4487 AVSS.n4200 AVSS.n4135 150
R4488 AVSS.n4196 AVSS.n4195 150
R4489 AVSS.n4192 AVSS.n4191 150
R4490 AVSS.n4188 AVSS.n4187 150
R4491 AVSS.n4202 AVSS.n4117 150
R4492 AVSS.n4139 AVSS.n4138 150
R4493 AVSS.n4143 AVSS.n4142 150
R4494 AVSS.n4147 AVSS.n4146 150
R4495 AVSS.n4014 AVSS.n4011 150
R4496 AVSS.n4018 AVSS.n4016 150
R4497 AVSS.n4022 AVSS.n4008 150
R4498 AVSS.n4025 AVSS.n4024 150
R4499 AVSS.n4043 AVSS.n4002 150
R4500 AVSS.n4039 AVSS.n4037 150
R4501 AVSS.n4035 AVSS.n4004 150
R4502 AVSS.n4031 AVSS.n4029 150
R4503 AVSS.n4029 AVSS.n4028 150
R4504 AVSS.n4058 AVSS.n4057 150
R4505 AVSS.n4054 AVSS.n4053 150
R4506 AVSS.n4051 AVSS.n4000 150
R4507 AVSS.n4047 AVSS.n4045 150
R4508 AVSS.n4065 AVSS.n3996 150
R4509 AVSS.n4069 AVSS.n4067 150
R4510 AVSS.n4073 AVSS.n3994 150
R4511 AVSS.n4076 AVSS.n4075 150
R4512 AVSS.n3803 AVSS.n3800 150
R4513 AVSS.n3807 AVSS.n3805 150
R4514 AVSS.n3811 AVSS.n3797 150
R4515 AVSS.n3814 AVSS.n3813 150
R4516 AVSS.n3832 AVSS.n3791 150
R4517 AVSS.n3828 AVSS.n3826 150
R4518 AVSS.n3824 AVSS.n3793 150
R4519 AVSS.n3820 AVSS.n3818 150
R4520 AVSS.n3818 AVSS.n3817 150
R4521 AVSS.n3847 AVSS.n3846 150
R4522 AVSS.n3843 AVSS.n3842 150
R4523 AVSS.n3840 AVSS.n3789 150
R4524 AVSS.n3836 AVSS.n3834 150
R4525 AVSS.n3854 AVSS.n3785 150
R4526 AVSS.n3858 AVSS.n3856 150
R4527 AVSS.n3862 AVSS.n3783 150
R4528 AVSS.n3865 AVSS.n3864 150
R4529 AVSS.n3494 AVSS.n3426 150
R4530 AVSS.n3498 AVSS.n3496 150
R4531 AVSS.n3502 AVSS.n3424 150
R4532 AVSS.n3505 AVSS.n3504 150
R4533 AVSS.n3488 AVSS.n3487 150
R4534 AVSS.n3484 AVSS.n3483 150
R4535 AVSS.n3481 AVSS.n3430 150
R4536 AVSS.n3477 AVSS.n3475 150
R4537 AVSS.n3473 AVSS.n3432 150
R4538 AVSS.n3469 AVSS.n3467 150
R4539 AVSS.n3465 AVSS.n3434 150
R4540 AVSS.n3461 AVSS.n3459 150
R4541 AVSS.n3459 AVSS.n3458 150
R4542 AVSS.n3444 AVSS.n3441 150
R4543 AVSS.n3448 AVSS.n3446 150
R4544 AVSS.n3452 AVSS.n3438 150
R4545 AVSS.n3455 AVSS.n3454 150
R4546 AVSS.n5793 AVSS.n5792 150
R4547 AVSS.n5789 AVSS.n5788 150
R4548 AVSS.n5785 AVSS.n5784 150
R4549 AVSS.n5781 AVSS.n5780 150
R4550 AVSS.n5777 AVSS.n5776 150
R4551 AVSS.n5773 AVSS.n5772 150
R4552 AVSS.n5769 AVSS.n5768 150
R4553 AVSS.n5765 AVSS.n5764 150
R4554 AVSS.n5815 AVSS.n5814 150
R4555 AVSS.n5749 AVSS.n5730 150
R4556 AVSS.n5753 AVSS.n5752 150
R4557 AVSS.n5757 AVSS.n5756 150
R4558 AVSS.n5811 AVSS.n5747 150
R4559 AVSS.n5807 AVSS.n5806 150
R4560 AVSS.n5803 AVSS.n5802 150
R4561 AVSS.n5799 AVSS.n5798 150
R4562 AVSS.n5521 AVSS.n5520 150
R4563 AVSS.n5517 AVSS.n5516 150
R4564 AVSS.n5513 AVSS.n5512 150
R4565 AVSS.n5509 AVSS.n5508 150
R4566 AVSS.n5505 AVSS.n5504 150
R4567 AVSS.n5501 AVSS.n5500 150
R4568 AVSS.n5497 AVSS.n5496 150
R4569 AVSS.n5493 AVSS.n5492 150
R4570 AVSS.n5543 AVSS.n5542 150
R4571 AVSS.n5477 AVSS.n5458 150
R4572 AVSS.n5481 AVSS.n5480 150
R4573 AVSS.n5485 AVSS.n5484 150
R4574 AVSS.n5539 AVSS.n5475 150
R4575 AVSS.n5535 AVSS.n5534 150
R4576 AVSS.n5531 AVSS.n5530 150
R4577 AVSS.n5527 AVSS.n5526 150
R4578 AVSS.n5360 AVSS.n5311 150
R4579 AVSS.n5364 AVSS.n5362 150
R4580 AVSS.n5368 AVSS.n5309 150
R4581 AVSS.n5372 AVSS.n5370 150
R4582 AVSS.n5352 AVSS.n5313 150
R4583 AVSS.n5348 AVSS.n5346 150
R4584 AVSS.n5344 AVSS.n5315 150
R4585 AVSS.n5340 AVSS.n5338 150
R4586 AVSS.n5336 AVSS.n5317 150
R4587 AVSS.n5332 AVSS.n5331 150
R4588 AVSS.n5329 AVSS.n5320 150
R4589 AVSS.n5325 AVSS.n5324 150
R4590 AVSS.n5377 AVSS.n5307 150
R4591 AVSS.n5381 AVSS.n5379 150
R4592 AVSS.n5385 AVSS.n5305 150
R4593 AVSS.n5388 AVSS.n5387 150
R4594 AVSS.n5161 AVSS.n5112 150
R4595 AVSS.n5165 AVSS.n5163 150
R4596 AVSS.n5169 AVSS.n5110 150
R4597 AVSS.n5173 AVSS.n5171 150
R4598 AVSS.n5153 AVSS.n5114 150
R4599 AVSS.n5149 AVSS.n5147 150
R4600 AVSS.n5145 AVSS.n5116 150
R4601 AVSS.n5141 AVSS.n5139 150
R4602 AVSS.n5137 AVSS.n5118 150
R4603 AVSS.n5133 AVSS.n5132 150
R4604 AVSS.n5130 AVSS.n5121 150
R4605 AVSS.n5126 AVSS.n5125 150
R4606 AVSS.n5178 AVSS.n5108 150
R4607 AVSS.n5182 AVSS.n5180 150
R4608 AVSS.n5186 AVSS.n5106 150
R4609 AVSS.n5189 AVSS.n5188 150
R4610 AVSS.n515 AVSS.n482 150
R4611 AVSS.n512 AVSS.n482 150
R4612 AVSS.n510 AVSS.n509 150
R4613 AVSS.n506 AVSS.n505 150
R4614 AVSS.n502 AVSS.n469 150
R4615 AVSS.n519 AVSS.n518 150
R4616 AVSS.n523 AVSS.n522 150
R4617 AVSS.n527 AVSS.n526 150
R4618 AVSS.n531 AVSS.n530 150
R4619 AVSS.n542 AVSS.n483 150
R4620 AVSS.n540 AVSS.n539 150
R4621 AVSS.n536 AVSS.n535 150
R4622 AVSS.n549 AVSS.n464 150
R4623 AVSS.n497 AVSS.n496 150
R4624 AVSS.n493 AVSS.n492 150
R4625 AVSS.n489 AVSS.n488 150
R4626 AVSS.n485 AVSS.n465 150
R4627 AVSS.n1445 AVSS.n1444 150
R4628 AVSS.n1449 AVSS.n1448 150
R4629 AVSS.n1453 AVSS.n1452 150
R4630 AVSS.n1457 AVSS.n1456 150
R4631 AVSS.n1472 AVSS.n1411 150
R4632 AVSS.n1470 AVSS.n1469 150
R4633 AVSS.n1466 AVSS.n1465 150
R4634 AVSS.n1462 AVSS.n1461 150
R4635 AVSS.n1428 AVSS.n1427 150
R4636 AVSS.n1432 AVSS.n1431 150
R4637 AVSS.n1436 AVSS.n1435 150
R4638 AVSS.n1440 AVSS.n1439 150
R4639 AVSS.n1424 AVSS.n1410 150
R4640 AVSS.n1421 AVSS.n1410 150
R4641 AVSS.n1419 AVSS.n1418 150
R4642 AVSS.n1415 AVSS.n1414 150
R4643 AVSS.n1478 AVSS.n1392 150
R4644 AVSS.n4865 AVSS.n4864 150
R4645 AVSS.n4869 AVSS.n4868 150
R4646 AVSS.n4873 AVSS.n4872 150
R4647 AVSS.n4877 AVSS.n4876 150
R4648 AVSS.n4892 AVSS.n4831 150
R4649 AVSS.n4890 AVSS.n4889 150
R4650 AVSS.n4886 AVSS.n4885 150
R4651 AVSS.n4882 AVSS.n4881 150
R4652 AVSS.n4848 AVSS.n4847 150
R4653 AVSS.n4852 AVSS.n4851 150
R4654 AVSS.n4856 AVSS.n4855 150
R4655 AVSS.n4860 AVSS.n4859 150
R4656 AVSS.n4844 AVSS.n4830 150
R4657 AVSS.n4841 AVSS.n4830 150
R4658 AVSS.n4839 AVSS.n4838 150
R4659 AVSS.n4835 AVSS.n4834 150
R4660 AVSS.n4898 AVSS.n4812 150
R4661 AVSS.n3177 AVSS.n3176 150
R4662 AVSS.n3181 AVSS.n3180 150
R4663 AVSS.n3185 AVSS.n3184 150
R4664 AVSS.n3189 AVSS.n3188 150
R4665 AVSS.n3209 AVSS.n3144 150
R4666 AVSS.n3205 AVSS.n3204 150
R4667 AVSS.n3201 AVSS.n3200 150
R4668 AVSS.n3197 AVSS.n3196 150
R4669 AVSS.n3147 AVSS.n3146 150
R4670 AVSS.n3151 AVSS.n3150 150
R4671 AVSS.n3155 AVSS.n3154 150
R4672 AVSS.n3157 AVSS.n3143 150
R4673 AVSS.n3161 AVSS.n3126 150
R4674 AVSS.n3165 AVSS.n3164 150
R4675 AVSS.n3169 AVSS.n3168 150
R4676 AVSS.n3173 AVSS.n3172 150
R4677 AVSS.n1253 AVSS.n1252 150
R4678 AVSS.n1257 AVSS.n1256 150
R4679 AVSS.n1261 AVSS.n1260 150
R4680 AVSS.n1265 AVSS.n1264 150
R4681 AVSS.n1285 AVSS.n1220 150
R4682 AVSS.n1281 AVSS.n1280 150
R4683 AVSS.n1277 AVSS.n1276 150
R4684 AVSS.n1273 AVSS.n1272 150
R4685 AVSS.n1223 AVSS.n1222 150
R4686 AVSS.n1227 AVSS.n1226 150
R4687 AVSS.n1231 AVSS.n1230 150
R4688 AVSS.n1233 AVSS.n1219 150
R4689 AVSS.n1237 AVSS.n1202 150
R4690 AVSS.n1241 AVSS.n1240 150
R4691 AVSS.n1245 AVSS.n1244 150
R4692 AVSS.n1249 AVSS.n1248 150
R4693 AVSS.n4574 AVSS.n4573 150
R4694 AVSS.n4570 AVSS.n4569 150
R4695 AVSS.n4566 AVSS.n4565 150
R4696 AVSS.n4562 AVSS.n4561 150
R4697 AVSS.n4613 AVSS.n4612 150
R4698 AVSS.n4546 AVSS.n4527 150
R4699 AVSS.n4550 AVSS.n4549 150
R4700 AVSS.n4554 AVSS.n4553 150
R4701 AVSS.n4609 AVSS.n4544 150
R4702 AVSS.n4605 AVSS.n4604 150
R4703 AVSS.n4601 AVSS.n4600 150
R4704 AVSS.n4597 AVSS.n4596 150
R4705 AVSS.n4590 AVSS.n4589 150
R4706 AVSS.n4586 AVSS.n4585 150
R4707 AVSS.n4582 AVSS.n4581 150
R4708 AVSS.n4578 AVSS.n4577 150
R4709 AVSS.n2715 AVSS.n2687 150
R4710 AVSS.n2719 AVSS.n2718 150
R4711 AVSS.n2723 AVSS.n2722 150
R4712 AVSS.n2727 AVSS.n2726 150
R4713 AVSS.n2731 AVSS.n2730 150
R4714 AVSS.n2735 AVSS.n2734 150
R4715 AVSS.n2739 AVSS.n2738 150
R4716 AVSS.n2743 AVSS.n2742 150
R4717 AVSS.n2763 AVSS.n2762 150
R4718 AVSS.n2759 AVSS.n2758 150
R4719 AVSS.n2755 AVSS.n2754 150
R4720 AVSS.n2751 AVSS.n2750 150
R4721 AVSS.n2708 AVSS.n2707 150
R4722 AVSS.n2712 AVSS.n2711 150
R4723 AVSS.n2769 AVSS.n2705 150
R4724 AVSS.n2765 AVSS.n2704 150
R4725 AVSS.n2616 AVSS.n2613 150
R4726 AVSS.n2620 AVSS.n2618 150
R4727 AVSS.n2624 AVSS.n2610 150
R4728 AVSS.n2627 AVSS.n2626 150
R4729 AVSS.n2645 AVSS.n2604 150
R4730 AVSS.n2641 AVSS.n2639 150
R4731 AVSS.n2637 AVSS.n2606 150
R4732 AVSS.n2633 AVSS.n2631 150
R4733 AVSS.n2631 AVSS.n2630 150
R4734 AVSS.n2660 AVSS.n2659 150
R4735 AVSS.n2656 AVSS.n2655 150
R4736 AVSS.n2653 AVSS.n2602 150
R4737 AVSS.n2649 AVSS.n2647 150
R4738 AVSS.n2667 AVSS.n2598 150
R4739 AVSS.n2671 AVSS.n2669 150
R4740 AVSS.n2675 AVSS.n2596 150
R4741 AVSS.n2678 AVSS.n2677 150
R4742 AVSS.n1699 AVSS.n1631 150
R4743 AVSS.n1703 AVSS.n1701 150
R4744 AVSS.n1707 AVSS.n1629 150
R4745 AVSS.n1710 AVSS.n1709 150
R4746 AVSS.n1693 AVSS.n1692 150
R4747 AVSS.n1689 AVSS.n1688 150
R4748 AVSS.n1686 AVSS.n1635 150
R4749 AVSS.n1682 AVSS.n1680 150
R4750 AVSS.n1678 AVSS.n1637 150
R4751 AVSS.n1674 AVSS.n1672 150
R4752 AVSS.n1670 AVSS.n1639 150
R4753 AVSS.n1666 AVSS.n1664 150
R4754 AVSS.n1664 AVSS.n1663 150
R4755 AVSS.n1649 AVSS.n1646 150
R4756 AVSS.n1653 AVSS.n1651 150
R4757 AVSS.n1657 AVSS.n1643 150
R4758 AVSS.n1660 AVSS.n1659 150
R4759 AVSS.n2032 AVSS.n2031 150
R4760 AVSS.n2036 AVSS.n2035 150
R4761 AVSS.n2040 AVSS.n2039 150
R4762 AVSS.n2044 AVSS.n2043 150
R4763 AVSS.n2059 AVSS.n1998 150
R4764 AVSS.n2057 AVSS.n2056 150
R4765 AVSS.n2053 AVSS.n2052 150
R4766 AVSS.n2049 AVSS.n2048 150
R4767 AVSS.n2015 AVSS.n2014 150
R4768 AVSS.n2019 AVSS.n2018 150
R4769 AVSS.n2023 AVSS.n2022 150
R4770 AVSS.n2027 AVSS.n2026 150
R4771 AVSS.n2011 AVSS.n1997 150
R4772 AVSS.n2008 AVSS.n1997 150
R4773 AVSS.n2006 AVSS.n2005 150
R4774 AVSS.n2002 AVSS.n2001 150
R4775 AVSS.n2065 AVSS.n1979 150
R4776 AVSS.n794 AVSS.n793 150
R4777 AVSS.n798 AVSS.n797 150
R4778 AVSS.n802 AVSS.n801 150
R4779 AVSS.n806 AVSS.n805 150
R4780 AVSS.n826 AVSS.n761 150
R4781 AVSS.n822 AVSS.n821 150
R4782 AVSS.n818 AVSS.n817 150
R4783 AVSS.n814 AVSS.n813 150
R4784 AVSS.n764 AVSS.n763 150
R4785 AVSS.n768 AVSS.n767 150
R4786 AVSS.n772 AVSS.n771 150
R4787 AVSS.n774 AVSS.n760 150
R4788 AVSS.n778 AVSS.n743 150
R4789 AVSS.n782 AVSS.n781 150
R4790 AVSS.n786 AVSS.n785 150
R4791 AVSS.n790 AVSS.n789 150
R4792 AVSS.n1041 AVSS.n1040 150
R4793 AVSS.n1037 AVSS.n1036 150
R4794 AVSS.n1033 AVSS.n1032 150
R4795 AVSS.n1029 AVSS.n1028 150
R4796 AVSS.n1025 AVSS.n1024 150
R4797 AVSS.n1021 AVSS.n1020 150
R4798 AVSS.n1017 AVSS.n1016 150
R4799 AVSS.n1013 AVSS.n1012 150
R4800 AVSS.n1063 AVSS.n1062 150
R4801 AVSS.n997 AVSS.n978 150
R4802 AVSS.n1001 AVSS.n1000 150
R4803 AVSS.n1005 AVSS.n1004 150
R4804 AVSS.n1059 AVSS.n995 150
R4805 AVSS.n1055 AVSS.n1054 150
R4806 AVSS.n1051 AVSS.n1050 150
R4807 AVSS.n1047 AVSS.n1046 150
R4808 AVSS.n2493 AVSS.n2423 150
R4809 AVSS.n2497 AVSS.n2495 150
R4810 AVSS.n2501 AVSS.n2421 150
R4811 AVSS.n2504 AVSS.n2503 150
R4812 AVSS.n2485 AVSS.n2425 150
R4813 AVSS.n2481 AVSS.n2479 150
R4814 AVSS.n2477 AVSS.n2427 150
R4815 AVSS.n2473 AVSS.n2471 150
R4816 AVSS.n2469 AVSS.n2429 150
R4817 AVSS.n2465 AVSS.n2464 150
R4818 AVSS.n2462 AVSS.n2432 150
R4819 AVSS.n2458 AVSS.n2457 150
R4820 AVSS.n2506 AVSS.n2419 150
R4821 AVSS.n2442 AVSS.n2440 150
R4822 AVSS.n2446 AVSS.n2437 150
R4823 AVSS.n2450 AVSS.n2448 150
R4824 AVSS.n1939 AVSS.n1906 150
R4825 AVSS.n1936 AVSS.n1906 150
R4826 AVSS.n1934 AVSS.n1933 150
R4827 AVSS.n1930 AVSS.n1929 150
R4828 AVSS.n1926 AVSS.n1893 150
R4829 AVSS.n1943 AVSS.n1942 150
R4830 AVSS.n1947 AVSS.n1946 150
R4831 AVSS.n1951 AVSS.n1950 150
R4832 AVSS.n1955 AVSS.n1954 150
R4833 AVSS.n1966 AVSS.n1907 150
R4834 AVSS.n1964 AVSS.n1963 150
R4835 AVSS.n1960 AVSS.n1959 150
R4836 AVSS.n1973 AVSS.n1888 150
R4837 AVSS.n1921 AVSS.n1920 150
R4838 AVSS.n1917 AVSS.n1916 150
R4839 AVSS.n1913 AVSS.n1912 150
R4840 AVSS.n1909 AVSS.n1889 150
R4841 AVSS.n2555 AVSS.n1771 150
R4842 AVSS.n2551 AVSS.n2550 150
R4843 AVSS.n2547 AVSS.n2546 150
R4844 AVSS.n2543 AVSS.n2542 150
R4845 AVSS.n1782 AVSS.n1781 150
R4846 AVSS.n1778 AVSS.n1777 150
R4847 AVSS.n1774 AVSS.n1773 150
R4848 AVSS.n2558 AVSS.n1752 150
R4849 AVSS.n1789 AVSS.n1753 150
R4850 AVSS.n1793 AVSS.n1792 150
R4851 AVSS.n1797 AVSS.n1796 150
R4852 AVSS.n1801 AVSS.n1800 150
R4853 AVSS.n1821 AVSS.n1820 150
R4854 AVSS.n1817 AVSS.n1816 150
R4855 AVSS.n1813 AVSS.n1812 150
R4856 AVSS.n1809 AVSS.n1808 150
R4857 AVSS.n3339 AVSS.n3338 150
R4858 AVSS.n3335 AVSS.n3334 150
R4859 AVSS.n3331 AVSS.n3330 150
R4860 AVSS.n3327 AVSS.n3307 150
R4861 AVSS.n3385 AVSS.n3325 150
R4862 AVSS.n3383 AVSS.n3382 150
R4863 AVSS.n3379 AVSS.n3378 150
R4864 AVSS.n3392 AVSS.n3306 150
R4865 AVSS.n3362 AVSS.n3361 150
R4866 AVSS.n3366 AVSS.n3365 150
R4867 AVSS.n3370 AVSS.n3369 150
R4868 AVSS.n3374 AVSS.n3373 150
R4869 AVSS.n3358 AVSS.n3324 150
R4870 AVSS.n3355 AVSS.n3324 150
R4871 AVSS.n3353 AVSS.n3352 150
R4872 AVSS.n3349 AVSS.n3348 150
R4873 AVSS.n3345 AVSS.n3311 150
R4874 AVSS.n6187 AVSS.n158 146.287
R4875 AVSS.n1321 AVSS.n1318 146.287
R4876 AVSS.n4960 AVSS.n1079 146.287
R4877 AVSS.n2185 AVSS.n2184 146.287
R4878 AVSS.n857 AVSS.n681 146.287
R4879 AVSS.n5615 AVSS.n5267 146.287
R4880 AVSS.n5444 AVSS.n5281 146.287
R4881 AVSS.n5218 AVSS.n418 146.287
R4882 AVSS.n5900 AVSS.n314 146.287
R4883 AVSS.n5676 AVSS.n5642 146.287
R4884 AVSS.n2253 AVSS.n2252 146.287
R4885 AVSS.n2390 AVSS.n2388 146.287
R4886 AVSS.n1565 AVSS.n1563 146.287
R4887 AVSS.n5015 AVSS.n634 146.287
R4888 AVSS.n3245 AVSS.n3242 146.287
R4889 AVSS.n4504 AVSS.n2789 146.287
R4890 AVSS.n4684 AVSS.n1736 146.287
R4891 AVSS.n4716 AVSS.n4715 146.287
R4892 AVSS.n4908 AVSS.n4907 146.287
R4893 AVSS.n1860 AVSS.n1859 146.287
R4894 AVSS.n4271 AVSS.n3901 146.287
R4895 AVSS.n4304 AVSS.n3690 146.287
R4896 AVSS.n4337 AVSS.n4336 146.287
R4897 AVSS.n6088 AVSS.n229 146.287
R4898 AVSS.n4420 AVSS.n4418 146.287
R4899 AVSS.t110 AVSS.n3527 141.339
R4900 AVSS.t108 AVSS.n3742 141.339
R4901 AVSS.t95 AVSS.n3953 141.339
R4902 AVSS.t102 AVSS.n216 141.339
R4903 AVSS.t85 AVSS.n167 141.339
R4904 AVSS.n6163 AVSS.n174 138.486
R4905 AVSS.n1346 AVSS.n1149 138.486
R4906 AVSS.n4939 AVSS.n1089 138.486
R4907 AVSS.n2164 AVSS.n2163 138.486
R4908 AVSS.n884 AVSS.n670 138.486
R4909 AVSS.n5848 AVSS.n5847 138.486
R4910 AVSS.n5420 AVSS.n5300 138.486
R4911 AVSS.n5224 AVSS.n5223 138.486
R4912 AVSS.n5879 AVSS.n324 138.486
R4913 AVSS.n5702 AVSS.n5631 138.486
R4914 AVSS.n2232 AVSS.n2231 138.486
R4915 AVSS.n2412 AVSS.n2411 138.486
R4916 AVSS.n1588 AVSS.n1587 138.486
R4917 AVSS.n4994 AVSS.n644 138.486
R4918 AVSS.n3271 AVSS.n3074 138.486
R4919 AVSS.n2900 AVSS.n2836 138.486
R4920 AVSS.n3040 AVSS.n3039 138.486
R4921 AVSS.n4474 AVSS.n2808 138.486
R4922 AVSS.n4932 AVSS.n1370 138.486
R4923 AVSS.n2584 AVSS.n1119 138.486
R4924 AVSS.n3968 AVSS.n3907 138.486
R4925 AVSS.n3757 AVSS.n3696 138.486
R4926 AVSS.n3620 AVSS.n3520 138.486
R4927 AVSS.n6112 AVSS.n223 138.486
R4928 AVSS.n4443 AVSS.n4442 138.486
R4929 AVSS.t9 AVSS.n293 130.019
R4930 AVSS.n5927 AVSS.n297 128.155
R4931 AVSS.n5992 AVSS.t46 128.137
R4932 AVSS.t5 AVSS.n5999 121.073
R4933 AVSS.n6013 AVSS.t117 121.073
R4934 AVSS.n6054 AVSS.t51 113.769
R4935 AVSS.t25 AVSS.n6054 113.769
R4936 AVSS.n350 AVSS.t90 107.15
R4937 AVSS.n1524 AVSS.t80 107.15
R4938 AVSS.n4773 AVSS.t78 107.15
R4939 AVSS.n4379 AVSS.t76 107.15
R4940 AVSS.t110 AVSS.n3605 107.15
R4941 AVSS.n6033 AVSS.t47 104.93
R4942 AVSS.t10 AVSS.n5964 101.525
R4943 AVSS.t47 AVSS.t0 98.6921
R4944 AVSS.n364 AVSS.t90 98.0316
R4945 AVSS.n1527 AVSS.t80 98.0316
R4946 AVSS.n4770 AVSS.t78 98.0316
R4947 AVSS.n4382 AVSS.t76 98.0316
R4948 AVSS.t110 AVSS.n3528 98.0316
R4949 AVSS.t15 AVSS.n6033 93.8322
R4950 AVSS.n5964 AVSS.n294 92.6428
R4951 AVSS.n5925 AVSS.n299 90.6806
R4952 AVSS.n5919 AVSS.n299 90.6806
R4953 AVSS.n5919 AVSS.n5918 90.6806
R4954 AVSS.n5918 AVSS.n5917 90.6806
R4955 AVSS.n5917 AVSS.n305 90.6806
R4956 AVSS.t23 AVSS.t35 83.7428
R4957 AVSS.t34 AVSS.t23 83.7428
R4958 AVSS.t38 AVSS.t34 83.7428
R4959 AVSS.t42 AVSS.t38 83.7428
R4960 AVSS.t40 AVSS.t11 83.7428
R4961 AVSS.t50 AVSS.t40 83.7428
R4962 AVSS.t126 AVSS.t50 83.7428
R4963 AVSS.t7 AVSS.t126 83.7428
R4964 AVSS.t14 AVSS.t44 83.7428
R4965 AVSS.t12 AVSS.t14 83.7428
R4966 AVSS.t36 AVSS.t12 83.7428
R4967 AVSS.t33 AVSS.t32 83.7428
R4968 AVSS.t32 AVSS.t39 83.7428
R4969 AVSS.t39 AVSS.t46 83.7428
R4970 AVSS.t130 AVSS.t30 83.7428
R4971 AVSS.t22 AVSS.t127 83.7428
R4972 AVSS.n6000 AVSS.t118 83.7172
R4973 AVSS.n6001 AVSS.t121 83.7172
R4974 AVSS.n6001 AVSS.t119 83.7172
R4975 AVSS.n6002 AVSS.t115 83.7172
R4976 AVSS.n6002 AVSS.t120 83.7172
R4977 AVSS.n6003 AVSS.t116 83.7172
R4978 AVSS.n3883 AVSS.n3872 83.5719
R4979 AVSS.n3873 AVSS.n188 83.5719
R4980 AVSS.n3878 AVSS.n187 83.5719
R4981 AVSS.n4094 AVSS.n4083 83.5719
R4982 AVSS.n4084 AVSS.n190 83.5719
R4983 AVSS.n4089 AVSS.n189 83.5719
R4984 AVSS.n4104 AVSS.n4103 83.5719
R4985 AVSS.n4099 AVSS.n192 83.5719
R4986 AVSS.n4109 AVSS.n191 83.5719
R4987 AVSS.n3650 AVSS.n3649 83.5719
R4988 AVSS.n3644 AVSS.n194 83.5719
R4989 AVSS.n3654 AVSS.n193 83.5719
R4990 AVSS.n3412 AVSS.n3411 83.5719
R4991 AVSS.n3401 AVSS.n2798 83.5719
R4992 AVSS.n3400 AVSS.n2797 83.5719
R4993 AVSS.n1615 AVSS.n1614 83.5719
R4994 AVSS.n1613 AVSS.n1612 83.5719
R4995 AVSS.n1602 AVSS.n1601 83.5719
R4996 AVSS.n5020 AVSS.n5019 83.5719
R4997 AVSS.n5018 AVSS.n5017 83.5719
R4998 AVSS.n570 AVSS.n569 83.5719
R4999 AVSS.n5038 AVSS.n454 83.5719
R5000 AVSS.n456 AVSS.n455 83.5719
R5001 AVSS.n5032 AVSS.n5031 83.5719
R5002 AVSS.n581 AVSS.n572 83.5719
R5003 AVSS.n591 AVSS.n590 83.5719
R5004 AVSS.n577 AVSS.n571 83.5719
R5005 AVSS.n1102 AVSS.n1093 83.5719
R5006 AVSS.n1112 AVSS.n1111 83.5719
R5007 AVSS.n1098 AVSS.n1092 83.5719
R5008 AVSS.n4487 AVSS.n4478 83.5719
R5009 AVSS.n4497 AVSS.n4496 83.5719
R5010 AVSS.n4483 AVSS.n4477 83.5719
R5011 AVSS.n6227 AVSS.n38 83.5719
R5012 AVSS.n6236 AVSS.n6235 83.5719
R5013 AVSS.n6238 AVSS.n6237 83.5719
R5014 AVSS.n6247 AVSS.n6246 83.5719
R5015 AVSS.n30 AVSS.n27 83.5719
R5016 AVSS.n6252 AVSS.n26 83.5719
R5017 AVSS.n6258 AVSS.n21 83.5719
R5018 AVSS.n6265 AVSS.n6264 83.5719
R5019 AVSS.n5051 AVSS.n20 83.5719
R5020 AVSS.n5057 AVSS.n450 83.5719
R5021 AVSS.n5064 AVSS.n5063 83.5719
R5022 AVSS.n5046 AVSS.n449 83.5719
R5023 AVSS.n268 AVSS.n267 83.5719
R5024 AVSS.n272 AVSS.n196 83.5719
R5025 AVSS.n271 AVSS.n195 83.5719
R5026 AVSS.t48 AVSS.t27 78.698
R5027 AVSS.t99 AVSS.n448 77.948
R5028 AVSS.t89 AVSS.n19 77.948
R5029 AVSS.n5582 AVSS.t92 77.948
R5030 AVSS.t106 AVSS.n37 77.948
R5031 AVSS.n5999 AVSS.n5998 76.6802
R5032 AVSS.n258 AVSS.n257 76.3222
R5033 AVSS.n255 AVSS.n254 76.3222
R5034 AVSS.n248 AVSS.n234 76.3222
R5035 AVSS.n247 AVSS.n246 76.3222
R5036 AVSS.n240 AVSS.n236 76.3222
R5037 AVSS.n239 AVSS.n238 76.3222
R5038 AVSS.n6208 AVSS.n150 76.3222
R5039 AVSS.n6206 AVSS.n6205 76.3222
R5040 AVSS.n6201 AVSS.n154 76.3222
R5041 AVSS.n6199 AVSS.n6198 76.3222
R5042 AVSS.n6194 AVSS.n157 76.3222
R5043 AVSS.n6192 AVSS.n6191 76.3222
R5044 AVSS.n1193 AVSS.n1165 76.3222
R5045 AVSS.n1191 AVSS.n1167 76.3222
R5046 AVSS.n1172 AVSS.n1171 76.3222
R5047 AVSS.n1185 AVSS.n1170 76.3222
R5048 AVSS.n1181 AVSS.n1169 76.3222
R5049 AVSS.n1177 AVSS.n1168 76.3222
R5050 AVSS.n1297 AVSS.n1296 76.3222
R5051 AVSS.n1298 AVSS.n1163 76.3222
R5052 AVSS.n1305 AVSS.n1304 76.3222
R5053 AVSS.n1306 AVSS.n1161 76.3222
R5054 AVSS.n1313 AVSS.n1312 76.3222
R5055 AVSS.n1317 AVSS.n1159 76.3222
R5056 AVSS.n1368 AVSS.n1367 76.3222
R5057 AVSS.n1363 AVSS.n1144 76.3222
R5058 AVSS.n1359 AVSS.n1143 76.3222
R5059 AVSS.n1355 AVSS.n1142 76.3222
R5060 AVSS.n1351 AVSS.n1141 76.3222
R5061 AVSS.n1347 AVSS.n1140 76.3222
R5062 AVSS.n4626 AVSS.n4625 76.3222
R5063 AVSS.n4629 AVSS.n4628 76.3222
R5064 AVSS.n4634 AVSS.n4633 76.3222
R5065 AVSS.n4637 AVSS.n4636 76.3222
R5066 AVSS.n4642 AVSS.n4641 76.3222
R5067 AVSS.n4645 AVSS.n4644 76.3222
R5068 AVSS.n4978 AVSS.n4977 76.3222
R5069 AVSS.n4975 AVSS.n4974 76.3222
R5070 AVSS.n4970 AVSS.n1075 76.3222
R5071 AVSS.n4968 AVSS.n4967 76.3222
R5072 AVSS.n4963 AVSS.n1078 76.3222
R5073 AVSS.n4961 AVSS.n4960 76.3222
R5074 AVSS.n4956 AVSS.n1081 76.3222
R5075 AVSS.n4954 AVSS.n4953 76.3222
R5076 AVSS.n4949 AVSS.n1085 76.3222
R5077 AVSS.n4947 AVSS.n4946 76.3222
R5078 AVSS.n4942 AVSS.n1088 76.3222
R5079 AVSS.n4940 AVSS.n4939 76.3222
R5080 AVSS.n4663 AVSS.n1127 76.3222
R5081 AVSS.n4659 AVSS.n1128 76.3222
R5082 AVSS.n4655 AVSS.n1129 76.3222
R5083 AVSS.n4651 AVSS.n1130 76.3222
R5084 AVSS.n1131 AVSS.n1091 76.3222
R5085 AVSS.n4934 AVSS.n1089 76.3222
R5086 AVSS.n2116 AVSS.n2115 76.3222
R5087 AVSS.n2119 AVSS.n2118 76.3222
R5088 AVSS.n2124 AVSS.n2123 76.3222
R5089 AVSS.n2127 AVSS.n2126 76.3222
R5090 AVSS.n2132 AVSS.n2131 76.3222
R5091 AVSS.n2135 AVSS.n2134 76.3222
R5092 AVSS.n2110 AVSS.n2109 76.3222
R5093 AVSS.n2107 AVSS.n2106 76.3222
R5094 AVSS.n2102 AVSS.n2094 76.3222
R5095 AVSS.n2100 AVSS.n2099 76.3222
R5096 AVSS.n2095 AVSS.n2071 76.3222
R5097 AVSS.n2186 AVSS.n2185 76.3222
R5098 AVSS.n2183 AVSS.n2182 76.3222
R5099 AVSS.n2178 AVSS.n2076 76.3222
R5100 AVSS.n2176 AVSS.n2175 76.3222
R5101 AVSS.n2171 AVSS.n2079 76.3222
R5102 AVSS.n2169 AVSS.n2168 76.3222
R5103 AVSS.n2164 AVSS.n2162 76.3222
R5104 AVSS.n2142 AVSS.n1138 76.3222
R5105 AVSS.n2146 AVSS.n1137 76.3222
R5106 AVSS.n2150 AVSS.n1136 76.3222
R5107 AVSS.n2154 AVSS.n1135 76.3222
R5108 AVSS.n2158 AVSS.n1134 76.3222
R5109 AVSS.n2163 AVSS.n1133 76.3222
R5110 AVSS.n836 AVSS.n632 76.3222
R5111 AVSS.n840 AVSS.n631 76.3222
R5112 AVSS.n844 AVSS.n630 76.3222
R5113 AVSS.n848 AVSS.n629 76.3222
R5114 AVSS.n852 AVSS.n628 76.3222
R5115 AVSS.n682 AVSS.n627 76.3222
R5116 AVSS.n735 AVSS.n648 76.3222
R5117 AVSS.n731 AVSS.n649 76.3222
R5118 AVSS.n727 AVSS.n650 76.3222
R5119 AVSS.n723 AVSS.n651 76.3222
R5120 AVSS.n719 AVSS.n652 76.3222
R5121 AVSS.n669 AVSS.n653 76.3222
R5122 AVSS.n692 AVSS.n691 76.3222
R5123 AVSS.n697 AVSS.n696 76.3222
R5124 AVSS.n700 AVSS.n699 76.3222
R5125 AVSS.n705 AVSS.n704 76.3222
R5126 AVSS.n708 AVSS.n707 76.3222
R5127 AVSS.n713 AVSS.n712 76.3222
R5128 AVSS.n5611 AVSS.n5260 76.3222
R5129 AVSS.n5607 AVSS.n5261 76.3222
R5130 AVSS.n5603 AVSS.n5262 76.3222
R5131 AVSS.n5599 AVSS.n5263 76.3222
R5132 AVSS.n5595 AVSS.n5264 76.3222
R5133 AVSS.n5847 AVSS.n5846 76.3222
R5134 AVSS.n5868 AVSS.n5254 76.3222
R5135 AVSS.n5864 AVSS.n5253 76.3222
R5136 AVSS.n5860 AVSS.n5252 76.3222
R5137 AVSS.n5856 AVSS.n5251 76.3222
R5138 AVSS.n5852 AVSS.n5250 76.3222
R5139 AVSS.n5848 AVSS.n5249 76.3222
R5140 AVSS.n5566 AVSS.n5447 76.3222
R5141 AVSS.n5564 AVSS.n5449 76.3222
R5142 AVSS.n5454 AVSS.n5453 76.3222
R5143 AVSS.n5558 AVSS.n5452 76.3222
R5144 AVSS.n5554 AVSS.n5451 76.3222
R5145 AVSS.n5550 AVSS.n5450 76.3222
R5146 AVSS.n5567 AVSS.n5566 76.3222
R5147 AVSS.n5564 AVSS.n5563 76.3222
R5148 AVSS.n5559 AVSS.n5453 76.3222
R5149 AVSS.n5555 AVSS.n5452 76.3222
R5150 AVSS.n5551 AVSS.n5451 76.3222
R5151 AVSS.n5450 AVSS.n5255 76.3222
R5152 AVSS.n6280 AVSS.n6279 76.3222
R5153 AVSS.n6283 AVSS.n6282 76.3222
R5154 AVSS.n6288 AVSS.n6287 76.3222
R5155 AVSS.n6291 AVSS.n6290 76.3222
R5156 AVSS.n6296 AVSS.n6295 76.3222
R5157 AVSS.n6299 AVSS.n6298 76.3222
R5158 AVSS.n5399 AVSS.n334 76.3222
R5159 AVSS.n5403 AVSS.n335 76.3222
R5160 AVSS.n5407 AVSS.n336 76.3222
R5161 AVSS.n5411 AVSS.n337 76.3222
R5162 AVSS.n5415 AVSS.n338 76.3222
R5163 AVSS.n5300 AVSS.n339 76.3222
R5164 AVSS.n5439 AVSS.n5281 76.3222
R5165 AVSS.n5438 AVSS.n5437 76.3222
R5166 AVSS.n5431 AVSS.n5296 76.3222
R5167 AVSS.n5430 AVSS.n5429 76.3222
R5168 AVSS.n5423 AVSS.n5298 76.3222
R5169 AVSS.n5422 AVSS.n5421 76.3222
R5170 AVSS.n5421 AVSS.n5420 76.3222
R5171 AVSS.n5424 AVSS.n5423 76.3222
R5172 AVSS.n5429 AVSS.n5428 76.3222
R5173 AVSS.n5432 AVSS.n5431 76.3222
R5174 AVSS.n5437 AVSS.n5436 76.3222
R5175 AVSS.n5440 AVSS.n5439 76.3222
R5176 AVSS.n6281 AVSS.n6280 76.3222
R5177 AVSS.n6282 AVSS.n9 76.3222
R5178 AVSS.n6289 AVSS.n6288 76.3222
R5179 AVSS.n6290 AVSS.n7 76.3222
R5180 AVSS.n6297 AVSS.n6296 76.3222
R5181 AVSS.n6300 AVSS.n6299 76.3222
R5182 AVSS.n5094 AVSS.n5093 76.3222
R5183 AVSS.n5089 AVSS.n426 76.3222
R5184 AVSS.n5086 AVSS.n425 76.3222
R5185 AVSS.n5082 AVSS.n424 76.3222
R5186 AVSS.n5078 AVSS.n423 76.3222
R5187 AVSS.n5097 AVSS.n5096 76.3222
R5188 AVSS.n5244 AVSS.n405 76.3222
R5189 AVSS.n5240 AVSS.n404 76.3222
R5190 AVSS.n5236 AVSS.n403 76.3222
R5191 AVSS.n5232 AVSS.n402 76.3222
R5192 AVSS.n5228 AVSS.n401 76.3222
R5193 AVSS.n5224 AVSS.n400 76.3222
R5194 AVSS.n418 AVSS.n411 76.3222
R5195 AVSS.n5213 AVSS.n412 76.3222
R5196 AVSS.n5209 AVSS.n413 76.3222
R5197 AVSS.n5205 AVSS.n414 76.3222
R5198 AVSS.n5201 AVSS.n415 76.3222
R5199 AVSS.n5222 AVSS.n410 76.3222
R5200 AVSS.n5223 AVSS.n5222 76.3222
R5201 AVSS.n5198 AVSS.n415 76.3222
R5202 AVSS.n5202 AVSS.n414 76.3222
R5203 AVSS.n5206 AVSS.n413 76.3222
R5204 AVSS.n5210 AVSS.n412 76.3222
R5205 AVSS.n5214 AVSS.n411 76.3222
R5206 AVSS.n391 AVSS.n341 76.3222
R5207 AVSS.n387 AVSS.n342 76.3222
R5208 AVSS.n383 AVSS.n343 76.3222
R5209 AVSS.n379 AVSS.n344 76.3222
R5210 AVSS.n345 AVSS.n327 76.3222
R5211 AVSS.n5874 AVSS.n324 76.3222
R5212 AVSS.n5896 AVSS.n316 76.3222
R5213 AVSS.n5894 AVSS.n5893 76.3222
R5214 AVSS.n5889 AVSS.n320 76.3222
R5215 AVSS.n5887 AVSS.n5886 76.3222
R5216 AVSS.n5882 AVSS.n323 76.3222
R5217 AVSS.n5880 AVSS.n5879 76.3222
R5218 AVSS.n5881 AVSS.n5880 76.3222
R5219 AVSS.n323 AVSS.n321 76.3222
R5220 AVSS.n5888 AVSS.n5887 76.3222
R5221 AVSS.n320 AVSS.n318 76.3222
R5222 AVSS.n5895 AVSS.n5894 76.3222
R5223 AVSS.n316 AVSS.n314 76.3222
R5224 AVSS.n5094 AVSS.n427 76.3222
R5225 AVSS.n5087 AVSS.n426 76.3222
R5226 AVSS.n5083 AVSS.n425 76.3222
R5227 AVSS.n5079 AVSS.n424 76.3222
R5228 AVSS.n423 AVSS.n422 76.3222
R5229 AVSS.n5096 AVSS.n406 76.3222
R5230 AVSS.n5846 AVSS.n5259 76.3222
R5231 AVSS.n5598 AVSS.n5264 76.3222
R5232 AVSS.n5602 AVSS.n5263 76.3222
R5233 AVSS.n5606 AVSS.n5262 76.3222
R5234 AVSS.n5610 AVSS.n5261 76.3222
R5235 AVSS.n5267 AVSS.n5260 76.3222
R5236 AVSS.n5723 AVSS.n328 76.3222
R5237 AVSS.n5719 AVSS.n329 76.3222
R5238 AVSS.n5715 AVSS.n330 76.3222
R5239 AVSS.n5711 AVSS.n331 76.3222
R5240 AVSS.n5707 AVSS.n332 76.3222
R5241 AVSS.n5703 AVSS.n333 76.3222
R5242 AVSS.n5842 AVSS.n5623 76.3222
R5243 AVSS.n5835 AVSS.n5622 76.3222
R5244 AVSS.n5831 AVSS.n5621 76.3222
R5245 AVSS.n5827 AVSS.n5620 76.3222
R5246 AVSS.n5823 AVSS.n5619 76.3222
R5247 AVSS.n5627 AVSS.n5618 76.3222
R5248 AVSS.n5842 AVSS.n5841 76.3222
R5249 AVSS.n5837 AVSS.n5622 76.3222
R5250 AVSS.n5834 AVSS.n5621 76.3222
R5251 AVSS.n5830 AVSS.n5620 76.3222
R5252 AVSS.n5826 AVSS.n5619 76.3222
R5253 AVSS.n5822 AVSS.n5618 76.3222
R5254 AVSS.n2273 AVSS.n607 76.3222
R5255 AVSS.n2269 AVSS.n608 76.3222
R5256 AVSS.n2265 AVSS.n609 76.3222
R5257 AVSS.n2261 AVSS.n610 76.3222
R5258 AVSS.n2257 AVSS.n611 76.3222
R5259 AVSS.n2253 AVSS.n612 76.3222
R5260 AVSS.n2251 AVSS.n2250 76.3222
R5261 AVSS.n2246 AVSS.n2204 76.3222
R5262 AVSS.n2244 AVSS.n2243 76.3222
R5263 AVSS.n2239 AVSS.n2207 76.3222
R5264 AVSS.n2237 AVSS.n2236 76.3222
R5265 AVSS.n2232 AVSS.n2230 76.3222
R5266 AVSS.n2210 AVSS.n970 76.3222
R5267 AVSS.n2214 AVSS.n969 76.3222
R5268 AVSS.n2218 AVSS.n968 76.3222
R5269 AVSS.n2222 AVSS.n967 76.3222
R5270 AVSS.n2226 AVSS.n966 76.3222
R5271 AVSS.n2231 AVSS.n965 76.3222
R5272 AVSS.n2280 AVSS.n2279 76.3222
R5273 AVSS.n2283 AVSS.n2282 76.3222
R5274 AVSS.n2288 AVSS.n2287 76.3222
R5275 AVSS.n2291 AVSS.n2290 76.3222
R5276 AVSS.n2296 AVSS.n2295 76.3222
R5277 AVSS.n2299 AVSS.n2298 76.3222
R5278 AVSS.n2368 AVSS.n625 76.3222
R5279 AVSS.n2372 AVSS.n624 76.3222
R5280 AVSS.n2376 AVSS.n623 76.3222
R5281 AVSS.n2380 AVSS.n622 76.3222
R5282 AVSS.n2384 AVSS.n621 76.3222
R5283 AVSS.n2388 AVSS.n620 76.3222
R5284 AVSS.n2389 AVSS.n2309 76.3222
R5285 AVSS.n2396 AVSS.n2395 76.3222
R5286 AVSS.n2397 AVSS.n2307 76.3222
R5287 AVSS.n2404 AVSS.n2403 76.3222
R5288 AVSS.n2408 AVSS.n2305 76.3222
R5289 AVSS.n2412 AVSS.n2410 76.3222
R5290 AVSS.n2334 AVSS.n655 76.3222
R5291 AVSS.n2330 AVSS.n656 76.3222
R5292 AVSS.n2326 AVSS.n657 76.3222
R5293 AVSS.n2322 AVSS.n658 76.3222
R5294 AVSS.n2318 AVSS.n659 76.3222
R5295 AVSS.n2411 AVSS.n660 76.3222
R5296 AVSS.n2362 AVSS.n2361 76.3222
R5297 AVSS.n2359 AVSS.n2311 76.3222
R5298 AVSS.n2355 AVSS.n2354 76.3222
R5299 AVSS.n2348 AVSS.n2313 76.3222
R5300 AVSS.n2347 AVSS.n2346 76.3222
R5301 AVSS.n2339 AVSS.n2315 76.3222
R5302 AVSS.n1543 AVSS.n614 76.3222
R5303 AVSS.n1547 AVSS.n615 76.3222
R5304 AVSS.n1551 AVSS.n616 76.3222
R5305 AVSS.n1555 AVSS.n617 76.3222
R5306 AVSS.n1559 AVSS.n618 76.3222
R5307 AVSS.n1563 AVSS.n619 76.3222
R5308 AVSS.n1508 AVSS.n662 76.3222
R5309 AVSS.n1504 AVSS.n663 76.3222
R5310 AVSS.n1500 AVSS.n664 76.3222
R5311 AVSS.n1496 AVSS.n665 76.3222
R5312 AVSS.n1590 AVSS.n666 76.3222
R5313 AVSS.n1588 AVSS.n667 76.3222
R5314 AVSS.n1564 AVSS.n1389 76.3222
R5315 AVSS.n1571 AVSS.n1570 76.3222
R5316 AVSS.n1572 AVSS.n1387 76.3222
R5317 AVSS.n1579 AVSS.n1578 76.3222
R5318 AVSS.n1580 AVSS.n1385 76.3222
R5319 AVSS.n1587 AVSS.n1586 76.3222
R5320 AVSS.n1586 AVSS.n1585 76.3222
R5321 AVSS.n1581 AVSS.n1580 76.3222
R5322 AVSS.n1578 AVSS.n1577 76.3222
R5323 AVSS.n1573 AVSS.n1572 76.3222
R5324 AVSS.n1570 AVSS.n1569 76.3222
R5325 AVSS.n1565 AVSS.n1564 76.3222
R5326 AVSS.n2361 AVSS.n2360 76.3222
R5327 AVSS.n2356 AVSS.n2311 76.3222
R5328 AVSS.n2354 AVSS.n2353 76.3222
R5329 AVSS.n2349 AVSS.n2348 76.3222
R5330 AVSS.n2346 AVSS.n2345 76.3222
R5331 AVSS.n2340 AVSS.n2339 76.3222
R5332 AVSS.n2410 AVSS.n2409 76.3222
R5333 AVSS.n2405 AVSS.n2305 76.3222
R5334 AVSS.n2403 AVSS.n2402 76.3222
R5335 AVSS.n2398 AVSS.n2397 76.3222
R5336 AVSS.n2395 AVSS.n2394 76.3222
R5337 AVSS.n2390 AVSS.n2389 76.3222
R5338 AVSS.n2281 AVSS.n2280 76.3222
R5339 AVSS.n2282 AVSS.n2199 76.3222
R5340 AVSS.n2289 AVSS.n2288 76.3222
R5341 AVSS.n2290 AVSS.n2197 76.3222
R5342 AVSS.n2297 AVSS.n2296 76.3222
R5343 AVSS.n2298 AVSS.n971 76.3222
R5344 AVSS.n2230 AVSS.n2208 76.3222
R5345 AVSS.n2238 AVSS.n2237 76.3222
R5346 AVSS.n2207 AVSS.n2205 76.3222
R5347 AVSS.n2245 AVSS.n2244 76.3222
R5348 AVSS.n2204 AVSS.n2202 76.3222
R5349 AVSS.n2252 AVSS.n2251 76.3222
R5350 AVSS.n691 AVSS.n689 76.3222
R5351 AVSS.n698 AVSS.n697 76.3222
R5352 AVSS.n699 AVSS.n687 76.3222
R5353 AVSS.n706 AVSS.n705 76.3222
R5354 AVSS.n707 AVSS.n685 76.3222
R5355 AVSS.n714 AVSS.n713 76.3222
R5356 AVSS.n1560 AVSS.n619 76.3222
R5357 AVSS.n1556 AVSS.n618 76.3222
R5358 AVSS.n1552 AVSS.n617 76.3222
R5359 AVSS.n1548 AVSS.n616 76.3222
R5360 AVSS.n1544 AVSS.n615 76.3222
R5361 AVSS.n1540 AVSS.n614 76.3222
R5362 AVSS.n2385 AVSS.n620 76.3222
R5363 AVSS.n2381 AVSS.n621 76.3222
R5364 AVSS.n2377 AVSS.n622 76.3222
R5365 AVSS.n2373 AVSS.n623 76.3222
R5366 AVSS.n2369 AVSS.n624 76.3222
R5367 AVSS.n2365 AVSS.n625 76.3222
R5368 AVSS.n2256 AVSS.n612 76.3222
R5369 AVSS.n2260 AVSS.n611 76.3222
R5370 AVSS.n2264 AVSS.n610 76.3222
R5371 AVSS.n2268 AVSS.n609 76.3222
R5372 AVSS.n2272 AVSS.n608 76.3222
R5373 AVSS.n2275 AVSS.n607 76.3222
R5374 AVSS.n853 AVSS.n627 76.3222
R5375 AVSS.n849 AVSS.n628 76.3222
R5376 AVSS.n845 AVSS.n629 76.3222
R5377 AVSS.n841 AVSS.n630 76.3222
R5378 AVSS.n837 AVSS.n631 76.3222
R5379 AVSS.n690 AVSS.n632 76.3222
R5380 AVSS.n5875 AVSS.n5874 76.3222
R5381 AVSS.n378 AVSS.n345 76.3222
R5382 AVSS.n382 AVSS.n344 76.3222
R5383 AVSS.n386 AVSS.n343 76.3222
R5384 AVSS.n390 AVSS.n342 76.3222
R5385 AVSS.n393 AVSS.n341 76.3222
R5386 AVSS.n5227 AVSS.n400 76.3222
R5387 AVSS.n5231 AVSS.n401 76.3222
R5388 AVSS.n5235 AVSS.n402 76.3222
R5389 AVSS.n5239 AVSS.n403 76.3222
R5390 AVSS.n5243 AVSS.n404 76.3222
R5391 AVSS.n407 AVSS.n405 76.3222
R5392 AVSS.n5416 AVSS.n339 76.3222
R5393 AVSS.n5412 AVSS.n338 76.3222
R5394 AVSS.n5408 AVSS.n337 76.3222
R5395 AVSS.n5404 AVSS.n336 76.3222
R5396 AVSS.n5400 AVSS.n335 76.3222
R5397 AVSS.n5396 AVSS.n334 76.3222
R5398 AVSS.n5851 AVSS.n5249 76.3222
R5399 AVSS.n5855 AVSS.n5250 76.3222
R5400 AVSS.n5859 AVSS.n5251 76.3222
R5401 AVSS.n5863 AVSS.n5252 76.3222
R5402 AVSS.n5867 AVSS.n5253 76.3222
R5403 AVSS.n5256 AVSS.n5254 76.3222
R5404 AVSS.n5706 AVSS.n333 76.3222
R5405 AVSS.n5710 AVSS.n332 76.3222
R5406 AVSS.n5714 AVSS.n331 76.3222
R5407 AVSS.n5718 AVSS.n330 76.3222
R5408 AVSS.n5722 AVSS.n329 76.3222
R5409 AVSS.n5628 AVSS.n328 76.3222
R5410 AVSS.n5011 AVSS.n637 76.3222
R5411 AVSS.n5009 AVSS.n5008 76.3222
R5412 AVSS.n5004 AVSS.n640 76.3222
R5413 AVSS.n5002 AVSS.n5001 76.3222
R5414 AVSS.n4997 AVSS.n643 76.3222
R5415 AVSS.n4995 AVSS.n4994 76.3222
R5416 AVSS.n960 AVSS.n891 76.3222
R5417 AVSS.n956 AVSS.n890 76.3222
R5418 AVSS.n952 AVSS.n889 76.3222
R5419 AVSS.n948 AVSS.n888 76.3222
R5420 AVSS.n887 AVSS.n647 76.3222
R5421 AVSS.n4989 AVSS.n644 76.3222
R5422 AVSS.n923 AVSS.n922 76.3222
R5423 AVSS.n926 AVSS.n925 76.3222
R5424 AVSS.n931 AVSS.n930 76.3222
R5425 AVSS.n934 AVSS.n933 76.3222
R5426 AVSS.n939 AVSS.n938 76.3222
R5427 AVSS.n942 AVSS.n941 76.3222
R5428 AVSS.n899 AVSS.n600 76.3222
R5429 AVSS.n917 AVSS.n601 76.3222
R5430 AVSS.n913 AVSS.n602 76.3222
R5431 AVSS.n909 AVSS.n603 76.3222
R5432 AVSS.n905 AVSS.n604 76.3222
R5433 AVSS.n901 AVSS.n605 76.3222
R5434 AVSS.n633 AVSS.n605 76.3222
R5435 AVSS.n902 AVSS.n604 76.3222
R5436 AVSS.n906 AVSS.n603 76.3222
R5437 AVSS.n910 AVSS.n602 76.3222
R5438 AVSS.n914 AVSS.n601 76.3222
R5439 AVSS.n918 AVSS.n600 76.3222
R5440 AVSS.n924 AVSS.n923 76.3222
R5441 AVSS.n925 AVSS.n897 76.3222
R5442 AVSS.n932 AVSS.n931 76.3222
R5443 AVSS.n933 AVSS.n895 76.3222
R5444 AVSS.n940 AVSS.n939 76.3222
R5445 AVSS.n941 AVSS.n892 76.3222
R5446 AVSS.n4996 AVSS.n4995 76.3222
R5447 AVSS.n643 AVSS.n641 76.3222
R5448 AVSS.n5003 AVSS.n5002 76.3222
R5449 AVSS.n640 AVSS.n638 76.3222
R5450 AVSS.n5010 AVSS.n5009 76.3222
R5451 AVSS.n637 AVSS.n634 76.3222
R5452 AVSS.n3221 AVSS.n3220 76.3222
R5453 AVSS.n3222 AVSS.n3089 76.3222
R5454 AVSS.n3229 AVSS.n3228 76.3222
R5455 AVSS.n3230 AVSS.n3087 76.3222
R5456 AVSS.n3237 AVSS.n3236 76.3222
R5457 AVSS.n3241 AVSS.n3085 76.3222
R5458 AVSS.n3293 AVSS.n3292 76.3222
R5459 AVSS.n3288 AVSS.n3069 76.3222
R5460 AVSS.n3284 AVSS.n3068 76.3222
R5461 AVSS.n3280 AVSS.n3067 76.3222
R5462 AVSS.n3276 AVSS.n3066 76.3222
R5463 AVSS.n3272 AVSS.n3065 76.3222
R5464 AVSS.n3118 AVSS.n3091 76.3222
R5465 AVSS.n3117 AVSS.n3116 76.3222
R5466 AVSS.n3110 AVSS.n3093 76.3222
R5467 AVSS.n3109 AVSS.n3108 76.3222
R5468 AVSS.n3102 AVSS.n3095 76.3222
R5469 AVSS.n3101 AVSS.n3100 76.3222
R5470 AVSS.n3119 AVSS.n3118 76.3222
R5471 AVSS.n3116 AVSS.n3115 76.3222
R5472 AVSS.n3111 AVSS.n3110 76.3222
R5473 AVSS.n3108 AVSS.n3107 76.3222
R5474 AVSS.n3103 AVSS.n3102 76.3222
R5475 AVSS.n3100 AVSS.n3099 76.3222
R5476 AVSS.n4521 AVSS.n2782 76.3222
R5477 AVSS.n4519 AVSS.n4518 76.3222
R5478 AVSS.n4514 AVSS.n2785 76.3222
R5479 AVSS.n4512 AVSS.n4511 76.3222
R5480 AVSS.n4507 AVSS.n2788 76.3222
R5481 AVSS.n4505 AVSS.n4504 76.3222
R5482 AVSS.n4675 AVSS.n4674 76.3222
R5483 AVSS.n2841 AVSS.n2778 76.3222
R5484 AVSS.n2846 AVSS.n2845 76.3222
R5485 AVSS.n2849 AVSS.n2848 76.3222
R5486 AVSS.n2854 AVSS.n2853 76.3222
R5487 AVSS.n2857 AVSS.n2856 76.3222
R5488 AVSS.n2864 AVSS.n2830 76.3222
R5489 AVSS.n2868 AVSS.n2831 76.3222
R5490 AVSS.n2872 AVSS.n2832 76.3222
R5491 AVSS.n2876 AVSS.n2833 76.3222
R5492 AVSS.n2879 AVSS.n2834 76.3222
R5493 AVSS.n2901 AVSS.n2900 76.3222
R5494 AVSS.n4499 AVSS.n2789 76.3222
R5495 AVSS.n2792 AVSS.n2791 76.3222
R5496 AVSS.n2884 AVSS.n2793 76.3222
R5497 AVSS.n2888 AVSS.n2794 76.3222
R5498 AVSS.n2892 AVSS.n2795 76.3222
R5499 AVSS.n2896 AVSS.n2796 76.3222
R5500 AVSS.n2836 AVSS.n2796 76.3222
R5501 AVSS.n2895 AVSS.n2795 76.3222
R5502 AVSS.n2891 AVSS.n2794 76.3222
R5503 AVSS.n2887 AVSS.n2793 76.3222
R5504 AVSS.n2883 AVSS.n2792 76.3222
R5505 AVSS.n4500 AVSS.n4499 76.3222
R5506 AVSS.n4676 AVSS.n4675 76.3222
R5507 AVSS.n2842 AVSS.n2841 76.3222
R5508 AVSS.n2847 AVSS.n2846 76.3222
R5509 AVSS.n2848 AVSS.n2839 76.3222
R5510 AVSS.n2855 AVSS.n2854 76.3222
R5511 AVSS.n2858 AVSS.n2857 76.3222
R5512 AVSS.n4701 AVSS.n1729 76.3222
R5513 AVSS.n4699 AVSS.n4698 76.3222
R5514 AVSS.n4694 AVSS.n1732 76.3222
R5515 AVSS.n4692 AVSS.n4691 76.3222
R5516 AVSS.n4687 AVSS.n1735 76.3222
R5517 AVSS.n4685 AVSS.n4684 76.3222
R5518 AVSS.n4707 AVSS.n4706 76.3222
R5519 AVSS.n2994 AVSS.n1725 76.3222
R5520 AVSS.n2999 AVSS.n2998 76.3222
R5521 AVSS.n3002 AVSS.n3001 76.3222
R5522 AVSS.n3007 AVSS.n3006 76.3222
R5523 AVSS.n3010 AVSS.n3009 76.3222
R5524 AVSS.n3060 AVSS.n2988 76.3222
R5525 AVSS.n3056 AVSS.n2987 76.3222
R5526 AVSS.n3052 AVSS.n2986 76.3222
R5527 AVSS.n3048 AVSS.n2985 76.3222
R5528 AVSS.n3044 AVSS.n2984 76.3222
R5529 AVSS.n3040 AVSS.n2983 76.3222
R5530 AVSS.n3018 AVSS.n1736 76.3222
R5531 AVSS.n3022 AVSS.n3021 76.3222
R5532 AVSS.n3025 AVSS.n3024 76.3222
R5533 AVSS.n3030 AVSS.n3029 76.3222
R5534 AVSS.n3033 AVSS.n3032 76.3222
R5535 AVSS.n3038 AVSS.n3037 76.3222
R5536 AVSS.n3039 AVSS.n3038 76.3222
R5537 AVSS.n3032 AVSS.n3014 76.3222
R5538 AVSS.n3031 AVSS.n3030 76.3222
R5539 AVSS.n3024 AVSS.n3016 76.3222
R5540 AVSS.n3023 AVSS.n3022 76.3222
R5541 AVSS.n3019 AVSS.n3018 76.3222
R5542 AVSS.n4708 AVSS.n4707 76.3222
R5543 AVSS.n2995 AVSS.n2994 76.3222
R5544 AVSS.n3000 AVSS.n2999 76.3222
R5545 AVSS.n3001 AVSS.n2992 76.3222
R5546 AVSS.n3008 AVSS.n3007 76.3222
R5547 AVSS.n3009 AVSS.n2989 76.3222
R5548 AVSS.n2936 AVSS.n2935 76.3222
R5549 AVSS.n2931 AVSS.n2918 76.3222
R5550 AVSS.n2929 AVSS.n2928 76.3222
R5551 AVSS.n2924 AVSS.n2921 76.3222
R5552 AVSS.n2922 AVSS.n1718 76.3222
R5553 AVSS.n4717 AVSS.n4716 76.3222
R5554 AVSS.n2939 AVSS.n2913 76.3222
R5555 AVSS.n2946 AVSS.n2945 76.3222
R5556 AVSS.n2947 AVSS.n2911 76.3222
R5557 AVSS.n2954 AVSS.n2953 76.3222
R5558 AVSS.n2958 AVSS.n2909 76.3222
R5559 AVSS.n2961 AVSS.n2960 76.3222
R5560 AVSS.n2967 AVSS.n2903 76.3222
R5561 AVSS.n2971 AVSS.n2904 76.3222
R5562 AVSS.n2975 AVSS.n2905 76.3222
R5563 AVSS.n2907 AVSS.n2906 76.3222
R5564 AVSS.n2981 AVSS.n2828 76.3222
R5565 AVSS.n4469 AVSS.n2808 76.3222
R5566 AVSS.n4715 AVSS.n1720 76.3222
R5567 AVSS.n2810 AVSS.n2803 76.3222
R5568 AVSS.n2814 AVSS.n2804 76.3222
R5569 AVSS.n2818 AVSS.n2805 76.3222
R5570 AVSS.n2822 AVSS.n2806 76.3222
R5571 AVSS.n4475 AVSS.n2807 76.3222
R5572 AVSS.n4475 AVSS.n4474 76.3222
R5573 AVSS.n2824 AVSS.n2806 76.3222
R5574 AVSS.n2821 AVSS.n2805 76.3222
R5575 AVSS.n2817 AVSS.n2804 76.3222
R5576 AVSS.n2813 AVSS.n2803 76.3222
R5577 AVSS.n2809 AVSS.n1720 76.3222
R5578 AVSS.n2940 AVSS.n2939 76.3222
R5579 AVSS.n2945 AVSS.n2944 76.3222
R5580 AVSS.n2948 AVSS.n2947 76.3222
R5581 AVSS.n2953 AVSS.n2952 76.3222
R5582 AVSS.n2955 AVSS.n2909 76.3222
R5583 AVSS.n2960 AVSS.n2959 76.3222
R5584 AVSS.n4718 AVSS.n4717 76.3222
R5585 AVSS.n2923 AVSS.n2922 76.3222
R5586 AVSS.n2921 AVSS.n2919 76.3222
R5587 AVSS.n2930 AVSS.n2929 76.3222
R5588 AVSS.n2918 AVSS.n2916 76.3222
R5589 AVSS.n2937 AVSS.n2936 76.3222
R5590 AVSS.n4686 AVSS.n4685 76.3222
R5591 AVSS.n1735 AVSS.n1733 76.3222
R5592 AVSS.n4693 AVSS.n4692 76.3222
R5593 AVSS.n1732 AVSS.n1730 76.3222
R5594 AVSS.n4700 AVSS.n4699 76.3222
R5595 AVSS.n1729 AVSS.n1727 76.3222
R5596 AVSS.n4506 AVSS.n4505 76.3222
R5597 AVSS.n2788 AVSS.n2786 76.3222
R5598 AVSS.n4513 AVSS.n4512 76.3222
R5599 AVSS.n2785 AVSS.n2783 76.3222
R5600 AVSS.n4520 AVSS.n4519 76.3222
R5601 AVSS.n2782 AVSS.n2780 76.3222
R5602 AVSS.n3238 AVSS.n3085 76.3222
R5603 AVSS.n3236 AVSS.n3235 76.3222
R5604 AVSS.n3231 AVSS.n3230 76.3222
R5605 AVSS.n3228 AVSS.n3227 76.3222
R5606 AVSS.n3223 AVSS.n3222 76.3222
R5607 AVSS.n3220 AVSS.n3219 76.3222
R5608 AVSS.n2159 AVSS.n1133 76.3222
R5609 AVSS.n2155 AVSS.n1134 76.3222
R5610 AVSS.n2151 AVSS.n1135 76.3222
R5611 AVSS.n2147 AVSS.n1136 76.3222
R5612 AVSS.n2143 AVSS.n1137 76.3222
R5613 AVSS.n2139 AVSS.n1138 76.3222
R5614 AVSS.n4935 AVSS.n4934 76.3222
R5615 AVSS.n4650 AVSS.n1131 76.3222
R5616 AVSS.n4654 AVSS.n1130 76.3222
R5617 AVSS.n4658 AVSS.n1129 76.3222
R5618 AVSS.n4662 AVSS.n1128 76.3222
R5619 AVSS.n4665 AVSS.n1127 76.3222
R5620 AVSS.n1350 AVSS.n1140 76.3222
R5621 AVSS.n1354 AVSS.n1141 76.3222
R5622 AVSS.n1358 AVSS.n1142 76.3222
R5623 AVSS.n1362 AVSS.n1143 76.3222
R5624 AVSS.n1146 AVSS.n1144 76.3222
R5625 AVSS.n1368 AVSS.n1145 76.3222
R5626 AVSS.n4754 AVSS.n4736 76.3222
R5627 AVSS.n4752 AVSS.n4751 76.3222
R5628 AVSS.n4747 AVSS.n4739 76.3222
R5629 AVSS.n4745 AVSS.n4744 76.3222
R5630 AVSS.n4740 AVSS.n1380 76.3222
R5631 AVSS.n4907 AVSS.n4906 76.3222
R5632 AVSS.n4911 AVSS.n1374 76.3222
R5633 AVSS.n4915 AVSS.n1375 76.3222
R5634 AVSS.n4919 AVSS.n1376 76.3222
R5635 AVSS.n1378 AVSS.n1377 76.3222
R5636 AVSS.n4925 AVSS.n1373 76.3222
R5637 AVSS.n4927 AVSS.n1370 76.3222
R5638 AVSS.n4785 AVSS.n1120 76.3222
R5639 AVSS.n4789 AVSS.n1121 76.3222
R5640 AVSS.n4793 AVSS.n1122 76.3222
R5641 AVSS.n4797 AVSS.n1123 76.3222
R5642 AVSS.n4801 AVSS.n1124 76.3222
R5643 AVSS.n4805 AVSS.n1125 76.3222
R5644 AVSS.n1369 AVSS.n1125 76.3222
R5645 AVSS.n4804 AVSS.n1124 76.3222
R5646 AVSS.n4800 AVSS.n1123 76.3222
R5647 AVSS.n4796 AVSS.n1122 76.3222
R5648 AVSS.n4792 AVSS.n1121 76.3222
R5649 AVSS.n4788 AVSS.n1120 76.3222
R5650 AVSS.n4928 AVSS.n4927 76.3222
R5651 AVSS.n4925 AVSS.n4924 76.3222
R5652 AVSS.n4920 AVSS.n1377 76.3222
R5653 AVSS.n4916 AVSS.n1376 76.3222
R5654 AVSS.n4912 AVSS.n1375 76.3222
R5655 AVSS.n4908 AVSS.n1374 76.3222
R5656 AVSS.n2117 AVSS.n2116 76.3222
R5657 AVSS.n2118 AVSS.n2087 76.3222
R5658 AVSS.n2125 AVSS.n2124 76.3222
R5659 AVSS.n2126 AVSS.n2085 76.3222
R5660 AVSS.n2133 AVSS.n2132 76.3222
R5661 AVSS.n2136 AVSS.n2135 76.3222
R5662 AVSS.n2162 AVSS.n2080 76.3222
R5663 AVSS.n2170 AVSS.n2169 76.3222
R5664 AVSS.n2079 AVSS.n2077 76.3222
R5665 AVSS.n2177 AVSS.n2176 76.3222
R5666 AVSS.n2076 AVSS.n2074 76.3222
R5667 AVSS.n2184 AVSS.n2183 76.3222
R5668 AVSS.n4627 AVSS.n4626 76.3222
R5669 AVSS.n4628 AVSS.n4622 76.3222
R5670 AVSS.n4635 AVSS.n4634 76.3222
R5671 AVSS.n4636 AVSS.n4620 76.3222
R5672 AVSS.n4643 AVSS.n4642 76.3222
R5673 AVSS.n4646 AVSS.n4645 76.3222
R5674 AVSS.n4941 AVSS.n4940 76.3222
R5675 AVSS.n1088 AVSS.n1086 76.3222
R5676 AVSS.n4948 AVSS.n4947 76.3222
R5677 AVSS.n1085 AVSS.n1083 76.3222
R5678 AVSS.n4955 AVSS.n4954 76.3222
R5679 AVSS.n1081 AVSS.n1079 76.3222
R5680 AVSS.n1194 AVSS.n1193 76.3222
R5681 AVSS.n1191 AVSS.n1190 76.3222
R5682 AVSS.n1186 AVSS.n1171 76.3222
R5683 AVSS.n1182 AVSS.n1170 76.3222
R5684 AVSS.n1178 AVSS.n1169 76.3222
R5685 AVSS.n1174 AVSS.n1168 76.3222
R5686 AVSS.n4906 AVSS.n4905 76.3222
R5687 AVSS.n4741 AVSS.n4740 76.3222
R5688 AVSS.n4746 AVSS.n4745 76.3222
R5689 AVSS.n4739 AVSS.n4737 76.3222
R5690 AVSS.n4753 AVSS.n4752 76.3222
R5691 AVSS.n4736 AVSS.n4734 76.3222
R5692 AVSS.n2187 AVSS.n2186 76.3222
R5693 AVSS.n2096 AVSS.n2095 76.3222
R5694 AVSS.n2101 AVSS.n2100 76.3222
R5695 AVSS.n2094 AVSS.n2092 76.3222
R5696 AVSS.n2108 AVSS.n2107 76.3222
R5697 AVSS.n2111 AVSS.n2110 76.3222
R5698 AVSS.n4962 AVSS.n4961 76.3222
R5699 AVSS.n1078 AVSS.n1076 76.3222
R5700 AVSS.n4969 AVSS.n4968 76.3222
R5701 AVSS.n1075 AVSS.n1073 76.3222
R5702 AVSS.n4976 AVSS.n4975 76.3222
R5703 AVSS.n4979 AVSS.n4978 76.3222
R5704 AVSS.n1314 AVSS.n1159 76.3222
R5705 AVSS.n1312 AVSS.n1311 76.3222
R5706 AVSS.n1307 AVSS.n1306 76.3222
R5707 AVSS.n1304 AVSS.n1303 76.3222
R5708 AVSS.n1299 AVSS.n1298 76.3222
R5709 AVSS.n1296 AVSS.n1295 76.3222
R5710 AVSS.n1591 AVSS.n667 76.3222
R5711 AVSS.n1495 AVSS.n666 76.3222
R5712 AVSS.n1499 AVSS.n665 76.3222
R5713 AVSS.n1503 AVSS.n664 76.3222
R5714 AVSS.n1507 AVSS.n663 76.3222
R5715 AVSS.n1510 AVSS.n662 76.3222
R5716 AVSS.n4990 AVSS.n4989 76.3222
R5717 AVSS.n947 AVSS.n887 76.3222
R5718 AVSS.n951 AVSS.n888 76.3222
R5719 AVSS.n955 AVSS.n889 76.3222
R5720 AVSS.n959 AVSS.n890 76.3222
R5721 AVSS.n893 AVSS.n891 76.3222
R5722 AVSS.n2317 AVSS.n660 76.3222
R5723 AVSS.n2321 AVSS.n659 76.3222
R5724 AVSS.n2325 AVSS.n658 76.3222
R5725 AVSS.n2329 AVSS.n657 76.3222
R5726 AVSS.n2333 AVSS.n656 76.3222
R5727 AVSS.n2336 AVSS.n655 76.3222
R5728 AVSS.n2227 AVSS.n965 76.3222
R5729 AVSS.n2223 AVSS.n966 76.3222
R5730 AVSS.n2219 AVSS.n967 76.3222
R5731 AVSS.n2215 AVSS.n968 76.3222
R5732 AVSS.n2211 AVSS.n969 76.3222
R5733 AVSS.n972 AVSS.n970 76.3222
R5734 AVSS.n718 AVSS.n653 76.3222
R5735 AVSS.n722 AVSS.n652 76.3222
R5736 AVSS.n726 AVSS.n651 76.3222
R5737 AVSS.n730 AVSS.n650 76.3222
R5738 AVSS.n734 AVSS.n649 76.3222
R5739 AVSS.n715 AVSS.n648 76.3222
R5740 AVSS.n2564 AVSS.n1742 76.3222
R5741 AVSS.n2568 AVSS.n1743 76.3222
R5742 AVSS.n2572 AVSS.n1744 76.3222
R5743 AVSS.n2575 AVSS.n1745 76.3222
R5744 AVSS.n2581 AVSS.n2580 76.3222
R5745 AVSS.n2584 AVSS.n2583 76.3222
R5746 AVSS.n1846 AVSS.n1113 76.3222
R5747 AVSS.n1841 AVSS.n1114 76.3222
R5748 AVSS.n1837 AVSS.n1115 76.3222
R5749 AVSS.n1833 AVSS.n1116 76.3222
R5750 AVSS.n1829 AVSS.n1117 76.3222
R5751 AVSS.n1825 AVSS.n1118 76.3222
R5752 AVSS.n2516 AVSS.n2515 76.3222
R5753 AVSS.n2519 AVSS.n2518 76.3222
R5754 AVSS.n2524 AVSS.n2523 76.3222
R5755 AVSS.n2527 AVSS.n2526 76.3222
R5756 AVSS.n2532 AVSS.n2531 76.3222
R5757 AVSS.n2535 AVSS.n2534 76.3222
R5758 AVSS.n1883 AVSS.n1853 76.3222
R5759 AVSS.n1882 AVSS.n1881 76.3222
R5760 AVSS.n1875 AVSS.n1855 76.3222
R5761 AVSS.n1874 AVSS.n1873 76.3222
R5762 AVSS.n1867 AVSS.n1857 76.3222
R5763 AVSS.n1866 AVSS.n1865 76.3222
R5764 AVSS.n1865 AVSS.n1864 76.3222
R5765 AVSS.n1868 AVSS.n1867 76.3222
R5766 AVSS.n1873 AVSS.n1872 76.3222
R5767 AVSS.n1876 AVSS.n1875 76.3222
R5768 AVSS.n1881 AVSS.n1880 76.3222
R5769 AVSS.n1884 AVSS.n1883 76.3222
R5770 AVSS.n2583 AVSS.n1741 76.3222
R5771 AVSS.n2581 AVSS.n1746 76.3222
R5772 AVSS.n2573 AVSS.n1745 76.3222
R5773 AVSS.n2569 AVSS.n1744 76.3222
R5774 AVSS.n2565 AVSS.n1743 76.3222
R5775 AVSS.n1859 AVSS.n1742 76.3222
R5776 AVSS.n2587 AVSS.n1118 76.3222
R5777 AVSS.n1826 AVSS.n1117 76.3222
R5778 AVSS.n1830 AVSS.n1116 76.3222
R5779 AVSS.n1834 AVSS.n1115 76.3222
R5780 AVSS.n1838 AVSS.n1114 76.3222
R5781 AVSS.n1842 AVSS.n1113 76.3222
R5782 AVSS.n2517 AVSS.n2516 76.3222
R5783 AVSS.n2518 AVSS.n1851 76.3222
R5784 AVSS.n2525 AVSS.n2524 76.3222
R5785 AVSS.n2526 AVSS.n1849 76.3222
R5786 AVSS.n2533 AVSS.n2532 76.3222
R5787 AVSS.n2536 AVSS.n2535 76.3222
R5788 AVSS.n4288 AVSS.n3894 76.3222
R5789 AVSS.n4286 AVSS.n4285 76.3222
R5790 AVSS.n4281 AVSS.n3897 76.3222
R5791 AVSS.n4279 AVSS.n4278 76.3222
R5792 AVSS.n4274 AVSS.n3900 76.3222
R5793 AVSS.n4272 AVSS.n4271 76.3222
R5794 AVSS.n4294 AVSS.n4293 76.3222
R5795 AVSS.n3923 AVSS.n3891 76.3222
R5796 AVSS.n3928 AVSS.n3927 76.3222
R5797 AVSS.n3931 AVSS.n3930 76.3222
R5798 AVSS.n3936 AVSS.n3935 76.3222
R5799 AVSS.n3939 AVSS.n3938 76.3222
R5800 AVSS.n3987 AVSS.n3901 76.3222
R5801 AVSS.n3986 AVSS.n3985 76.3222
R5802 AVSS.n3979 AVSS.n3903 76.3222
R5803 AVSS.n3978 AVSS.n3977 76.3222
R5804 AVSS.n3971 AVSS.n3905 76.3222
R5805 AVSS.n3970 AVSS.n3969 76.3222
R5806 AVSS.n3969 AVSS.n3968 76.3222
R5807 AVSS.n3972 AVSS.n3971 76.3222
R5808 AVSS.n3977 AVSS.n3976 76.3222
R5809 AVSS.n3980 AVSS.n3979 76.3222
R5810 AVSS.n3985 AVSS.n3984 76.3222
R5811 AVSS.n3988 AVSS.n3987 76.3222
R5812 AVSS.n4295 AVSS.n4294 76.3222
R5813 AVSS.n3924 AVSS.n3923 76.3222
R5814 AVSS.n3929 AVSS.n3928 76.3222
R5815 AVSS.n3930 AVSS.n3921 76.3222
R5816 AVSS.n3937 AVSS.n3936 76.3222
R5817 AVSS.n3940 AVSS.n3939 76.3222
R5818 AVSS.n4321 AVSS.n3683 76.3222
R5819 AVSS.n4319 AVSS.n4318 76.3222
R5820 AVSS.n4314 AVSS.n3686 76.3222
R5821 AVSS.n4312 AVSS.n4311 76.3222
R5822 AVSS.n4307 AVSS.n3689 76.3222
R5823 AVSS.n4305 AVSS.n4304 76.3222
R5824 AVSS.n4327 AVSS.n4326 76.3222
R5825 AVSS.n3712 AVSS.n3680 76.3222
R5826 AVSS.n3717 AVSS.n3716 76.3222
R5827 AVSS.n3720 AVSS.n3719 76.3222
R5828 AVSS.n3725 AVSS.n3724 76.3222
R5829 AVSS.n3728 AVSS.n3727 76.3222
R5830 AVSS.n3776 AVSS.n3690 76.3222
R5831 AVSS.n3775 AVSS.n3774 76.3222
R5832 AVSS.n3768 AVSS.n3692 76.3222
R5833 AVSS.n3767 AVSS.n3766 76.3222
R5834 AVSS.n3760 AVSS.n3694 76.3222
R5835 AVSS.n3759 AVSS.n3758 76.3222
R5836 AVSS.n3758 AVSS.n3757 76.3222
R5837 AVSS.n3761 AVSS.n3760 76.3222
R5838 AVSS.n3766 AVSS.n3765 76.3222
R5839 AVSS.n3769 AVSS.n3768 76.3222
R5840 AVSS.n3774 AVSS.n3773 76.3222
R5841 AVSS.n3777 AVSS.n3776 76.3222
R5842 AVSS.n4328 AVSS.n4327 76.3222
R5843 AVSS.n3713 AVSS.n3712 76.3222
R5844 AVSS.n3718 AVSS.n3717 76.3222
R5845 AVSS.n3719 AVSS.n3710 76.3222
R5846 AVSS.n3726 AVSS.n3725 76.3222
R5847 AVSS.n3729 AVSS.n3728 76.3222
R5848 AVSS.n3558 AVSS.n3557 76.3222
R5849 AVSS.n3553 AVSS.n3540 76.3222
R5850 AVSS.n3551 AVSS.n3550 76.3222
R5851 AVSS.n3546 AVSS.n3543 76.3222
R5852 AVSS.n3544 AVSS.n3513 76.3222
R5853 AVSS.n4338 AVSS.n4337 76.3222
R5854 AVSS.n4336 AVSS.n3514 76.3222
R5855 AVSS.n3638 AVSS.n3637 76.3222
R5856 AVSS.n3631 AVSS.n3516 76.3222
R5857 AVSS.n3630 AVSS.n3629 76.3222
R5858 AVSS.n3623 AVSS.n3518 76.3222
R5859 AVSS.n3622 AVSS.n3621 76.3222
R5860 AVSS.n3621 AVSS.n3620 76.3222
R5861 AVSS.n3624 AVSS.n3623 76.3222
R5862 AVSS.n3629 AVSS.n3628 76.3222
R5863 AVSS.n3632 AVSS.n3631 76.3222
R5864 AVSS.n3637 AVSS.n3636 76.3222
R5865 AVSS.n3639 AVSS.n3514 76.3222
R5866 AVSS.n4339 AVSS.n4338 76.3222
R5867 AVSS.n3545 AVSS.n3544 76.3222
R5868 AVSS.n3543 AVSS.n3541 76.3222
R5869 AVSS.n3552 AVSS.n3551 76.3222
R5870 AVSS.n3540 AVSS.n3538 76.3222
R5871 AVSS.n3559 AVSS.n3558 76.3222
R5872 AVSS.n4306 AVSS.n4305 76.3222
R5873 AVSS.n3689 AVSS.n3687 76.3222
R5874 AVSS.n4313 AVSS.n4312 76.3222
R5875 AVSS.n3686 AVSS.n3684 76.3222
R5876 AVSS.n4320 AVSS.n4319 76.3222
R5877 AVSS.n3683 AVSS.n3681 76.3222
R5878 AVSS.n4273 AVSS.n4272 76.3222
R5879 AVSS.n3900 AVSS.n3898 76.3222
R5880 AVSS.n4280 AVSS.n4279 76.3222
R5881 AVSS.n3897 AVSS.n3895 76.3222
R5882 AVSS.n4287 AVSS.n4286 76.3222
R5883 AVSS.n3894 AVSS.n3892 76.3222
R5884 AVSS.n6193 AVSS.n6192 76.3222
R5885 AVSS.n157 AVSS.n155 76.3222
R5886 AVSS.n6200 AVSS.n6199 76.3222
R5887 AVSS.n154 AVSS.n152 76.3222
R5888 AVSS.n6207 AVSS.n6206 76.3222
R5889 AVSS.n256 AVSS.n150 76.3222
R5890 AVSS.n4470 AVSS.n4469 76.3222
R5891 AVSS.n2981 AVSS.n2980 76.3222
R5892 AVSS.n2976 AVSS.n2906 76.3222
R5893 AVSS.n2972 AVSS.n2905 76.3222
R5894 AVSS.n2968 AVSS.n2904 76.3222
R5895 AVSS.n2964 AVSS.n2903 76.3222
R5896 AVSS.n3043 AVSS.n2983 76.3222
R5897 AVSS.n3047 AVSS.n2984 76.3222
R5898 AVSS.n3051 AVSS.n2985 76.3222
R5899 AVSS.n3055 AVSS.n2986 76.3222
R5900 AVSS.n3059 AVSS.n2987 76.3222
R5901 AVSS.n2990 AVSS.n2988 76.3222
R5902 AVSS.n2901 AVSS.n2835 76.3222
R5903 AVSS.n2877 AVSS.n2834 76.3222
R5904 AVSS.n2873 AVSS.n2833 76.3222
R5905 AVSS.n2869 AVSS.n2832 76.3222
R5906 AVSS.n2865 AVSS.n2831 76.3222
R5907 AVSS.n2861 AVSS.n2830 76.3222
R5908 AVSS.n3275 AVSS.n3065 76.3222
R5909 AVSS.n3279 AVSS.n3066 76.3222
R5910 AVSS.n3283 AVSS.n3067 76.3222
R5911 AVSS.n3287 AVSS.n3068 76.3222
R5912 AVSS.n3071 AVSS.n3069 76.3222
R5913 AVSS.n3293 AVSS.n3070 76.3222
R5914 AVSS.n6090 AVSS.n6089 76.3222
R5915 AVSS.n6091 AVSS.n227 76.3222
R5916 AVSS.n6098 AVSS.n6097 76.3222
R5917 AVSS.n6099 AVSS.n225 76.3222
R5918 AVSS.n6106 AVSS.n6105 76.3222
R5919 AVSS.n6107 AVSS.n223 76.3222
R5920 AVSS.n4261 AVSS.n4260 76.3222
R5921 AVSS.n4229 AVSS.n4228 76.3222
R5922 AVSS.n4222 AVSS.n4208 76.3222
R5923 AVSS.n4221 AVSS.n4220 76.3222
R5924 AVSS.n4214 AVSS.n4210 76.3222
R5925 AVSS.n4213 AVSS.n4212 76.3222
R5926 AVSS.n4259 AVSS.n4230 76.3222
R5927 AVSS.n4255 AVSS.n4254 76.3222
R5928 AVSS.n4248 AVSS.n4232 76.3222
R5929 AVSS.n4247 AVSS.n4246 76.3222
R5930 AVSS.n4240 AVSS.n4234 76.3222
R5931 AVSS.n4239 AVSS.n4238 76.3222
R5932 AVSS.n4238 AVSS.n4237 76.3222
R5933 AVSS.n4241 AVSS.n4240 76.3222
R5934 AVSS.n4246 AVSS.n4245 76.3222
R5935 AVSS.n4249 AVSS.n4248 76.3222
R5936 AVSS.n4254 AVSS.n4253 76.3222
R5937 AVSS.n4256 AVSS.n4230 76.3222
R5938 AVSS.n4262 AVSS.n4261 76.3222
R5939 AVSS.n4228 AVSS.n4227 76.3222
R5940 AVSS.n4223 AVSS.n4222 76.3222
R5941 AVSS.n4220 AVSS.n4219 76.3222
R5942 AVSS.n4215 AVSS.n4214 76.3222
R5943 AVSS.n4212 AVSS.n211 76.3222
R5944 AVSS.n6108 AVSS.n6107 76.3222
R5945 AVSS.n6105 AVSS.n6104 76.3222
R5946 AVSS.n6100 AVSS.n6099 76.3222
R5947 AVSS.n6097 AVSS.n6096 76.3222
R5948 AVSS.n6092 AVSS.n6091 76.3222
R5949 AVSS.n6089 AVSS.n6088 76.3222
R5950 AVSS.n259 AVSS.n258 76.3222
R5951 AVSS.n254 AVSS.n253 76.3222
R5952 AVSS.n249 AVSS.n248 76.3222
R5953 AVSS.n246 AVSS.n245 76.3222
R5954 AVSS.n241 AVSS.n240 76.3222
R5955 AVSS.n238 AVSS.n186 76.3222
R5956 AVSS.n4394 AVSS.n4357 76.3222
R5957 AVSS.n4401 AVSS.n4400 76.3222
R5958 AVSS.n4402 AVSS.n4355 76.3222
R5959 AVSS.n4409 AVSS.n4408 76.3222
R5960 AVSS.n4410 AVSS.n4353 76.3222
R5961 AVSS.n4418 AVSS.n4417 76.3222
R5962 AVSS.n4419 AVSS.n4351 76.3222
R5963 AVSS.n4426 AVSS.n4425 76.3222
R5964 AVSS.n4427 AVSS.n4349 76.3222
R5965 AVSS.n4434 AVSS.n4433 76.3222
R5966 AVSS.n4435 AVSS.n4347 76.3222
R5967 AVSS.n4442 AVSS.n4441 76.3222
R5968 AVSS.n4463 AVSS.n3299 76.3222
R5969 AVSS.n4459 AVSS.n3298 76.3222
R5970 AVSS.n4455 AVSS.n3297 76.3222
R5971 AVSS.n4451 AVSS.n3296 76.3222
R5972 AVSS.n4447 AVSS.n3295 76.3222
R5973 AVSS.n4443 AVSS.n3294 76.3222
R5974 AVSS.n4417 AVSS.n4416 76.3222
R5975 AVSS.n4411 AVSS.n4410 76.3222
R5976 AVSS.n4408 AVSS.n4407 76.3222
R5977 AVSS.n4403 AVSS.n4402 76.3222
R5978 AVSS.n4400 AVSS.n4399 76.3222
R5979 AVSS.n4395 AVSS.n4394 76.3222
R5980 AVSS.n4441 AVSS.n4440 76.3222
R5981 AVSS.n4436 AVSS.n4435 76.3222
R5982 AVSS.n4433 AVSS.n4432 76.3222
R5983 AVSS.n4428 AVSS.n4427 76.3222
R5984 AVSS.n4425 AVSS.n4424 76.3222
R5985 AVSS.n4420 AVSS.n4419 76.3222
R5986 AVSS.n4446 AVSS.n3294 76.3222
R5987 AVSS.n4450 AVSS.n3295 76.3222
R5988 AVSS.n4454 AVSS.n3296 76.3222
R5989 AVSS.n4458 AVSS.n3297 76.3222
R5990 AVSS.n4462 AVSS.n3298 76.3222
R5991 AVSS.n3301 AVSS.n3299 76.3222
R5992 AVSS.n135 AVSS.n72 76.062
R5993 AVSS.n137 AVSS.n72 76.062
R5994 AVSS.n4187 AVSS.n4131 76.062
R5995 AVSS.n4184 AVSS.n4131 76.062
R5996 AVSS.n4045 AVSS.n4044 76.062
R5997 AVSS.n4044 AVSS.n4043 76.062
R5998 AVSS.n3834 AVSS.n3833 76.062
R5999 AVSS.n3833 AVSS.n3832 76.062
R6000 AVSS.n3475 AVSS.n3474 76.062
R6001 AVSS.n3474 AVSS.n3473 76.062
R6002 AVSS.n5815 AVSS.n5729 76.062
R6003 AVSS.n5798 AVSS.n5729 76.062
R6004 AVSS.n5543 AVSS.n5457 76.062
R6005 AVSS.n5526 AVSS.n5457 76.062
R6006 AVSS.n5372 AVSS.n5371 76.062
R6007 AVSS.n5371 AVSS.n5307 76.062
R6008 AVSS.n5173 AVSS.n5172 76.062
R6009 AVSS.n5172 AVSS.n5108 76.062
R6010 AVSS.n3210 AVSS.n3209 76.062
R6011 AVSS.n3210 AVSS.n3143 76.062
R6012 AVSS.n1286 AVSS.n1285 76.062
R6013 AVSS.n1286 AVSS.n1219 76.062
R6014 AVSS.n4613 AVSS.n4526 76.062
R6015 AVSS.n4596 AVSS.n4526 76.062
R6016 AVSS.n2763 AVSS.n2700 76.062
R6017 AVSS.n2765 AVSS.n2700 76.062
R6018 AVSS.n2647 AVSS.n2646 76.062
R6019 AVSS.n2646 AVSS.n2645 76.062
R6020 AVSS.n1680 AVSS.n1679 76.062
R6021 AVSS.n1679 AVSS.n1678 76.062
R6022 AVSS.n827 AVSS.n826 76.062
R6023 AVSS.n827 AVSS.n760 76.062
R6024 AVSS.n1063 AVSS.n977 76.062
R6025 AVSS.n1046 AVSS.n977 76.062
R6026 AVSS.n2505 AVSS.n2504 76.062
R6027 AVSS.n2506 AVSS.n2505 76.062
R6028 AVSS.n2542 AVSS.n1766 76.062
R6029 AVSS.n1821 AVSS.n1766 76.062
R6030 AVSS.n5992 AVSS.t10 74.6623
R6031 AVSS.n518 AVSS.n477 74.5978
R6032 AVSS.n515 AVSS.n477 74.5978
R6033 AVSS.n1427 AVSS.n1405 74.5978
R6034 AVSS.n1424 AVSS.n1405 74.5978
R6035 AVSS.n4847 AVSS.n4825 74.5978
R6036 AVSS.n4844 AVSS.n4825 74.5978
R6037 AVSS.n2014 AVSS.n1992 74.5978
R6038 AVSS.n2011 AVSS.n1992 74.5978
R6039 AVSS.n1942 AVSS.n1901 74.5978
R6040 AVSS.n1939 AVSS.n1901 74.5978
R6041 AVSS.n3361 AVSS.n3319 74.5978
R6042 AVSS.n3358 AVSS.n3319 74.5978
R6043 AVSS.n3885 AVSS.n3872 73.3165
R6044 AVSS.n4096 AVSS.n4083 73.3165
R6045 AVSS.n4103 AVSS.n4102 73.3165
R6046 AVSS.n3649 AVSS.n3648 73.3165
R6047 AVSS.n3413 AVSS.n3412 73.3165
R6048 AVSS.n1616 AVSS.n1615 73.3165
R6049 AVSS.n5021 AVSS.n5020 73.3165
R6050 AVSS.n5040 AVSS.n454 73.3165
R6051 AVSS.n583 AVSS.n572 73.3165
R6052 AVSS.n1104 AVSS.n1093 73.3165
R6053 AVSS.n4489 AVSS.n4478 73.3165
R6054 AVSS.n6230 AVSS.n38 73.3165
R6055 AVSS.n6246 AVSS.n6245 73.3165
R6056 AVSS.n6259 AVSS.n21 73.3165
R6057 AVSS.n5058 AVSS.n450 73.3165
R6058 AVSS.n269 AVSS.n268 73.3165
R6059 AVSS.n3876 AVSS.n187 73.19
R6060 AVSS.n4087 AVSS.n189 73.19
R6061 AVSS.n4111 AVSS.n191 73.19
R6062 AVSS.n3664 AVSS.n193 73.19
R6063 AVSS.n3403 AVSS.n2797 73.19
R6064 AVSS.n1603 AVSS.n1602 73.19
R6065 AVSS.n570 AVSS.n561 73.19
R6066 AVSS.n5031 AVSS.n5030 73.19
R6067 AVSS.n586 AVSS.n571 73.19
R6068 AVSS.n1107 AVSS.n1092 73.19
R6069 AVSS.n4492 AVSS.n4477 73.19
R6070 AVSS.n6237 AVSS.n33 73.19
R6071 AVSS.n6254 AVSS.n26 73.19
R6072 AVSS.n5053 AVSS.n20 73.19
R6073 AVSS.n5045 AVSS.n449 73.19
R6074 AVSS.n277 AVSS.n195 73.19
R6075 AVSS.t10 AVSS 70.6265
R6076 AVSS.n4169 AVSS.n4125 69.3109
R6077 AVSS.n4167 AVSS.n4125 69.3109
R6078 AVSS.n4028 AVSS.n4006 69.3109
R6079 AVSS.n4025 AVSS.n4006 69.3109
R6080 AVSS.n3817 AVSS.n3795 69.3109
R6081 AVSS.n3814 AVSS.n3795 69.3109
R6082 AVSS.n3458 AVSS.n3436 69.3109
R6083 AVSS.n3455 AVSS.n3436 69.3109
R6084 AVSS.n549 AVSS.n548 69.3109
R6085 AVSS.n548 AVSS.n465 69.3109
R6086 AVSS.n1461 AVSS.n1401 69.3109
R6087 AVSS.n1457 AVSS.n1401 69.3109
R6088 AVSS.n4881 AVSS.n4821 69.3109
R6089 AVSS.n4877 AVSS.n4821 69.3109
R6090 AVSS.n2630 AVSS.n2608 69.3109
R6091 AVSS.n2627 AVSS.n2608 69.3109
R6092 AVSS.n1663 AVSS.n1641 69.3109
R6093 AVSS.n1660 AVSS.n1641 69.3109
R6094 AVSS.n2048 AVSS.n1988 69.3109
R6095 AVSS.n2044 AVSS.n1988 69.3109
R6096 AVSS.n1973 AVSS.n1972 69.3109
R6097 AVSS.n1972 AVSS.n1889 69.3109
R6098 AVSS.n3392 AVSS.n3391 69.3109
R6099 AVSS.n3391 AVSS.n3307 69.3109
R6100 AVSS.n5873 AVSS.n399 67.477
R6101 AVSS.n4933 AVSS.n1132 67.477
R6102 AVSS.n4988 AVSS.n886 67.477
R6103 AVSS.n4468 AVSS.n2982 67.477
R6104 AVSS.n3606 AVSS.t110 67.1938
R6105 AVSS.n3743 AVSS.t108 67.1938
R6106 AVSS.n3954 AVSS.t95 67.1938
R6107 AVSS.n6123 AVSS.t102 67.1938
R6108 AVSS.t85 AVSS.n168 67.1938
R6109 AVSS.n5016 AVSS.n399 66.8089
R6110 AVSS.n1719 AVSS.n1132 66.8089
R6111 AVSS.n1071 AVSS.n886 66.8089
R6112 AVSS.n2982 AVSS.n151 66.8089
R6113 AVSS.n5952 AVSS.n5951 66.3172
R6114 AVSS.n5950 AVSS.n5949 66.3172
R6115 AVSS.t83 AVSS.n73 65.8183
R6116 AVSS.t83 AVSS.n74 65.8183
R6117 AVSS.t83 AVSS.n75 65.8183
R6118 AVSS.t83 AVSS.n142 65.8183
R6119 AVSS.t83 AVSS.n62 65.8183
R6120 AVSS.t83 AVSS.n61 65.8183
R6121 AVSS.t83 AVSS.n69 65.8183
R6122 AVSS.t83 AVSS.n60 65.8183
R6123 AVSS.t83 AVSS.n66 65.8183
R6124 AVSS.t83 AVSS.n65 65.8183
R6125 AVSS.t83 AVSS.n64 65.8183
R6126 AVSS.t83 AVSS.n63 65.8183
R6127 AVSS.t83 AVSS.n68 65.8183
R6128 AVSS.t83 AVSS.n70 65.8183
R6129 AVSS.t83 AVSS.n71 65.8183
R6130 AVSS.n143 AVSS.t83 65.8183
R6131 AVSS.t101 AVSS.n4129 65.8183
R6132 AVSS.t101 AVSS.n4128 65.8183
R6133 AVSS.t101 AVSS.n4127 65.8183
R6134 AVSS.t101 AVSS.n4126 65.8183
R6135 AVSS.t101 AVSS.n4122 65.8183
R6136 AVSS.t101 AVSS.n4130 65.8183
R6137 AVSS.t101 AVSS.n4119 65.8183
R6138 AVSS.t101 AVSS.n4201 65.8183
R6139 AVSS.t101 AVSS.n4134 65.8183
R6140 AVSS.t101 AVSS.n4133 65.8183
R6141 AVSS.t101 AVSS.n4132 65.8183
R6142 AVSS.t101 AVSS.n4123 65.8183
R6143 AVSS.t101 AVSS.n4121 65.8183
R6144 AVSS.t101 AVSS.n4120 65.8183
R6145 AVSS.t101 AVSS.n4118 65.8183
R6146 AVSS.n4023 AVSS.t94 65.8183
R6147 AVSS.n4017 AVSS.t94 65.8183
R6148 AVSS.n4015 AVSS.t94 65.8183
R6149 AVSS.n4010 AVSS.t94 65.8183
R6150 AVSS.n4030 AVSS.t94 65.8183
R6151 AVSS.n4036 AVSS.t94 65.8183
R6152 AVSS.n4038 AVSS.t94 65.8183
R6153 AVSS.n4059 AVSS.t94 65.8183
R6154 AVSS.n3998 AVSS.t94 65.8183
R6155 AVSS.n4052 AVSS.t94 65.8183
R6156 AVSS.n4046 AVSS.t94 65.8183
R6157 AVSS.n4077 AVSS.t94 65.8183
R6158 AVSS.n4074 AVSS.t94 65.8183
R6159 AVSS.n4068 AVSS.t94 65.8183
R6160 AVSS.n4066 AVSS.t94 65.8183
R6161 AVSS.n3812 AVSS.t107 65.8183
R6162 AVSS.n3806 AVSS.t107 65.8183
R6163 AVSS.n3804 AVSS.t107 65.8183
R6164 AVSS.n3799 AVSS.t107 65.8183
R6165 AVSS.n3819 AVSS.t107 65.8183
R6166 AVSS.n3825 AVSS.t107 65.8183
R6167 AVSS.n3827 AVSS.t107 65.8183
R6168 AVSS.n3848 AVSS.t107 65.8183
R6169 AVSS.n3787 AVSS.t107 65.8183
R6170 AVSS.n3841 AVSS.t107 65.8183
R6171 AVSS.n3835 AVSS.t107 65.8183
R6172 AVSS.n3866 AVSS.t107 65.8183
R6173 AVSS.n3863 AVSS.t107 65.8183
R6174 AVSS.n3857 AVSS.t107 65.8183
R6175 AVSS.n3855 AVSS.t107 65.8183
R6176 AVSS.n3453 AVSS.t109 65.8183
R6177 AVSS.n3447 AVSS.t109 65.8183
R6178 AVSS.n3445 AVSS.t109 65.8183
R6179 AVSS.n3440 AVSS.t109 65.8183
R6180 AVSS.n3460 AVSS.t109 65.8183
R6181 AVSS.n3466 AVSS.t109 65.8183
R6182 AVSS.n3468 AVSS.t109 65.8183
R6183 AVSS.n3489 AVSS.t109 65.8183
R6184 AVSS.n3428 AVSS.t109 65.8183
R6185 AVSS.n3482 AVSS.t109 65.8183
R6186 AVSS.n3476 AVSS.t109 65.8183
R6187 AVSS.n3506 AVSS.t109 65.8183
R6188 AVSS.n3503 AVSS.t109 65.8183
R6189 AVSS.n3497 AVSS.t109 65.8183
R6190 AVSS.n3495 AVSS.t109 65.8183
R6191 AVSS.t105 AVSS.n5812 65.8183
R6192 AVSS.t105 AVSS.n5745 65.8183
R6193 AVSS.t105 AVSS.n5744 65.8183
R6194 AVSS.t105 AVSS.n5743 65.8183
R6195 AVSS.t105 AVSS.n5735 65.8183
R6196 AVSS.t105 AVSS.n5733 65.8183
R6197 AVSS.t105 AVSS.n5731 65.8183
R6198 AVSS.t105 AVSS.n5742 65.8183
R6199 AVSS.t105 AVSS.n5741 65.8183
R6200 AVSS.t105 AVSS.n5740 65.8183
R6201 AVSS.t105 AVSS.n5739 65.8183
R6202 AVSS.t105 AVSS.n5738 65.8183
R6203 AVSS.t105 AVSS.n5736 65.8183
R6204 AVSS.t105 AVSS.n5734 65.8183
R6205 AVSS.t105 AVSS.n5732 65.8183
R6206 AVSS.n5813 AVSS.t105 65.8183
R6207 AVSS.t91 AVSS.n5540 65.8183
R6208 AVSS.t91 AVSS.n5473 65.8183
R6209 AVSS.t91 AVSS.n5472 65.8183
R6210 AVSS.t91 AVSS.n5471 65.8183
R6211 AVSS.t91 AVSS.n5463 65.8183
R6212 AVSS.t91 AVSS.n5461 65.8183
R6213 AVSS.t91 AVSS.n5459 65.8183
R6214 AVSS.t91 AVSS.n5470 65.8183
R6215 AVSS.t91 AVSS.n5469 65.8183
R6216 AVSS.t91 AVSS.n5468 65.8183
R6217 AVSS.t91 AVSS.n5467 65.8183
R6218 AVSS.t91 AVSS.n5466 65.8183
R6219 AVSS.t91 AVSS.n5464 65.8183
R6220 AVSS.t91 AVSS.n5462 65.8183
R6221 AVSS.t91 AVSS.n5460 65.8183
R6222 AVSS.n5541 AVSS.t91 65.8183
R6223 AVSS.n5355 AVSS.t88 65.8183
R6224 AVSS.n5361 AVSS.t88 65.8183
R6225 AVSS.n5363 AVSS.t88 65.8183
R6226 AVSS.n5369 AVSS.t88 65.8183
R6227 AVSS.n5339 AVSS.t88 65.8183
R6228 AVSS.n5345 AVSS.t88 65.8183
R6229 AVSS.n5347 AVSS.t88 65.8183
R6230 AVSS.n5353 AVSS.t88 65.8183
R6231 AVSS.n5323 AVSS.t88 65.8183
R6232 AVSS.n5322 AVSS.t88 65.8183
R6233 AVSS.n5330 AVSS.t88 65.8183
R6234 AVSS.n5319 AVSS.t88 65.8183
R6235 AVSS.n5389 AVSS.t88 65.8183
R6236 AVSS.n5386 AVSS.t88 65.8183
R6237 AVSS.n5380 AVSS.t88 65.8183
R6238 AVSS.n5378 AVSS.t88 65.8183
R6239 AVSS.n5156 AVSS.t98 65.8183
R6240 AVSS.n5162 AVSS.t98 65.8183
R6241 AVSS.n5164 AVSS.t98 65.8183
R6242 AVSS.n5170 AVSS.t98 65.8183
R6243 AVSS.n5140 AVSS.t98 65.8183
R6244 AVSS.n5146 AVSS.t98 65.8183
R6245 AVSS.n5148 AVSS.t98 65.8183
R6246 AVSS.n5154 AVSS.t98 65.8183
R6247 AVSS.n5124 AVSS.t98 65.8183
R6248 AVSS.n5123 AVSS.t98 65.8183
R6249 AVSS.n5131 AVSS.t98 65.8183
R6250 AVSS.n5120 AVSS.t98 65.8183
R6251 AVSS.n5190 AVSS.t98 65.8183
R6252 AVSS.n5187 AVSS.t98 65.8183
R6253 AVSS.n5181 AVSS.t98 65.8183
R6254 AVSS.n5179 AVSS.t98 65.8183
R6255 AVSS.t103 AVSS.n470 65.8183
R6256 AVSS.t103 AVSS.n471 65.8183
R6257 AVSS.t103 AVSS.n472 65.8183
R6258 AVSS.t103 AVSS.n473 65.8183
R6259 AVSS.t103 AVSS.n468 65.8183
R6260 AVSS.t103 AVSS.n467 65.8183
R6261 AVSS.t103 AVSS.n466 65.8183
R6262 AVSS.t103 AVSS.n478 65.8183
R6263 AVSS.t103 AVSS.n479 65.8183
R6264 AVSS.t103 AVSS.n480 65.8183
R6265 AVSS.t103 AVSS.n481 65.8183
R6266 AVSS.t103 AVSS.n474 65.8183
R6267 AVSS.t103 AVSS.n475 65.8183
R6268 AVSS.t103 AVSS.n476 65.8183
R6269 AVSS.t103 AVSS.n547 65.8183
R6270 AVSS.t86 AVSS.n1397 65.8183
R6271 AVSS.t86 AVSS.n1398 65.8183
R6272 AVSS.t86 AVSS.n1399 65.8183
R6273 AVSS.t86 AVSS.n1400 65.8183
R6274 AVSS.t86 AVSS.n1396 65.8183
R6275 AVSS.t86 AVSS.n1395 65.8183
R6276 AVSS.t86 AVSS.n1394 65.8183
R6277 AVSS.t86 AVSS.n1406 65.8183
R6278 AVSS.t86 AVSS.n1407 65.8183
R6279 AVSS.t86 AVSS.n1408 65.8183
R6280 AVSS.t86 AVSS.n1409 65.8183
R6281 AVSS.t86 AVSS.n1402 65.8183
R6282 AVSS.t86 AVSS.n1403 65.8183
R6283 AVSS.t86 AVSS.n1404 65.8183
R6284 AVSS.t86 AVSS.n1477 65.8183
R6285 AVSS.t93 AVSS.n4817 65.8183
R6286 AVSS.t93 AVSS.n4818 65.8183
R6287 AVSS.t93 AVSS.n4819 65.8183
R6288 AVSS.t93 AVSS.n4820 65.8183
R6289 AVSS.t93 AVSS.n4816 65.8183
R6290 AVSS.t93 AVSS.n4815 65.8183
R6291 AVSS.t93 AVSS.n4814 65.8183
R6292 AVSS.t93 AVSS.n4826 65.8183
R6293 AVSS.t93 AVSS.n4827 65.8183
R6294 AVSS.t93 AVSS.n4828 65.8183
R6295 AVSS.t93 AVSS.n4829 65.8183
R6296 AVSS.t93 AVSS.n4822 65.8183
R6297 AVSS.t93 AVSS.n4823 65.8183
R6298 AVSS.t93 AVSS.n4824 65.8183
R6299 AVSS.t93 AVSS.n4897 65.8183
R6300 AVSS.t100 AVSS.n3142 65.8183
R6301 AVSS.t100 AVSS.n3141 65.8183
R6302 AVSS.t100 AVSS.n3140 65.8183
R6303 AVSS.t100 AVSS.n3139 65.8183
R6304 AVSS.t100 AVSS.n3132 65.8183
R6305 AVSS.t100 AVSS.n3130 65.8183
R6306 AVSS.t100 AVSS.n3128 65.8183
R6307 AVSS.n3211 AVSS.t100 65.8183
R6308 AVSS.t100 AVSS.n3138 65.8183
R6309 AVSS.t100 AVSS.n3137 65.8183
R6310 AVSS.t100 AVSS.n3136 65.8183
R6311 AVSS.t100 AVSS.n3135 65.8183
R6312 AVSS.t100 AVSS.n3133 65.8183
R6313 AVSS.t100 AVSS.n3131 65.8183
R6314 AVSS.t100 AVSS.n3129 65.8183
R6315 AVSS.t100 AVSS.n3127 65.8183
R6316 AVSS.t96 AVSS.n1218 65.8183
R6317 AVSS.t96 AVSS.n1217 65.8183
R6318 AVSS.t96 AVSS.n1216 65.8183
R6319 AVSS.t96 AVSS.n1215 65.8183
R6320 AVSS.t96 AVSS.n1208 65.8183
R6321 AVSS.t96 AVSS.n1206 65.8183
R6322 AVSS.t96 AVSS.n1204 65.8183
R6323 AVSS.n1287 AVSS.t96 65.8183
R6324 AVSS.t96 AVSS.n1214 65.8183
R6325 AVSS.t96 AVSS.n1213 65.8183
R6326 AVSS.t96 AVSS.n1212 65.8183
R6327 AVSS.t96 AVSS.n1211 65.8183
R6328 AVSS.t96 AVSS.n1209 65.8183
R6329 AVSS.t96 AVSS.n1207 65.8183
R6330 AVSS.t96 AVSS.n1205 65.8183
R6331 AVSS.t96 AVSS.n1203 65.8183
R6332 AVSS.t112 AVSS.n4610 65.8183
R6333 AVSS.t112 AVSS.n4542 65.8183
R6334 AVSS.t112 AVSS.n4541 65.8183
R6335 AVSS.t112 AVSS.n4540 65.8183
R6336 AVSS.t112 AVSS.n4532 65.8183
R6337 AVSS.t112 AVSS.n4530 65.8183
R6338 AVSS.t112 AVSS.n4528 65.8183
R6339 AVSS.t112 AVSS.n4539 65.8183
R6340 AVSS.t112 AVSS.n4538 65.8183
R6341 AVSS.t112 AVSS.n4537 65.8183
R6342 AVSS.t112 AVSS.n4536 65.8183
R6343 AVSS.t112 AVSS.n4535 65.8183
R6344 AVSS.t112 AVSS.n4533 65.8183
R6345 AVSS.t112 AVSS.n4531 65.8183
R6346 AVSS.t112 AVSS.n4529 65.8183
R6347 AVSS.n4611 AVSS.t112 65.8183
R6348 AVSS.t75 AVSS.n2701 65.8183
R6349 AVSS.t75 AVSS.n2702 65.8183
R6350 AVSS.t75 AVSS.n2703 65.8183
R6351 AVSS.t75 AVSS.n2770 65.8183
R6352 AVSS.t75 AVSS.n2690 65.8183
R6353 AVSS.t75 AVSS.n2689 65.8183
R6354 AVSS.t75 AVSS.n2697 65.8183
R6355 AVSS.t75 AVSS.n2688 65.8183
R6356 AVSS.t75 AVSS.n2694 65.8183
R6357 AVSS.t75 AVSS.n2693 65.8183
R6358 AVSS.t75 AVSS.n2692 65.8183
R6359 AVSS.t75 AVSS.n2691 65.8183
R6360 AVSS.t75 AVSS.n2696 65.8183
R6361 AVSS.t75 AVSS.n2698 65.8183
R6362 AVSS.t75 AVSS.n2699 65.8183
R6363 AVSS.n2771 AVSS.t75 65.8183
R6364 AVSS.n2625 AVSS.t111 65.8183
R6365 AVSS.n2619 AVSS.t111 65.8183
R6366 AVSS.n2617 AVSS.t111 65.8183
R6367 AVSS.n2612 AVSS.t111 65.8183
R6368 AVSS.n2632 AVSS.t111 65.8183
R6369 AVSS.n2638 AVSS.t111 65.8183
R6370 AVSS.n2640 AVSS.t111 65.8183
R6371 AVSS.n2661 AVSS.t111 65.8183
R6372 AVSS.n2600 AVSS.t111 65.8183
R6373 AVSS.n2654 AVSS.t111 65.8183
R6374 AVSS.n2648 AVSS.t111 65.8183
R6375 AVSS.n2679 AVSS.t111 65.8183
R6376 AVSS.n2676 AVSS.t111 65.8183
R6377 AVSS.n2670 AVSS.t111 65.8183
R6378 AVSS.n2668 AVSS.t111 65.8183
R6379 AVSS.n1658 AVSS.t113 65.8183
R6380 AVSS.n1652 AVSS.t113 65.8183
R6381 AVSS.n1650 AVSS.t113 65.8183
R6382 AVSS.n1645 AVSS.t113 65.8183
R6383 AVSS.n1665 AVSS.t113 65.8183
R6384 AVSS.n1671 AVSS.t113 65.8183
R6385 AVSS.n1673 AVSS.t113 65.8183
R6386 AVSS.n1694 AVSS.t113 65.8183
R6387 AVSS.n1633 AVSS.t113 65.8183
R6388 AVSS.n1687 AVSS.t113 65.8183
R6389 AVSS.n1681 AVSS.t113 65.8183
R6390 AVSS.n1711 AVSS.t113 65.8183
R6391 AVSS.n1708 AVSS.t113 65.8183
R6392 AVSS.n1702 AVSS.t113 65.8183
R6393 AVSS.n1700 AVSS.t113 65.8183
R6394 AVSS.t77 AVSS.n1984 65.8183
R6395 AVSS.t77 AVSS.n1985 65.8183
R6396 AVSS.t77 AVSS.n1986 65.8183
R6397 AVSS.t77 AVSS.n1987 65.8183
R6398 AVSS.t77 AVSS.n1983 65.8183
R6399 AVSS.t77 AVSS.n1982 65.8183
R6400 AVSS.t77 AVSS.n1981 65.8183
R6401 AVSS.t77 AVSS.n1993 65.8183
R6402 AVSS.t77 AVSS.n1994 65.8183
R6403 AVSS.t77 AVSS.n1995 65.8183
R6404 AVSS.t77 AVSS.n1996 65.8183
R6405 AVSS.t77 AVSS.n1989 65.8183
R6406 AVSS.t77 AVSS.n1990 65.8183
R6407 AVSS.t77 AVSS.n1991 65.8183
R6408 AVSS.t77 AVSS.n2064 65.8183
R6409 AVSS.t87 AVSS.n759 65.8183
R6410 AVSS.t87 AVSS.n758 65.8183
R6411 AVSS.t87 AVSS.n757 65.8183
R6412 AVSS.t87 AVSS.n756 65.8183
R6413 AVSS.t87 AVSS.n749 65.8183
R6414 AVSS.t87 AVSS.n747 65.8183
R6415 AVSS.t87 AVSS.n745 65.8183
R6416 AVSS.n828 AVSS.t87 65.8183
R6417 AVSS.t87 AVSS.n755 65.8183
R6418 AVSS.t87 AVSS.n754 65.8183
R6419 AVSS.t87 AVSS.n753 65.8183
R6420 AVSS.t87 AVSS.n752 65.8183
R6421 AVSS.t87 AVSS.n750 65.8183
R6422 AVSS.t87 AVSS.n748 65.8183
R6423 AVSS.t87 AVSS.n746 65.8183
R6424 AVSS.t87 AVSS.n744 65.8183
R6425 AVSS.t79 AVSS.n1060 65.8183
R6426 AVSS.t79 AVSS.n993 65.8183
R6427 AVSS.t79 AVSS.n992 65.8183
R6428 AVSS.t79 AVSS.n991 65.8183
R6429 AVSS.t79 AVSS.n983 65.8183
R6430 AVSS.t79 AVSS.n981 65.8183
R6431 AVSS.t79 AVSS.n979 65.8183
R6432 AVSS.t79 AVSS.n990 65.8183
R6433 AVSS.t79 AVSS.n989 65.8183
R6434 AVSS.t79 AVSS.n988 65.8183
R6435 AVSS.t79 AVSS.n987 65.8183
R6436 AVSS.t79 AVSS.n986 65.8183
R6437 AVSS.t79 AVSS.n984 65.8183
R6438 AVSS.t79 AVSS.n982 65.8183
R6439 AVSS.t79 AVSS.n980 65.8183
R6440 AVSS.n1061 AVSS.t79 65.8183
R6441 AVSS.n2488 AVSS.t114 65.8183
R6442 AVSS.n2494 AVSS.t114 65.8183
R6443 AVSS.n2496 AVSS.t114 65.8183
R6444 AVSS.n2502 AVSS.t114 65.8183
R6445 AVSS.n2472 AVSS.t114 65.8183
R6446 AVSS.n2478 AVSS.t114 65.8183
R6447 AVSS.n2480 AVSS.t114 65.8183
R6448 AVSS.n2486 AVSS.t114 65.8183
R6449 AVSS.n2456 AVSS.t114 65.8183
R6450 AVSS.n2434 AVSS.t114 65.8183
R6451 AVSS.n2463 AVSS.t114 65.8183
R6452 AVSS.n2431 AVSS.t114 65.8183
R6453 AVSS.n2449 AVSS.t114 65.8183
R6454 AVSS.n2447 AVSS.t114 65.8183
R6455 AVSS.n2441 AVSS.t114 65.8183
R6456 AVSS.n2439 AVSS.t114 65.8183
R6457 AVSS.t81 AVSS.n1894 65.8183
R6458 AVSS.t81 AVSS.n1895 65.8183
R6459 AVSS.t81 AVSS.n1896 65.8183
R6460 AVSS.t81 AVSS.n1897 65.8183
R6461 AVSS.t81 AVSS.n1892 65.8183
R6462 AVSS.t81 AVSS.n1891 65.8183
R6463 AVSS.t81 AVSS.n1890 65.8183
R6464 AVSS.t81 AVSS.n1902 65.8183
R6465 AVSS.t81 AVSS.n1903 65.8183
R6466 AVSS.t81 AVSS.n1904 65.8183
R6467 AVSS.t81 AVSS.n1905 65.8183
R6468 AVSS.t81 AVSS.n1898 65.8183
R6469 AVSS.t81 AVSS.n1899 65.8183
R6470 AVSS.t81 AVSS.n1900 65.8183
R6471 AVSS.t81 AVSS.n1971 65.8183
R6472 AVSS.t82 AVSS.n2556 65.8183
R6473 AVSS.t82 AVSS.n1769 65.8183
R6474 AVSS.t82 AVSS.n1768 65.8183
R6475 AVSS.t82 AVSS.n1767 65.8183
R6476 AVSS.t82 AVSS.n1759 65.8183
R6477 AVSS.t82 AVSS.n1757 65.8183
R6478 AVSS.t82 AVSS.n1755 65.8183
R6479 AVSS.t82 AVSS.n1765 65.8183
R6480 AVSS.t82 AVSS.n1764 65.8183
R6481 AVSS.t82 AVSS.n1763 65.8183
R6482 AVSS.t82 AVSS.n1762 65.8183
R6483 AVSS.t82 AVSS.n1761 65.8183
R6484 AVSS.t82 AVSS.n1760 65.8183
R6485 AVSS.t82 AVSS.n1758 65.8183
R6486 AVSS.t82 AVSS.n1756 65.8183
R6487 AVSS.t82 AVSS.n1754 65.8183
R6488 AVSS.t97 AVSS.n3312 65.8183
R6489 AVSS.t97 AVSS.n3313 65.8183
R6490 AVSS.t97 AVSS.n3314 65.8183
R6491 AVSS.t97 AVSS.n3315 65.8183
R6492 AVSS.t97 AVSS.n3310 65.8183
R6493 AVSS.t97 AVSS.n3309 65.8183
R6494 AVSS.t97 AVSS.n3308 65.8183
R6495 AVSS.t97 AVSS.n3320 65.8183
R6496 AVSS.t97 AVSS.n3321 65.8183
R6497 AVSS.t97 AVSS.n3322 65.8183
R6498 AVSS.t97 AVSS.n3323 65.8183
R6499 AVSS.t97 AVSS.n3316 65.8183
R6500 AVSS.t97 AVSS.n3317 65.8183
R6501 AVSS.t97 AVSS.n3318 65.8183
R6502 AVSS.t97 AVSS.n3390 65.8183
R6503 AVSS.t83 AVSS.n67 64.1729
R6504 AVSS.t105 AVSS.n5737 64.1729
R6505 AVSS.t91 AVSS.n5465 64.1729
R6506 AVSS.n5337 AVSS.t88 64.1729
R6507 AVSS.n5138 AVSS.t98 64.1729
R6508 AVSS.t100 AVSS.n3134 64.1729
R6509 AVSS.t96 AVSS.n1210 64.1729
R6510 AVSS.t112 AVSS.n4534 64.1729
R6511 AVSS.t75 AVSS.n2695 64.1729
R6512 AVSS.t87 AVSS.n751 64.1729
R6513 AVSS.t79 AVSS.n985 64.1729
R6514 AVSS.n2470 AVSS.t114 64.1729
R6515 AVSS.n2557 AVSS.t82 64.1729
R6516 AVSS.t104 AVSS.n305 61.4615
R6517 AVSS.n5964 AVSS.t9 59.1566
R6518 AVSS.n5959 AVSS.n5958 58.5005
R6519 AVSS.n5960 AVSS.n5959 58.5005
R6520 AVSS.n5948 AVSS.n5947 58.5005
R6521 AVSS.n5947 AVSS.n5942 58.5005
R6522 AVSS.t101 AVSS.n4125 57.8461
R6523 AVSS.n4006 AVSS.t94 57.8461
R6524 AVSS.n3795 AVSS.t107 57.8461
R6525 AVSS.n3436 AVSS.t109 57.8461
R6526 AVSS.n548 AVSS.t103 57.8461
R6527 AVSS.t86 AVSS.n1401 57.8461
R6528 AVSS.t93 AVSS.n4821 57.8461
R6529 AVSS.n2608 AVSS.t111 57.8461
R6530 AVSS.n1641 AVSS.t113 57.8461
R6531 AVSS.t77 AVSS.n1988 57.8461
R6532 AVSS.n1972 AVSS.t81 57.8461
R6533 AVSS.n3391 AVSS.t97 57.8461
R6534 AVSS.n99 AVSS.n67 56.6572
R6535 AVSS.n102 AVSS.n67 56.6572
R6536 AVSS.n5780 AVSS.n5737 56.6572
R6537 AVSS.n5777 AVSS.n5737 56.6572
R6538 AVSS.n5508 AVSS.n5465 56.6572
R6539 AVSS.n5505 AVSS.n5465 56.6572
R6540 AVSS.n5338 AVSS.n5337 56.6572
R6541 AVSS.n5337 AVSS.n5336 56.6572
R6542 AVSS.n5139 AVSS.n5138 56.6572
R6543 AVSS.n5138 AVSS.n5137 56.6572
R6544 AVSS.n3173 AVSS.n3134 56.6572
R6545 AVSS.n3176 AVSS.n3134 56.6572
R6546 AVSS.n1249 AVSS.n1210 56.6572
R6547 AVSS.n1252 AVSS.n1210 56.6572
R6548 AVSS.n4577 AVSS.n4534 56.6572
R6549 AVSS.n4574 AVSS.n4534 56.6572
R6550 AVSS.n2727 AVSS.n2695 56.6572
R6551 AVSS.n2730 AVSS.n2695 56.6572
R6552 AVSS.n790 AVSS.n751 56.6572
R6553 AVSS.n793 AVSS.n751 56.6572
R6554 AVSS.n1028 AVSS.n985 56.6572
R6555 AVSS.n1025 AVSS.n985 56.6572
R6556 AVSS.n2471 AVSS.n2470 56.6572
R6557 AVSS.n2470 AVSS.n2469 56.6572
R6558 AVSS.n2558 AVSS.n2557 56.6572
R6559 AVSS.n2557 AVSS.n1753 56.6572
R6560 AVSS.n6034 AVSS.n5940 56.1999
R6561 AVSS.t103 AVSS.n477 55.2026
R6562 AVSS.t86 AVSS.n1405 55.2026
R6563 AVSS.t93 AVSS.n4825 55.2026
R6564 AVSS.t77 AVSS.n1992 55.2026
R6565 AVSS.t81 AVSS.n1901 55.2026
R6566 AVSS.t97 AVSS.n3319 55.2026
R6567 AVSS.t83 AVSS.n72 54.4705
R6568 AVSS.t101 AVSS.n4131 54.4705
R6569 AVSS.n4044 AVSS.t94 54.4705
R6570 AVSS.n3833 AVSS.t107 54.4705
R6571 AVSS.n3474 AVSS.t109 54.4705
R6572 AVSS.t105 AVSS.n5729 54.4705
R6573 AVSS.t91 AVSS.n5457 54.4705
R6574 AVSS.n5371 AVSS.t88 54.4705
R6575 AVSS.n5172 AVSS.t98 54.4705
R6576 AVSS.t100 AVSS.n3210 54.4705
R6577 AVSS.t96 AVSS.n1286 54.4705
R6578 AVSS.t112 AVSS.n4526 54.4705
R6579 AVSS.t75 AVSS.n2700 54.4705
R6580 AVSS.n2646 AVSS.t111 54.4705
R6581 AVSS.n1679 AVSS.t113 54.4705
R6582 AVSS.t87 AVSS.n827 54.4705
R6583 AVSS.t79 AVSS.n977 54.4705
R6584 AVSS.n2505 AVSS.t114 54.4705
R6585 AVSS.t82 AVSS.n1766 54.4705
R6586 AVSS.n144 AVSS.n143 53.3664
R6587 AVSS.n87 AVSS.n71 53.3664
R6588 AVSS.n91 AVSS.n70 53.3664
R6589 AVSS.n95 AVSS.n68 53.3664
R6590 AVSS.n106 AVSS.n63 53.3664
R6591 AVSS.n110 AVSS.n64 53.3664
R6592 AVSS.n114 AVSS.n65 53.3664
R6593 AVSS.n118 AVSS.n66 53.3664
R6594 AVSS.n134 AVSS.n60 53.3664
R6595 AVSS.n130 AVSS.n69 53.3664
R6596 AVSS.n126 AVSS.n61 53.3664
R6597 AVSS.n122 AVSS.n62 53.3664
R6598 AVSS.n79 AVSS.n73 53.3664
R6599 AVSS.n80 AVSS.n74 53.3664
R6600 AVSS.n84 AVSS.n75 53.3664
R6601 AVSS.n142 AVSS.n141 53.3664
R6602 AVSS.n73 AVSS.n58 53.3664
R6603 AVSS.n83 AVSS.n74 53.3664
R6604 AVSS.n77 AVSS.n75 53.3664
R6605 AVSS.n142 AVSS.n76 53.3664
R6606 AVSS.n119 AVSS.n62 53.3664
R6607 AVSS.n123 AVSS.n61 53.3664
R6608 AVSS.n127 AVSS.n69 53.3664
R6609 AVSS.n131 AVSS.n60 53.3664
R6610 AVSS.n115 AVSS.n66 53.3664
R6611 AVSS.n111 AVSS.n65 53.3664
R6612 AVSS.n107 AVSS.n64 53.3664
R6613 AVSS.n103 AVSS.n63 53.3664
R6614 AVSS.n98 AVSS.n68 53.3664
R6615 AVSS.n94 AVSS.n70 53.3664
R6616 AVSS.n90 AVSS.n71 53.3664
R6617 AVSS.n143 AVSS.n59 53.3664
R6618 AVSS.n4154 AVSS.n4126 53.3664
R6619 AVSS.n4158 AVSS.n4127 53.3664
R6620 AVSS.n4162 AVSS.n4128 53.3664
R6621 AVSS.n4166 AVSS.n4129 53.3664
R6622 AVSS.n4163 AVSS.n4129 53.3664
R6623 AVSS.n4159 AVSS.n4128 53.3664
R6624 AVSS.n4155 AVSS.n4127 53.3664
R6625 AVSS.n4151 AVSS.n4126 53.3664
R6626 AVSS.n4183 AVSS.n4119 53.3664
R6627 AVSS.n4179 AVSS.n4130 53.3664
R6628 AVSS.n4175 AVSS.n4122 53.3664
R6629 AVSS.n4172 AVSS.n4122 53.3664
R6630 AVSS.n4176 AVSS.n4130 53.3664
R6631 AVSS.n4180 AVSS.n4119 53.3664
R6632 AVSS.n4201 AVSS.n4116 53.3664
R6633 AVSS.n4135 AVSS.n4134 53.3664
R6634 AVSS.n4195 AVSS.n4133 53.3664
R6635 AVSS.n4191 AVSS.n4132 53.3664
R6636 AVSS.n4201 AVSS.n4200 53.3664
R6637 AVSS.n4196 AVSS.n4134 53.3664
R6638 AVSS.n4192 AVSS.n4133 53.3664
R6639 AVSS.n4188 AVSS.n4132 53.3664
R6640 AVSS.n4118 AVSS.n4117 53.3664
R6641 AVSS.n4139 AVSS.n4120 53.3664
R6642 AVSS.n4143 AVSS.n4121 53.3664
R6643 AVSS.n4147 AVSS.n4123 53.3664
R6644 AVSS.n4150 AVSS.n4123 53.3664
R6645 AVSS.n4146 AVSS.n4121 53.3664
R6646 AVSS.n4142 AVSS.n4120 53.3664
R6647 AVSS.n4138 AVSS.n4118 53.3664
R6648 AVSS.n4011 AVSS.n4010 53.3664
R6649 AVSS.n4016 AVSS.n4015 53.3664
R6650 AVSS.n4017 AVSS.n4008 53.3664
R6651 AVSS.n4024 AVSS.n4023 53.3664
R6652 AVSS.n4023 AVSS.n4022 53.3664
R6653 AVSS.n4018 AVSS.n4017 53.3664
R6654 AVSS.n4015 AVSS.n4014 53.3664
R6655 AVSS.n4010 AVSS.n3992 53.3664
R6656 AVSS.n4038 AVSS.n4002 53.3664
R6657 AVSS.n4037 AVSS.n4036 53.3664
R6658 AVSS.n4030 AVSS.n4004 53.3664
R6659 AVSS.n4031 AVSS.n4030 53.3664
R6660 AVSS.n4036 AVSS.n4035 53.3664
R6661 AVSS.n4039 AVSS.n4038 53.3664
R6662 AVSS.n4060 AVSS.n4059 53.3664
R6663 AVSS.n4057 AVSS.n3998 53.3664
R6664 AVSS.n4053 AVSS.n4052 53.3664
R6665 AVSS.n4046 AVSS.n4000 53.3664
R6666 AVSS.n4059 AVSS.n4058 53.3664
R6667 AVSS.n4054 AVSS.n3998 53.3664
R6668 AVSS.n4052 AVSS.n4051 53.3664
R6669 AVSS.n4047 AVSS.n4046 53.3664
R6670 AVSS.n4066 AVSS.n4065 53.3664
R6671 AVSS.n4069 AVSS.n4068 53.3664
R6672 AVSS.n4074 AVSS.n4073 53.3664
R6673 AVSS.n4077 AVSS.n4076 53.3664
R6674 AVSS.n4078 AVSS.n4077 53.3664
R6675 AVSS.n4075 AVSS.n4074 53.3664
R6676 AVSS.n4068 AVSS.n3994 53.3664
R6677 AVSS.n4067 AVSS.n4066 53.3664
R6678 AVSS.n3800 AVSS.n3799 53.3664
R6679 AVSS.n3805 AVSS.n3804 53.3664
R6680 AVSS.n3806 AVSS.n3797 53.3664
R6681 AVSS.n3813 AVSS.n3812 53.3664
R6682 AVSS.n3812 AVSS.n3811 53.3664
R6683 AVSS.n3807 AVSS.n3806 53.3664
R6684 AVSS.n3804 AVSS.n3803 53.3664
R6685 AVSS.n3799 AVSS.n3781 53.3664
R6686 AVSS.n3827 AVSS.n3791 53.3664
R6687 AVSS.n3826 AVSS.n3825 53.3664
R6688 AVSS.n3819 AVSS.n3793 53.3664
R6689 AVSS.n3820 AVSS.n3819 53.3664
R6690 AVSS.n3825 AVSS.n3824 53.3664
R6691 AVSS.n3828 AVSS.n3827 53.3664
R6692 AVSS.n3849 AVSS.n3848 53.3664
R6693 AVSS.n3846 AVSS.n3787 53.3664
R6694 AVSS.n3842 AVSS.n3841 53.3664
R6695 AVSS.n3835 AVSS.n3789 53.3664
R6696 AVSS.n3848 AVSS.n3847 53.3664
R6697 AVSS.n3843 AVSS.n3787 53.3664
R6698 AVSS.n3841 AVSS.n3840 53.3664
R6699 AVSS.n3836 AVSS.n3835 53.3664
R6700 AVSS.n3855 AVSS.n3854 53.3664
R6701 AVSS.n3858 AVSS.n3857 53.3664
R6702 AVSS.n3863 AVSS.n3862 53.3664
R6703 AVSS.n3866 AVSS.n3865 53.3664
R6704 AVSS.n3867 AVSS.n3866 53.3664
R6705 AVSS.n3864 AVSS.n3863 53.3664
R6706 AVSS.n3857 AVSS.n3783 53.3664
R6707 AVSS.n3856 AVSS.n3855 53.3664
R6708 AVSS.n3495 AVSS.n3494 53.3664
R6709 AVSS.n3498 AVSS.n3497 53.3664
R6710 AVSS.n3503 AVSS.n3502 53.3664
R6711 AVSS.n3506 AVSS.n3505 53.3664
R6712 AVSS.n3490 AVSS.n3489 53.3664
R6713 AVSS.n3487 AVSS.n3428 53.3664
R6714 AVSS.n3483 AVSS.n3482 53.3664
R6715 AVSS.n3476 AVSS.n3430 53.3664
R6716 AVSS.n3468 AVSS.n3432 53.3664
R6717 AVSS.n3467 AVSS.n3466 53.3664
R6718 AVSS.n3460 AVSS.n3434 53.3664
R6719 AVSS.n3441 AVSS.n3440 53.3664
R6720 AVSS.n3446 AVSS.n3445 53.3664
R6721 AVSS.n3447 AVSS.n3438 53.3664
R6722 AVSS.n3454 AVSS.n3453 53.3664
R6723 AVSS.n3453 AVSS.n3452 53.3664
R6724 AVSS.n3448 AVSS.n3447 53.3664
R6725 AVSS.n3445 AVSS.n3444 53.3664
R6726 AVSS.n3440 AVSS.n3422 53.3664
R6727 AVSS.n3461 AVSS.n3460 53.3664
R6728 AVSS.n3466 AVSS.n3465 53.3664
R6729 AVSS.n3469 AVSS.n3468 53.3664
R6730 AVSS.n3489 AVSS.n3488 53.3664
R6731 AVSS.n3484 AVSS.n3428 53.3664
R6732 AVSS.n3482 AVSS.n3481 53.3664
R6733 AVSS.n3477 AVSS.n3476 53.3664
R6734 AVSS.n3507 AVSS.n3506 53.3664
R6735 AVSS.n3504 AVSS.n3503 53.3664
R6736 AVSS.n3497 AVSS.n3424 53.3664
R6737 AVSS.n3496 AVSS.n3495 53.3664
R6738 AVSS.n5795 AVSS.n5742 53.3664
R6739 AVSS.n5792 AVSS.n5731 53.3664
R6740 AVSS.n5788 AVSS.n5733 53.3664
R6741 AVSS.n5784 AVSS.n5735 53.3664
R6742 AVSS.n5773 AVSS.n5738 53.3664
R6743 AVSS.n5769 AVSS.n5739 53.3664
R6744 AVSS.n5765 AVSS.n5740 53.3664
R6745 AVSS.n5761 AVSS.n5741 53.3664
R6746 AVSS.n5814 AVSS.n5813 53.3664
R6747 AVSS.n5749 AVSS.n5732 53.3664
R6748 AVSS.n5753 AVSS.n5734 53.3664
R6749 AVSS.n5757 AVSS.n5736 53.3664
R6750 AVSS.n5812 AVSS.n5811 53.3664
R6751 AVSS.n5747 AVSS.n5745 53.3664
R6752 AVSS.n5806 AVSS.n5744 53.3664
R6753 AVSS.n5802 AVSS.n5743 53.3664
R6754 AVSS.n5812 AVSS.n5746 53.3664
R6755 AVSS.n5807 AVSS.n5745 53.3664
R6756 AVSS.n5803 AVSS.n5744 53.3664
R6757 AVSS.n5799 AVSS.n5743 53.3664
R6758 AVSS.n5781 AVSS.n5735 53.3664
R6759 AVSS.n5785 AVSS.n5733 53.3664
R6760 AVSS.n5789 AVSS.n5731 53.3664
R6761 AVSS.n5793 AVSS.n5742 53.3664
R6762 AVSS.n5764 AVSS.n5741 53.3664
R6763 AVSS.n5768 AVSS.n5740 53.3664
R6764 AVSS.n5772 AVSS.n5739 53.3664
R6765 AVSS.n5776 AVSS.n5738 53.3664
R6766 AVSS.n5760 AVSS.n5736 53.3664
R6767 AVSS.n5756 AVSS.n5734 53.3664
R6768 AVSS.n5752 AVSS.n5732 53.3664
R6769 AVSS.n5813 AVSS.n5730 53.3664
R6770 AVSS.n5523 AVSS.n5470 53.3664
R6771 AVSS.n5520 AVSS.n5459 53.3664
R6772 AVSS.n5516 AVSS.n5461 53.3664
R6773 AVSS.n5512 AVSS.n5463 53.3664
R6774 AVSS.n5501 AVSS.n5466 53.3664
R6775 AVSS.n5497 AVSS.n5467 53.3664
R6776 AVSS.n5493 AVSS.n5468 53.3664
R6777 AVSS.n5489 AVSS.n5469 53.3664
R6778 AVSS.n5542 AVSS.n5541 53.3664
R6779 AVSS.n5477 AVSS.n5460 53.3664
R6780 AVSS.n5481 AVSS.n5462 53.3664
R6781 AVSS.n5485 AVSS.n5464 53.3664
R6782 AVSS.n5540 AVSS.n5539 53.3664
R6783 AVSS.n5475 AVSS.n5473 53.3664
R6784 AVSS.n5534 AVSS.n5472 53.3664
R6785 AVSS.n5530 AVSS.n5471 53.3664
R6786 AVSS.n5540 AVSS.n5474 53.3664
R6787 AVSS.n5535 AVSS.n5473 53.3664
R6788 AVSS.n5531 AVSS.n5472 53.3664
R6789 AVSS.n5527 AVSS.n5471 53.3664
R6790 AVSS.n5509 AVSS.n5463 53.3664
R6791 AVSS.n5513 AVSS.n5461 53.3664
R6792 AVSS.n5517 AVSS.n5459 53.3664
R6793 AVSS.n5521 AVSS.n5470 53.3664
R6794 AVSS.n5492 AVSS.n5469 53.3664
R6795 AVSS.n5496 AVSS.n5468 53.3664
R6796 AVSS.n5500 AVSS.n5467 53.3664
R6797 AVSS.n5504 AVSS.n5466 53.3664
R6798 AVSS.n5488 AVSS.n5464 53.3664
R6799 AVSS.n5484 AVSS.n5462 53.3664
R6800 AVSS.n5480 AVSS.n5460 53.3664
R6801 AVSS.n5541 AVSS.n5458 53.3664
R6802 AVSS.n5355 AVSS.n5311 53.3664
R6803 AVSS.n5361 AVSS.n5360 53.3664
R6804 AVSS.n5364 AVSS.n5363 53.3664
R6805 AVSS.n5369 AVSS.n5368 53.3664
R6806 AVSS.n5356 AVSS.n5355 53.3664
R6807 AVSS.n5362 AVSS.n5361 53.3664
R6808 AVSS.n5363 AVSS.n5309 53.3664
R6809 AVSS.n5370 AVSS.n5369 53.3664
R6810 AVSS.n5354 AVSS.n5353 53.3664
R6811 AVSS.n5347 AVSS.n5313 53.3664
R6812 AVSS.n5346 AVSS.n5345 53.3664
R6813 AVSS.n5339 AVSS.n5315 53.3664
R6814 AVSS.n5340 AVSS.n5339 53.3664
R6815 AVSS.n5345 AVSS.n5344 53.3664
R6816 AVSS.n5348 AVSS.n5347 53.3664
R6817 AVSS.n5353 AVSS.n5352 53.3664
R6818 AVSS.n5332 AVSS.n5319 53.3664
R6819 AVSS.n5330 AVSS.n5329 53.3664
R6820 AVSS.n5325 AVSS.n5322 53.3664
R6821 AVSS.n5323 AVSS.n5303 53.3664
R6822 AVSS.n5324 AVSS.n5323 53.3664
R6823 AVSS.n5322 AVSS.n5320 53.3664
R6824 AVSS.n5331 AVSS.n5330 53.3664
R6825 AVSS.n5319 AVSS.n5317 53.3664
R6826 AVSS.n5378 AVSS.n5377 53.3664
R6827 AVSS.n5381 AVSS.n5380 53.3664
R6828 AVSS.n5386 AVSS.n5385 53.3664
R6829 AVSS.n5389 AVSS.n5388 53.3664
R6830 AVSS.n5390 AVSS.n5389 53.3664
R6831 AVSS.n5387 AVSS.n5386 53.3664
R6832 AVSS.n5380 AVSS.n5305 53.3664
R6833 AVSS.n5379 AVSS.n5378 53.3664
R6834 AVSS.n5156 AVSS.n5112 53.3664
R6835 AVSS.n5162 AVSS.n5161 53.3664
R6836 AVSS.n5165 AVSS.n5164 53.3664
R6837 AVSS.n5170 AVSS.n5169 53.3664
R6838 AVSS.n5157 AVSS.n5156 53.3664
R6839 AVSS.n5163 AVSS.n5162 53.3664
R6840 AVSS.n5164 AVSS.n5110 53.3664
R6841 AVSS.n5171 AVSS.n5170 53.3664
R6842 AVSS.n5155 AVSS.n5154 53.3664
R6843 AVSS.n5148 AVSS.n5114 53.3664
R6844 AVSS.n5147 AVSS.n5146 53.3664
R6845 AVSS.n5140 AVSS.n5116 53.3664
R6846 AVSS.n5141 AVSS.n5140 53.3664
R6847 AVSS.n5146 AVSS.n5145 53.3664
R6848 AVSS.n5149 AVSS.n5148 53.3664
R6849 AVSS.n5154 AVSS.n5153 53.3664
R6850 AVSS.n5133 AVSS.n5120 53.3664
R6851 AVSS.n5131 AVSS.n5130 53.3664
R6852 AVSS.n5126 AVSS.n5123 53.3664
R6853 AVSS.n5124 AVSS.n5104 53.3664
R6854 AVSS.n5125 AVSS.n5124 53.3664
R6855 AVSS.n5123 AVSS.n5121 53.3664
R6856 AVSS.n5132 AVSS.n5131 53.3664
R6857 AVSS.n5120 AVSS.n5118 53.3664
R6858 AVSS.n5179 AVSS.n5178 53.3664
R6859 AVSS.n5182 AVSS.n5181 53.3664
R6860 AVSS.n5187 AVSS.n5186 53.3664
R6861 AVSS.n5190 AVSS.n5189 53.3664
R6862 AVSS.n5191 AVSS.n5190 53.3664
R6863 AVSS.n5188 AVSS.n5187 53.3664
R6864 AVSS.n5181 AVSS.n5106 53.3664
R6865 AVSS.n5180 AVSS.n5179 53.3664
R6866 AVSS.n512 AVSS.n466 53.3664
R6867 AVSS.n509 AVSS.n467 53.3664
R6868 AVSS.n505 AVSS.n468 53.3664
R6869 AVSS.n519 AVSS.n478 53.3664
R6870 AVSS.n523 AVSS.n479 53.3664
R6871 AVSS.n527 AVSS.n480 53.3664
R6872 AVSS.n531 AVSS.n481 53.3664
R6873 AVSS.n547 AVSS.n546 53.3664
R6874 AVSS.n542 AVSS.n476 53.3664
R6875 AVSS.n539 AVSS.n475 53.3664
R6876 AVSS.n535 AVSS.n474 53.3664
R6877 AVSS.n497 AVSS.n473 53.3664
R6878 AVSS.n493 AVSS.n472 53.3664
R6879 AVSS.n489 AVSS.n471 53.3664
R6880 AVSS.n485 AVSS.n470 53.3664
R6881 AVSS.n488 AVSS.n470 53.3664
R6882 AVSS.n492 AVSS.n471 53.3664
R6883 AVSS.n496 AVSS.n472 53.3664
R6884 AVSS.n499 AVSS.n473 53.3664
R6885 AVSS.n502 AVSS.n468 53.3664
R6886 AVSS.n506 AVSS.n467 53.3664
R6887 AVSS.n510 AVSS.n466 53.3664
R6888 AVSS.n522 AVSS.n478 53.3664
R6889 AVSS.n526 AVSS.n479 53.3664
R6890 AVSS.n530 AVSS.n480 53.3664
R6891 AVSS.n484 AVSS.n481 53.3664
R6892 AVSS.n474 AVSS.n464 53.3664
R6893 AVSS.n536 AVSS.n475 53.3664
R6894 AVSS.n540 AVSS.n476 53.3664
R6895 AVSS.n547 AVSS.n483 53.3664
R6896 AVSS.n1444 AVSS.n1400 53.3664
R6897 AVSS.n1448 AVSS.n1399 53.3664
R6898 AVSS.n1452 AVSS.n1398 53.3664
R6899 AVSS.n1456 AVSS.n1397 53.3664
R6900 AVSS.n1453 AVSS.n1397 53.3664
R6901 AVSS.n1449 AVSS.n1398 53.3664
R6902 AVSS.n1445 AVSS.n1399 53.3664
R6903 AVSS.n1400 AVSS.n1393 53.3664
R6904 AVSS.n1477 AVSS.n1476 53.3664
R6905 AVSS.n1472 AVSS.n1404 53.3664
R6906 AVSS.n1469 AVSS.n1403 53.3664
R6907 AVSS.n1465 AVSS.n1402 53.3664
R6908 AVSS.n1428 AVSS.n1406 53.3664
R6909 AVSS.n1432 AVSS.n1407 53.3664
R6910 AVSS.n1436 AVSS.n1408 53.3664
R6911 AVSS.n1440 AVSS.n1409 53.3664
R6912 AVSS.n1421 AVSS.n1394 53.3664
R6913 AVSS.n1418 AVSS.n1395 53.3664
R6914 AVSS.n1414 AVSS.n1396 53.3664
R6915 AVSS.n1396 AVSS.n1392 53.3664
R6916 AVSS.n1415 AVSS.n1395 53.3664
R6917 AVSS.n1419 AVSS.n1394 53.3664
R6918 AVSS.n1431 AVSS.n1406 53.3664
R6919 AVSS.n1435 AVSS.n1407 53.3664
R6920 AVSS.n1439 AVSS.n1408 53.3664
R6921 AVSS.n1412 AVSS.n1409 53.3664
R6922 AVSS.n1462 AVSS.n1402 53.3664
R6923 AVSS.n1466 AVSS.n1403 53.3664
R6924 AVSS.n1470 AVSS.n1404 53.3664
R6925 AVSS.n1477 AVSS.n1411 53.3664
R6926 AVSS.n4864 AVSS.n4820 53.3664
R6927 AVSS.n4868 AVSS.n4819 53.3664
R6928 AVSS.n4872 AVSS.n4818 53.3664
R6929 AVSS.n4876 AVSS.n4817 53.3664
R6930 AVSS.n4873 AVSS.n4817 53.3664
R6931 AVSS.n4869 AVSS.n4818 53.3664
R6932 AVSS.n4865 AVSS.n4819 53.3664
R6933 AVSS.n4820 AVSS.n4813 53.3664
R6934 AVSS.n4897 AVSS.n4896 53.3664
R6935 AVSS.n4892 AVSS.n4824 53.3664
R6936 AVSS.n4889 AVSS.n4823 53.3664
R6937 AVSS.n4885 AVSS.n4822 53.3664
R6938 AVSS.n4848 AVSS.n4826 53.3664
R6939 AVSS.n4852 AVSS.n4827 53.3664
R6940 AVSS.n4856 AVSS.n4828 53.3664
R6941 AVSS.n4860 AVSS.n4829 53.3664
R6942 AVSS.n4841 AVSS.n4814 53.3664
R6943 AVSS.n4838 AVSS.n4815 53.3664
R6944 AVSS.n4834 AVSS.n4816 53.3664
R6945 AVSS.n4816 AVSS.n4812 53.3664
R6946 AVSS.n4835 AVSS.n4815 53.3664
R6947 AVSS.n4839 AVSS.n4814 53.3664
R6948 AVSS.n4851 AVSS.n4826 53.3664
R6949 AVSS.n4855 AVSS.n4827 53.3664
R6950 AVSS.n4859 AVSS.n4828 53.3664
R6951 AVSS.n4832 AVSS.n4829 53.3664
R6952 AVSS.n4882 AVSS.n4822 53.3664
R6953 AVSS.n4886 AVSS.n4823 53.3664
R6954 AVSS.n4890 AVSS.n4824 53.3664
R6955 AVSS.n4897 AVSS.n4831 53.3664
R6956 AVSS.n3180 AVSS.n3135 53.3664
R6957 AVSS.n3184 AVSS.n3136 53.3664
R6958 AVSS.n3188 AVSS.n3137 53.3664
R6959 AVSS.n3192 AVSS.n3138 53.3664
R6960 AVSS.n3144 AVSS.n3127 53.3664
R6961 AVSS.n3204 AVSS.n3129 53.3664
R6962 AVSS.n3200 AVSS.n3131 53.3664
R6963 AVSS.n3196 AVSS.n3133 53.3664
R6964 AVSS.n3146 AVSS.n3142 53.3664
R6965 AVSS.n3147 AVSS.n3141 53.3664
R6966 AVSS.n3151 AVSS.n3140 53.3664
R6967 AVSS.n3155 AVSS.n3139 53.3664
R6968 AVSS.n3142 AVSS.n3125 53.3664
R6969 AVSS.n3150 AVSS.n3141 53.3664
R6970 AVSS.n3154 AVSS.n3140 53.3664
R6971 AVSS.n3157 AVSS.n3139 53.3664
R6972 AVSS.n3212 AVSS.n3211 53.3664
R6973 AVSS.n3161 AVSS.n3128 53.3664
R6974 AVSS.n3165 AVSS.n3130 53.3664
R6975 AVSS.n3169 AVSS.n3132 53.3664
R6976 AVSS.n3172 AVSS.n3132 53.3664
R6977 AVSS.n3168 AVSS.n3130 53.3664
R6978 AVSS.n3164 AVSS.n3128 53.3664
R6979 AVSS.n3211 AVSS.n3126 53.3664
R6980 AVSS.n3189 AVSS.n3138 53.3664
R6981 AVSS.n3185 AVSS.n3137 53.3664
R6982 AVSS.n3181 AVSS.n3136 53.3664
R6983 AVSS.n3177 AVSS.n3135 53.3664
R6984 AVSS.n3193 AVSS.n3133 53.3664
R6985 AVSS.n3197 AVSS.n3131 53.3664
R6986 AVSS.n3201 AVSS.n3129 53.3664
R6987 AVSS.n3205 AVSS.n3127 53.3664
R6988 AVSS.n1256 AVSS.n1211 53.3664
R6989 AVSS.n1260 AVSS.n1212 53.3664
R6990 AVSS.n1264 AVSS.n1213 53.3664
R6991 AVSS.n1268 AVSS.n1214 53.3664
R6992 AVSS.n1220 AVSS.n1203 53.3664
R6993 AVSS.n1280 AVSS.n1205 53.3664
R6994 AVSS.n1276 AVSS.n1207 53.3664
R6995 AVSS.n1272 AVSS.n1209 53.3664
R6996 AVSS.n1222 AVSS.n1218 53.3664
R6997 AVSS.n1223 AVSS.n1217 53.3664
R6998 AVSS.n1227 AVSS.n1216 53.3664
R6999 AVSS.n1231 AVSS.n1215 53.3664
R7000 AVSS.n1218 AVSS.n1201 53.3664
R7001 AVSS.n1226 AVSS.n1217 53.3664
R7002 AVSS.n1230 AVSS.n1216 53.3664
R7003 AVSS.n1233 AVSS.n1215 53.3664
R7004 AVSS.n1288 AVSS.n1287 53.3664
R7005 AVSS.n1237 AVSS.n1204 53.3664
R7006 AVSS.n1241 AVSS.n1206 53.3664
R7007 AVSS.n1245 AVSS.n1208 53.3664
R7008 AVSS.n1248 AVSS.n1208 53.3664
R7009 AVSS.n1244 AVSS.n1206 53.3664
R7010 AVSS.n1240 AVSS.n1204 53.3664
R7011 AVSS.n1287 AVSS.n1202 53.3664
R7012 AVSS.n1265 AVSS.n1214 53.3664
R7013 AVSS.n1261 AVSS.n1213 53.3664
R7014 AVSS.n1257 AVSS.n1212 53.3664
R7015 AVSS.n1253 AVSS.n1211 53.3664
R7016 AVSS.n1269 AVSS.n1209 53.3664
R7017 AVSS.n1273 AVSS.n1207 53.3664
R7018 AVSS.n1277 AVSS.n1205 53.3664
R7019 AVSS.n1281 AVSS.n1203 53.3664
R7020 AVSS.n4570 AVSS.n4535 53.3664
R7021 AVSS.n4566 AVSS.n4536 53.3664
R7022 AVSS.n4562 AVSS.n4537 53.3664
R7023 AVSS.n4558 AVSS.n4538 53.3664
R7024 AVSS.n4612 AVSS.n4611 53.3664
R7025 AVSS.n4546 AVSS.n4529 53.3664
R7026 AVSS.n4550 AVSS.n4531 53.3664
R7027 AVSS.n4554 AVSS.n4533 53.3664
R7028 AVSS.n4610 AVSS.n4609 53.3664
R7029 AVSS.n4544 AVSS.n4542 53.3664
R7030 AVSS.n4604 AVSS.n4541 53.3664
R7031 AVSS.n4600 AVSS.n4540 53.3664
R7032 AVSS.n4610 AVSS.n4543 53.3664
R7033 AVSS.n4605 AVSS.n4542 53.3664
R7034 AVSS.n4601 AVSS.n4541 53.3664
R7035 AVSS.n4597 AVSS.n4540 53.3664
R7036 AVSS.n4592 AVSS.n4539 53.3664
R7037 AVSS.n4589 AVSS.n4528 53.3664
R7038 AVSS.n4585 AVSS.n4530 53.3664
R7039 AVSS.n4581 AVSS.n4532 53.3664
R7040 AVSS.n4578 AVSS.n4532 53.3664
R7041 AVSS.n4582 AVSS.n4530 53.3664
R7042 AVSS.n4586 AVSS.n4528 53.3664
R7043 AVSS.n4590 AVSS.n4539 53.3664
R7044 AVSS.n4561 AVSS.n4538 53.3664
R7045 AVSS.n4565 AVSS.n4537 53.3664
R7046 AVSS.n4569 AVSS.n4536 53.3664
R7047 AVSS.n4573 AVSS.n4535 53.3664
R7048 AVSS.n4557 AVSS.n4533 53.3664
R7049 AVSS.n4553 AVSS.n4531 53.3664
R7050 AVSS.n4549 AVSS.n4529 53.3664
R7051 AVSS.n4611 AVSS.n4527 53.3664
R7052 AVSS.n2772 AVSS.n2771 53.3664
R7053 AVSS.n2715 AVSS.n2699 53.3664
R7054 AVSS.n2719 AVSS.n2698 53.3664
R7055 AVSS.n2723 AVSS.n2696 53.3664
R7056 AVSS.n2734 AVSS.n2691 53.3664
R7057 AVSS.n2738 AVSS.n2692 53.3664
R7058 AVSS.n2742 AVSS.n2693 53.3664
R7059 AVSS.n2746 AVSS.n2694 53.3664
R7060 AVSS.n2762 AVSS.n2688 53.3664
R7061 AVSS.n2758 AVSS.n2697 53.3664
R7062 AVSS.n2754 AVSS.n2689 53.3664
R7063 AVSS.n2750 AVSS.n2690 53.3664
R7064 AVSS.n2707 AVSS.n2701 53.3664
R7065 AVSS.n2708 AVSS.n2702 53.3664
R7066 AVSS.n2712 AVSS.n2703 53.3664
R7067 AVSS.n2770 AVSS.n2769 53.3664
R7068 AVSS.n2701 AVSS.n2686 53.3664
R7069 AVSS.n2711 AVSS.n2702 53.3664
R7070 AVSS.n2705 AVSS.n2703 53.3664
R7071 AVSS.n2770 AVSS.n2704 53.3664
R7072 AVSS.n2747 AVSS.n2690 53.3664
R7073 AVSS.n2751 AVSS.n2689 53.3664
R7074 AVSS.n2755 AVSS.n2697 53.3664
R7075 AVSS.n2759 AVSS.n2688 53.3664
R7076 AVSS.n2743 AVSS.n2694 53.3664
R7077 AVSS.n2739 AVSS.n2693 53.3664
R7078 AVSS.n2735 AVSS.n2692 53.3664
R7079 AVSS.n2731 AVSS.n2691 53.3664
R7080 AVSS.n2726 AVSS.n2696 53.3664
R7081 AVSS.n2722 AVSS.n2698 53.3664
R7082 AVSS.n2718 AVSS.n2699 53.3664
R7083 AVSS.n2771 AVSS.n2687 53.3664
R7084 AVSS.n2613 AVSS.n2612 53.3664
R7085 AVSS.n2618 AVSS.n2617 53.3664
R7086 AVSS.n2619 AVSS.n2610 53.3664
R7087 AVSS.n2626 AVSS.n2625 53.3664
R7088 AVSS.n2625 AVSS.n2624 53.3664
R7089 AVSS.n2620 AVSS.n2619 53.3664
R7090 AVSS.n2617 AVSS.n2616 53.3664
R7091 AVSS.n2612 AVSS.n2594 53.3664
R7092 AVSS.n2640 AVSS.n2604 53.3664
R7093 AVSS.n2639 AVSS.n2638 53.3664
R7094 AVSS.n2632 AVSS.n2606 53.3664
R7095 AVSS.n2633 AVSS.n2632 53.3664
R7096 AVSS.n2638 AVSS.n2637 53.3664
R7097 AVSS.n2641 AVSS.n2640 53.3664
R7098 AVSS.n2662 AVSS.n2661 53.3664
R7099 AVSS.n2659 AVSS.n2600 53.3664
R7100 AVSS.n2655 AVSS.n2654 53.3664
R7101 AVSS.n2648 AVSS.n2602 53.3664
R7102 AVSS.n2661 AVSS.n2660 53.3664
R7103 AVSS.n2656 AVSS.n2600 53.3664
R7104 AVSS.n2654 AVSS.n2653 53.3664
R7105 AVSS.n2649 AVSS.n2648 53.3664
R7106 AVSS.n2668 AVSS.n2667 53.3664
R7107 AVSS.n2671 AVSS.n2670 53.3664
R7108 AVSS.n2676 AVSS.n2675 53.3664
R7109 AVSS.n2679 AVSS.n2678 53.3664
R7110 AVSS.n2680 AVSS.n2679 53.3664
R7111 AVSS.n2677 AVSS.n2676 53.3664
R7112 AVSS.n2670 AVSS.n2596 53.3664
R7113 AVSS.n2669 AVSS.n2668 53.3664
R7114 AVSS.n1700 AVSS.n1699 53.3664
R7115 AVSS.n1703 AVSS.n1702 53.3664
R7116 AVSS.n1708 AVSS.n1707 53.3664
R7117 AVSS.n1711 AVSS.n1710 53.3664
R7118 AVSS.n1695 AVSS.n1694 53.3664
R7119 AVSS.n1692 AVSS.n1633 53.3664
R7120 AVSS.n1688 AVSS.n1687 53.3664
R7121 AVSS.n1681 AVSS.n1635 53.3664
R7122 AVSS.n1673 AVSS.n1637 53.3664
R7123 AVSS.n1672 AVSS.n1671 53.3664
R7124 AVSS.n1665 AVSS.n1639 53.3664
R7125 AVSS.n1646 AVSS.n1645 53.3664
R7126 AVSS.n1651 AVSS.n1650 53.3664
R7127 AVSS.n1652 AVSS.n1643 53.3664
R7128 AVSS.n1659 AVSS.n1658 53.3664
R7129 AVSS.n1658 AVSS.n1657 53.3664
R7130 AVSS.n1653 AVSS.n1652 53.3664
R7131 AVSS.n1650 AVSS.n1649 53.3664
R7132 AVSS.n1645 AVSS.n1627 53.3664
R7133 AVSS.n1666 AVSS.n1665 53.3664
R7134 AVSS.n1671 AVSS.n1670 53.3664
R7135 AVSS.n1674 AVSS.n1673 53.3664
R7136 AVSS.n1694 AVSS.n1693 53.3664
R7137 AVSS.n1689 AVSS.n1633 53.3664
R7138 AVSS.n1687 AVSS.n1686 53.3664
R7139 AVSS.n1682 AVSS.n1681 53.3664
R7140 AVSS.n1712 AVSS.n1711 53.3664
R7141 AVSS.n1709 AVSS.n1708 53.3664
R7142 AVSS.n1702 AVSS.n1629 53.3664
R7143 AVSS.n1701 AVSS.n1700 53.3664
R7144 AVSS.n2031 AVSS.n1987 53.3664
R7145 AVSS.n2035 AVSS.n1986 53.3664
R7146 AVSS.n2039 AVSS.n1985 53.3664
R7147 AVSS.n2043 AVSS.n1984 53.3664
R7148 AVSS.n2040 AVSS.n1984 53.3664
R7149 AVSS.n2036 AVSS.n1985 53.3664
R7150 AVSS.n2032 AVSS.n1986 53.3664
R7151 AVSS.n1987 AVSS.n1980 53.3664
R7152 AVSS.n2064 AVSS.n2063 53.3664
R7153 AVSS.n2059 AVSS.n1991 53.3664
R7154 AVSS.n2056 AVSS.n1990 53.3664
R7155 AVSS.n2052 AVSS.n1989 53.3664
R7156 AVSS.n2015 AVSS.n1993 53.3664
R7157 AVSS.n2019 AVSS.n1994 53.3664
R7158 AVSS.n2023 AVSS.n1995 53.3664
R7159 AVSS.n2027 AVSS.n1996 53.3664
R7160 AVSS.n2008 AVSS.n1981 53.3664
R7161 AVSS.n2005 AVSS.n1982 53.3664
R7162 AVSS.n2001 AVSS.n1983 53.3664
R7163 AVSS.n1983 AVSS.n1979 53.3664
R7164 AVSS.n2002 AVSS.n1982 53.3664
R7165 AVSS.n2006 AVSS.n1981 53.3664
R7166 AVSS.n2018 AVSS.n1993 53.3664
R7167 AVSS.n2022 AVSS.n1994 53.3664
R7168 AVSS.n2026 AVSS.n1995 53.3664
R7169 AVSS.n1999 AVSS.n1996 53.3664
R7170 AVSS.n2049 AVSS.n1989 53.3664
R7171 AVSS.n2053 AVSS.n1990 53.3664
R7172 AVSS.n2057 AVSS.n1991 53.3664
R7173 AVSS.n2064 AVSS.n1998 53.3664
R7174 AVSS.n797 AVSS.n752 53.3664
R7175 AVSS.n801 AVSS.n753 53.3664
R7176 AVSS.n805 AVSS.n754 53.3664
R7177 AVSS.n809 AVSS.n755 53.3664
R7178 AVSS.n761 AVSS.n744 53.3664
R7179 AVSS.n821 AVSS.n746 53.3664
R7180 AVSS.n817 AVSS.n748 53.3664
R7181 AVSS.n813 AVSS.n750 53.3664
R7182 AVSS.n763 AVSS.n759 53.3664
R7183 AVSS.n764 AVSS.n758 53.3664
R7184 AVSS.n768 AVSS.n757 53.3664
R7185 AVSS.n772 AVSS.n756 53.3664
R7186 AVSS.n759 AVSS.n742 53.3664
R7187 AVSS.n767 AVSS.n758 53.3664
R7188 AVSS.n771 AVSS.n757 53.3664
R7189 AVSS.n774 AVSS.n756 53.3664
R7190 AVSS.n829 AVSS.n828 53.3664
R7191 AVSS.n778 AVSS.n745 53.3664
R7192 AVSS.n782 AVSS.n747 53.3664
R7193 AVSS.n786 AVSS.n749 53.3664
R7194 AVSS.n789 AVSS.n749 53.3664
R7195 AVSS.n785 AVSS.n747 53.3664
R7196 AVSS.n781 AVSS.n745 53.3664
R7197 AVSS.n828 AVSS.n743 53.3664
R7198 AVSS.n806 AVSS.n755 53.3664
R7199 AVSS.n802 AVSS.n754 53.3664
R7200 AVSS.n798 AVSS.n753 53.3664
R7201 AVSS.n794 AVSS.n752 53.3664
R7202 AVSS.n810 AVSS.n750 53.3664
R7203 AVSS.n814 AVSS.n748 53.3664
R7204 AVSS.n818 AVSS.n746 53.3664
R7205 AVSS.n822 AVSS.n744 53.3664
R7206 AVSS.n1043 AVSS.n990 53.3664
R7207 AVSS.n1040 AVSS.n979 53.3664
R7208 AVSS.n1036 AVSS.n981 53.3664
R7209 AVSS.n1032 AVSS.n983 53.3664
R7210 AVSS.n1021 AVSS.n986 53.3664
R7211 AVSS.n1017 AVSS.n987 53.3664
R7212 AVSS.n1013 AVSS.n988 53.3664
R7213 AVSS.n1009 AVSS.n989 53.3664
R7214 AVSS.n1062 AVSS.n1061 53.3664
R7215 AVSS.n997 AVSS.n980 53.3664
R7216 AVSS.n1001 AVSS.n982 53.3664
R7217 AVSS.n1005 AVSS.n984 53.3664
R7218 AVSS.n1060 AVSS.n1059 53.3664
R7219 AVSS.n995 AVSS.n993 53.3664
R7220 AVSS.n1054 AVSS.n992 53.3664
R7221 AVSS.n1050 AVSS.n991 53.3664
R7222 AVSS.n1060 AVSS.n994 53.3664
R7223 AVSS.n1055 AVSS.n993 53.3664
R7224 AVSS.n1051 AVSS.n992 53.3664
R7225 AVSS.n1047 AVSS.n991 53.3664
R7226 AVSS.n1029 AVSS.n983 53.3664
R7227 AVSS.n1033 AVSS.n981 53.3664
R7228 AVSS.n1037 AVSS.n979 53.3664
R7229 AVSS.n1041 AVSS.n990 53.3664
R7230 AVSS.n1012 AVSS.n989 53.3664
R7231 AVSS.n1016 AVSS.n988 53.3664
R7232 AVSS.n1020 AVSS.n987 53.3664
R7233 AVSS.n1024 AVSS.n986 53.3664
R7234 AVSS.n1008 AVSS.n984 53.3664
R7235 AVSS.n1004 AVSS.n982 53.3664
R7236 AVSS.n1000 AVSS.n980 53.3664
R7237 AVSS.n1061 AVSS.n978 53.3664
R7238 AVSS.n2488 AVSS.n2423 53.3664
R7239 AVSS.n2494 AVSS.n2493 53.3664
R7240 AVSS.n2497 AVSS.n2496 53.3664
R7241 AVSS.n2502 AVSS.n2501 53.3664
R7242 AVSS.n2489 AVSS.n2488 53.3664
R7243 AVSS.n2495 AVSS.n2494 53.3664
R7244 AVSS.n2496 AVSS.n2421 53.3664
R7245 AVSS.n2503 AVSS.n2502 53.3664
R7246 AVSS.n2487 AVSS.n2486 53.3664
R7247 AVSS.n2480 AVSS.n2425 53.3664
R7248 AVSS.n2479 AVSS.n2478 53.3664
R7249 AVSS.n2472 AVSS.n2427 53.3664
R7250 AVSS.n2473 AVSS.n2472 53.3664
R7251 AVSS.n2478 AVSS.n2477 53.3664
R7252 AVSS.n2481 AVSS.n2480 53.3664
R7253 AVSS.n2486 AVSS.n2485 53.3664
R7254 AVSS.n2465 AVSS.n2431 53.3664
R7255 AVSS.n2463 AVSS.n2462 53.3664
R7256 AVSS.n2458 AVSS.n2434 53.3664
R7257 AVSS.n2456 AVSS.n2455 53.3664
R7258 AVSS.n2457 AVSS.n2456 53.3664
R7259 AVSS.n2434 AVSS.n2432 53.3664
R7260 AVSS.n2464 AVSS.n2463 53.3664
R7261 AVSS.n2431 AVSS.n2429 53.3664
R7262 AVSS.n2439 AVSS.n2419 53.3664
R7263 AVSS.n2442 AVSS.n2441 53.3664
R7264 AVSS.n2447 AVSS.n2446 53.3664
R7265 AVSS.n2450 AVSS.n2449 53.3664
R7266 AVSS.n2449 AVSS.n2435 53.3664
R7267 AVSS.n2448 AVSS.n2447 53.3664
R7268 AVSS.n2441 AVSS.n2437 53.3664
R7269 AVSS.n2440 AVSS.n2439 53.3664
R7270 AVSS.n1936 AVSS.n1890 53.3664
R7271 AVSS.n1933 AVSS.n1891 53.3664
R7272 AVSS.n1929 AVSS.n1892 53.3664
R7273 AVSS.n1943 AVSS.n1902 53.3664
R7274 AVSS.n1947 AVSS.n1903 53.3664
R7275 AVSS.n1951 AVSS.n1904 53.3664
R7276 AVSS.n1955 AVSS.n1905 53.3664
R7277 AVSS.n1971 AVSS.n1970 53.3664
R7278 AVSS.n1966 AVSS.n1900 53.3664
R7279 AVSS.n1963 AVSS.n1899 53.3664
R7280 AVSS.n1959 AVSS.n1898 53.3664
R7281 AVSS.n1921 AVSS.n1897 53.3664
R7282 AVSS.n1917 AVSS.n1896 53.3664
R7283 AVSS.n1913 AVSS.n1895 53.3664
R7284 AVSS.n1909 AVSS.n1894 53.3664
R7285 AVSS.n1912 AVSS.n1894 53.3664
R7286 AVSS.n1916 AVSS.n1895 53.3664
R7287 AVSS.n1920 AVSS.n1896 53.3664
R7288 AVSS.n1923 AVSS.n1897 53.3664
R7289 AVSS.n1926 AVSS.n1892 53.3664
R7290 AVSS.n1930 AVSS.n1891 53.3664
R7291 AVSS.n1934 AVSS.n1890 53.3664
R7292 AVSS.n1946 AVSS.n1902 53.3664
R7293 AVSS.n1950 AVSS.n1903 53.3664
R7294 AVSS.n1954 AVSS.n1904 53.3664
R7295 AVSS.n1908 AVSS.n1905 53.3664
R7296 AVSS.n1898 AVSS.n1888 53.3664
R7297 AVSS.n1960 AVSS.n1899 53.3664
R7298 AVSS.n1964 AVSS.n1900 53.3664
R7299 AVSS.n1971 AVSS.n1907 53.3664
R7300 AVSS.n2556 AVSS.n2555 53.3664
R7301 AVSS.n1771 AVSS.n1769 53.3664
R7302 AVSS.n2550 AVSS.n1768 53.3664
R7303 AVSS.n2546 AVSS.n1767 53.3664
R7304 AVSS.n2556 AVSS.n1770 53.3664
R7305 AVSS.n2551 AVSS.n1769 53.3664
R7306 AVSS.n2547 AVSS.n1768 53.3664
R7307 AVSS.n2543 AVSS.n1767 53.3664
R7308 AVSS.n1784 AVSS.n1765 53.3664
R7309 AVSS.n1781 AVSS.n1755 53.3664
R7310 AVSS.n1777 AVSS.n1757 53.3664
R7311 AVSS.n1773 AVSS.n1759 53.3664
R7312 AVSS.n1759 AVSS.n1752 53.3664
R7313 AVSS.n1774 AVSS.n1757 53.3664
R7314 AVSS.n1778 AVSS.n1755 53.3664
R7315 AVSS.n1782 AVSS.n1765 53.3664
R7316 AVSS.n1792 AVSS.n1761 53.3664
R7317 AVSS.n1796 AVSS.n1762 53.3664
R7318 AVSS.n1800 AVSS.n1763 53.3664
R7319 AVSS.n1804 AVSS.n1764 53.3664
R7320 AVSS.n1801 AVSS.n1764 53.3664
R7321 AVSS.n1797 AVSS.n1763 53.3664
R7322 AVSS.n1793 AVSS.n1762 53.3664
R7323 AVSS.n1789 AVSS.n1761 53.3664
R7324 AVSS.n1820 AVSS.n1754 53.3664
R7325 AVSS.n1816 AVSS.n1756 53.3664
R7326 AVSS.n1812 AVSS.n1758 53.3664
R7327 AVSS.n1808 AVSS.n1760 53.3664
R7328 AVSS.n1805 AVSS.n1760 53.3664
R7329 AVSS.n1809 AVSS.n1758 53.3664
R7330 AVSS.n1813 AVSS.n1756 53.3664
R7331 AVSS.n1817 AVSS.n1754 53.3664
R7332 AVSS.n3339 AVSS.n3315 53.3664
R7333 AVSS.n3335 AVSS.n3314 53.3664
R7334 AVSS.n3331 AVSS.n3313 53.3664
R7335 AVSS.n3327 AVSS.n3312 53.3664
R7336 AVSS.n3330 AVSS.n3312 53.3664
R7337 AVSS.n3334 AVSS.n3313 53.3664
R7338 AVSS.n3338 AVSS.n3314 53.3664
R7339 AVSS.n3341 AVSS.n3315 53.3664
R7340 AVSS.n3390 AVSS.n3389 53.3664
R7341 AVSS.n3385 AVSS.n3318 53.3664
R7342 AVSS.n3382 AVSS.n3317 53.3664
R7343 AVSS.n3378 AVSS.n3316 53.3664
R7344 AVSS.n3362 AVSS.n3320 53.3664
R7345 AVSS.n3366 AVSS.n3321 53.3664
R7346 AVSS.n3370 AVSS.n3322 53.3664
R7347 AVSS.n3374 AVSS.n3323 53.3664
R7348 AVSS.n3355 AVSS.n3308 53.3664
R7349 AVSS.n3352 AVSS.n3309 53.3664
R7350 AVSS.n3348 AVSS.n3310 53.3664
R7351 AVSS.n3345 AVSS.n3310 53.3664
R7352 AVSS.n3349 AVSS.n3309 53.3664
R7353 AVSS.n3353 AVSS.n3308 53.3664
R7354 AVSS.n3365 AVSS.n3320 53.3664
R7355 AVSS.n3369 AVSS.n3321 53.3664
R7356 AVSS.n3373 AVSS.n3322 53.3664
R7357 AVSS.n3326 AVSS.n3323 53.3664
R7358 AVSS.n3316 AVSS.n3306 53.3664
R7359 AVSS.n3379 AVSS.n3317 53.3664
R7360 AVSS.n3383 AVSS.n3318 53.3664
R7361 AVSS.n3390 AVSS.n3325 53.3664
R7362 AVSS.t10 AVSS.n5961 51.7263
R7363 AVSS.t80 AVSS.n5016 51.443
R7364 AVSS.t76 AVSS.n1719 51.443
R7365 AVSS.t78 AVSS.n1071 51.443
R7366 AVSS.t84 AVSS.n151 51.443
R7367 AVSS.n5873 AVSS.t90 50.7749
R7368 AVSS.n4933 AVSS.t78 50.7749
R7369 AVSS.n4988 AVSS.t80 50.7749
R7370 AVSS.n4468 AVSS.t76 50.7749
R7371 AVSS.n5957 AVSS.n5944 48.7505
R7372 AVSS.n5944 AVSS.n5940 48.7505
R7373 AVSS.n5945 AVSS.n5943 48.7505
R7374 AVSS.n5943 AVSS.n5941 48.7505
R7375 AVSS.n6024 AVSS.n6008 48.7505
R7376 AVSS.n6019 AVSS.n6008 48.7505
R7377 AVSS.n6012 AVSS.n6011 48.7505
R7378 AVSS.n6019 AVSS.n6012 48.7505
R7379 AVSS.n6014 AVSS.n6013 48.4298
R7380 AVSS.n5978 AVSS.t42 45.9074
R7381 AVSS.t24 AVSS.t28 45.4029
R7382 AVSS.n5970 AVSS.t18 43.4116
R7383 AVSS.n5971 AVSS.t129 43.4116
R7384 AVSS.n6049 AVSS.t21 43.3991
R7385 AVSS.n6041 AVSS.t124 43.3991
R7386 AVSS.n290 AVSS.t29 43.2506
R7387 AVSS.n5975 AVSS.t8 43.2316
R7388 AVSS.n5973 AVSS.t125 43.2316
R7389 AVSS.n6045 AVSS.t31 43.2191
R7390 AVSS.n6048 AVSS.t26 43.1466
R7391 AVSS AVSS.t52 43.1141
R7392 AVSS AVSS.t49 43.0816
R7393 AVSS.n5983 AVSS.t45 42.9563
R7394 AVSS.n288 AVSS.t43 42.9316
R7395 AVSS AVSS.t41 42.9316
R7396 AVSS AVSS.t122 42.9197
R7397 AVSS.n6016 AVSS.n6014 42.8806
R7398 AVSS.n5979 AVSS.t36 41.8716
R7399 AVSS.n5979 AVSS.t33 41.8716
R7400 AVSS.n6018 AVSS.t24 41.8716
R7401 AVSS.n6021 AVSS.n6020 41.8716
R7402 AVSS.t127 AVSS.n6019 41.3672
R7403 AVSS.n6053 AVSS.n6052 39.0005
R7404 AVSS.n6054 AVSS.n6053 39.0005
R7405 AVSS.n6017 AVSS.n5933 39.0005
R7406 AVSS.n6018 AVSS.n6017 39.0005
R7407 AVSS.t28 AVSS.t130 38.3403
R7408 AVSS.t11 AVSS.n5978 37.8359
R7409 AVSS.n5986 AVSS.n5975 35.8673
R7410 AVSS.n5973 AVSS.n5969 35.8266
R7411 AVSS.n5970 AVSS.n5969 35.8266
R7412 AVSS.n6020 AVSS.n5928 34.3046
R7413 AVSS.n6021 AVSS.t48 32.7911
R7414 AVSS.t30 AVSS.n6016 31.7822
R7415 AVSS.n5995 AVSS.n5962 30.79
R7416 AVSS.n5966 AVSS.n5962 30.79
R7417 AVSS.n6060 AVSS.n6059 30.79
R7418 AVSS.n6059 AVSS.n6058 30.79
R7419 AVSS.n5963 AVSS.n5961 30.79
R7420 AVSS.n5981 AVSS.n5980 30.79
R7421 AVSS.n5980 AVSS.n5979 30.79
R7422 AVSS.n5984 AVSS.n5983 29.256
R7423 AVSS.n5977 AVSS.n5976 29.1418
R7424 AVSS.n5976 AVSS.n290 29.1418
R7425 AVSS.n138 AVSS.n136 27.5561
R7426 AVSS.n4186 AVSS.n4185 27.5561
R7427 AVSS.n4042 AVSS.n4001 27.5561
R7428 AVSS.n3831 AVSS.n3790 27.5561
R7429 AVSS.n3472 AVSS.n3431 27.5561
R7430 AVSS.n545 AVSS.n533 27.5561
R7431 AVSS.n1475 AVSS.n1442 27.5561
R7432 AVSS.n4895 AVSS.n4862 27.5561
R7433 AVSS.n2766 AVSS.n2764 27.5561
R7434 AVSS.n2644 AVSS.n2603 27.5561
R7435 AVSS.n1677 AVSS.n1636 27.5561
R7436 AVSS.n2062 AVSS.n2029 27.5561
R7437 AVSS.n1969 AVSS.n1957 27.5561
R7438 AVSS.n3388 AVSS.n3376 27.5561
R7439 AVSS.n5985 AVSS.n5984 26.7233
R7440 AVSS.n3492 AVSS.n3491 26.6672
R7441 AVSS.n5797 AVSS.n5796 26.6672
R7442 AVSS.n5525 AVSS.n5524 26.6672
R7443 AVSS.n5357 AVSS.n5312 26.6672
R7444 AVSS.n5158 AVSS.n5113 26.6672
R7445 AVSS.n517 AVSS.n516 26.6672
R7446 AVSS.n1426 AVSS.n1425 26.6672
R7447 AVSS.n4846 AVSS.n4845 26.6672
R7448 AVSS.n1697 AVSS.n1696 26.6672
R7449 AVSS.n2013 AVSS.n2012 26.6672
R7450 AVSS.n1045 AVSS.n1044 26.6672
R7451 AVSS.n2490 AVSS.n2424 26.6672
R7452 AVSS.n1941 AVSS.n1940 26.6672
R7453 AVSS.n3360 AVSS.n3359 26.6672
R7454 AVSS.n3872 AVSS.n188 26.074
R7455 AVSS.n4083 AVSS.n190 26.074
R7456 AVSS.n4103 AVSS.n192 26.074
R7457 AVSS.n3649 AVSS.n194 26.074
R7458 AVSS.n3412 AVSS.n2798 26.074
R7459 AVSS.n1615 AVSS.n1613 26.074
R7460 AVSS.n5020 AVSS.n5018 26.074
R7461 AVSS.n455 AVSS.n454 26.074
R7462 AVSS.n591 AVSS.n572 26.074
R7463 AVSS.n1112 AVSS.n1093 26.074
R7464 AVSS.n4497 AVSS.n4478 26.074
R7465 AVSS.n6236 AVSS.n38 26.074
R7466 AVSS.n6246 AVSS.n30 26.074
R7467 AVSS.n6265 AVSS.n21 26.074
R7468 AVSS.n5064 AVSS.n450 26.074
R7469 AVSS.n268 AVSS.n196 26.074
R7470 AVSS.t84 AVSS.n187 25.7843
R7471 AVSS.t84 AVSS.n189 25.7843
R7472 AVSS.t84 AVSS.n191 25.7843
R7473 AVSS.t84 AVSS.n193 25.7843
R7474 AVSS.t76 AVSS.n2797 25.7843
R7475 AVSS.n1602 AVSS.t78 25.7843
R7476 AVSS.t80 AVSS.n570 25.7843
R7477 AVSS.n5031 AVSS.t104 25.7843
R7478 AVSS.t80 AVSS.n571 25.7843
R7479 AVSS.t78 AVSS.n1092 25.7843
R7480 AVSS.t76 AVSS.n4477 25.7843
R7481 AVSS.n6237 AVSS.t106 25.7843
R7482 AVSS.t92 AVSS.n26 25.7843
R7483 AVSS.t89 AVSS.n20 25.7843
R7484 AVSS.t99 AVSS.n449 25.7843
R7485 AVSS.t84 AVSS.n195 25.7843
R7486 AVSS.n6036 AVSS.n6035 25.4353
R7487 AVSS.n6035 AVSS.n6034 25.4353
R7488 AVSS.n6032 AVSS.n6031 25.4353
R7489 AVSS.n6033 AVSS.n6032 25.4353
R7490 AVSS.n120 AVSS.n117 23.6449
R7491 AVSS.n4170 AVSS.n4168 23.6449
R7492 AVSS.n4027 AVSS.n4026 23.6449
R7493 AVSS.n3816 AVSS.n3815 23.6449
R7494 AVSS.n3457 AVSS.n3456 23.6449
R7495 AVSS.n5762 AVSS.n5759 23.6449
R7496 AVSS.n5490 AVSS.n5487 23.6449
R7497 AVSS.n3194 AVSS.n3191 23.6449
R7498 AVSS.n1270 AVSS.n1267 23.6449
R7499 AVSS.n4559 AVSS.n4556 23.6449
R7500 AVSS.n2748 AVSS.n2745 23.6449
R7501 AVSS.n2629 AVSS.n2628 23.6449
R7502 AVSS.n1662 AVSS.n1661 23.6449
R7503 AVSS.n811 AVSS.n808 23.6449
R7504 AVSS.n1010 AVSS.n1007 23.6449
R7505 AVSS.n5988 AVSS.n295 23.4005
R7506 AVSS.n5968 AVSS.n5967 23.4005
R7507 AVSS.n5978 AVSS.n5967 23.4005
R7508 AVSS.n5911 AVSS.t104 21.2535
R7509 AVSS.n5986 AVSS.n5985 20.832
R7510 AVSS.n5817 AVSS.n5816 20.0894
R7511 AVSS.n5545 AVSS.n5544 20.0894
R7512 AVSS.n5375 AVSS.n5374 20.0894
R7513 AVSS.n5176 AVSS.n5175 20.0894
R7514 AVSS.n3208 AVSS.n3160 20.0894
R7515 AVSS.n1284 AVSS.n1236 20.0894
R7516 AVSS.n4615 AVSS.n4614 20.0894
R7517 AVSS.n825 AVSS.n777 20.0894
R7518 AVSS.n1065 AVSS.n1064 20.0894
R7519 AVSS.n2508 AVSS.n2507 20.0894
R7520 AVSS.n2540 AVSS.n1822 20.0894
R7521 AVSS.n1294 AVSS.n1196 17.455
R7522 AVSS.n4624 AVSS.n1068 17.455
R7523 AVSS.n2114 AVSS.n2113 17.455
R7524 AVSS.n5570 AVSS.n5569 17.455
R7525 AVSS.n6278 AVSS.n6277 17.455
R7526 AVSS.n5092 AVSS.n5076 17.455
R7527 AVSS.n5923 AVSS.n302 17.455
R7528 AVSS.n5840 AVSS.n5625 17.455
R7529 AVSS.n693 AVSS.n683 17.455
R7530 AVSS.n2278 AVSS.n2277 17.455
R7531 AVSS.n2364 AVSS.n2363 17.455
R7532 AVSS.n1539 AVSS.n1538 17.455
R7533 AVSS.n921 AVSS.n920 17.455
R7534 AVSS.n3218 AVSS.n3121 17.455
R7535 AVSS.n4672 AVSS.n2776 17.455
R7536 AVSS.n4704 AVSS.n1723 17.455
R7537 AVSS.n2941 AVSS.n2914 17.455
R7538 AVSS.n4757 AVSS.n4733 17.455
R7539 AVSS.n2514 AVSS.n2512 17.455
R7540 AVSS.n232 AVSS.n148 17.455
R7541 AVSS.n4291 AVSS.n3889 17.455
R7542 AVSS.n4324 AVSS.n3678 17.455
R7543 AVSS.n3563 AVSS.n3536 17.455
R7544 AVSS.n4258 AVSS.n4206 17.455
R7545 AVSS.n4360 AVSS.n4358 17.455
R7546 AVSS.n101 AVSS.n100 17.4227
R7547 AVSS.n5779 AVSS.n5778 17.4227
R7548 AVSS.n5507 AVSS.n5506 17.4227
R7549 AVSS.n5335 AVSS.n5316 17.4227
R7550 AVSS.n5136 AVSS.n5117 17.4227
R7551 AVSS.n501 AVSS.n500 17.4227
R7552 AVSS.n3175 AVSS.n3174 17.4227
R7553 AVSS.n1251 AVSS.n1250 17.4227
R7554 AVSS.n4576 AVSS.n4575 17.4227
R7555 AVSS.n2729 AVSS.n2728 17.4227
R7556 AVSS.n792 AVSS.n791 17.4227
R7557 AVSS.n1027 AVSS.n1026 17.4227
R7558 AVSS.n2468 AVSS.n2428 17.4227
R7559 AVSS.n1925 AVSS.n1924 17.4227
R7560 AVSS.n5951 AVSS.t19 17.4005
R7561 AVSS.n5951 AVSS.t3 17.4005
R7562 AVSS.n5949 AVSS.t1 17.4005
R7563 AVSS.n5949 AVSS.t4 17.4005
R7564 AVSS.n1175 AVSS.n1173 16.9379
R7565 AVSS.n4648 AVSS.n4647 16.9379
R7566 AVSS.n2138 AVSS.n2137 16.9379
R7567 AVSS.n5871 AVSS.n5257 16.9379
R7568 AVSS.n6301 AVSS.n3 16.9379
R7569 AVSS.n5247 AVSS.n408 16.9379
R7570 AVSS.n396 AVSS.n395 16.9379
R7571 AVSS.n5629 AVSS.n5626 16.9379
R7572 AVSS.n716 AVSS.n684 16.9379
R7573 AVSS.n4986 AVSS.n973 16.9379
R7574 AVSS.n2341 AVSS.n2338 16.9379
R7575 AVSS.n1513 AVSS.n1512 16.9379
R7576 AVSS.n963 AVSS.n944 16.9379
R7577 AVSS.n3098 AVSS.n3097 16.9379
R7578 AVSS.n2860 AVSS.n2859 16.9379
R7579 AVSS.n3063 AVSS.n3012 16.9379
R7580 AVSS.n2963 AVSS.n2962 16.9379
R7581 AVSS.n4786 AVSS.n4724 16.9379
R7582 AVSS.n2537 AVSS.n1845 16.9379
R7583 AVSS.n6140 AVSS.n185 16.9379
R7584 AVSS.n3942 AVSS.n3941 16.9379
R7585 AVSS.n3731 AVSS.n3730 16.9379
R7586 AVSS.n3594 AVSS.n3593 16.9379
R7587 AVSS.n6135 AVSS.n213 16.9379
R7588 AVSS.n4466 AVSS.n3302 16.9379
R7589 AVSS.n146 AVSS.n145 16.7116
R7590 AVSS.n4204 AVSS.n4203 16.7116
R7591 AVSS.n4063 AVSS.n4062 16.7116
R7592 AVSS.n3852 AVSS.n3851 16.7116
R7593 AVSS.n3214 AVSS.n3213 16.7116
R7594 AVSS.n1290 AVSS.n1289 16.7116
R7595 AVSS.n4594 AVSS.n4593 16.7116
R7596 AVSS.n2774 AVSS.n2773 16.7116
R7597 AVSS.n2665 AVSS.n2664 16.7116
R7598 AVSS.n831 AVSS.n830 16.7116
R7599 AVSS.n1786 AVSS.n1785 16.7116
R7600 AVSS.t5 AVSS.t2 16.4491
R7601 AVSS.n78 AVSS.n56 16.0005
R7602 AVSS.n81 AVSS.n78 16.0005
R7603 AVSS.n82 AVSS.n81 16.0005
R7604 AVSS.n85 AVSS.n82 16.0005
R7605 AVSS.n86 AVSS.n85 16.0005
R7606 AVSS.n140 AVSS.n86 16.0005
R7607 AVSS.n140 AVSS.n139 16.0005
R7608 AVSS.n139 AVSS.n138 16.0005
R7609 AVSS.n136 AVSS.n133 16.0005
R7610 AVSS.n133 AVSS.n132 16.0005
R7611 AVSS.n132 AVSS.n129 16.0005
R7612 AVSS.n129 AVSS.n128 16.0005
R7613 AVSS.n128 AVSS.n125 16.0005
R7614 AVSS.n125 AVSS.n124 16.0005
R7615 AVSS.n124 AVSS.n121 16.0005
R7616 AVSS.n121 AVSS.n120 16.0005
R7617 AVSS.n104 AVSS.n101 16.0005
R7618 AVSS.n105 AVSS.n104 16.0005
R7619 AVSS.n108 AVSS.n105 16.0005
R7620 AVSS.n109 AVSS.n108 16.0005
R7621 AVSS.n112 AVSS.n109 16.0005
R7622 AVSS.n116 AVSS.n113 16.0005
R7623 AVSS.n117 AVSS.n116 16.0005
R7624 AVSS.n145 AVSS.n57 16.0005
R7625 AVSS.n88 AVSS.n57 16.0005
R7626 AVSS.n89 AVSS.n88 16.0005
R7627 AVSS.n92 AVSS.n89 16.0005
R7628 AVSS.n93 AVSS.n92 16.0005
R7629 AVSS.n96 AVSS.n93 16.0005
R7630 AVSS.n97 AVSS.n96 16.0005
R7631 AVSS.n100 AVSS.n97 16.0005
R7632 AVSS.n4199 AVSS.n4114 16.0005
R7633 AVSS.n4199 AVSS.n4198 16.0005
R7634 AVSS.n4198 AVSS.n4197 16.0005
R7635 AVSS.n4197 AVSS.n4194 16.0005
R7636 AVSS.n4194 AVSS.n4193 16.0005
R7637 AVSS.n4193 AVSS.n4190 16.0005
R7638 AVSS.n4190 AVSS.n4189 16.0005
R7639 AVSS.n4189 AVSS.n4186 16.0005
R7640 AVSS.n4185 AVSS.n4182 16.0005
R7641 AVSS.n4182 AVSS.n4181 16.0005
R7642 AVSS.n4181 AVSS.n4178 16.0005
R7643 AVSS.n4178 AVSS.n4177 16.0005
R7644 AVSS.n4177 AVSS.n4174 16.0005
R7645 AVSS.n4174 AVSS.n4173 16.0005
R7646 AVSS.n4173 AVSS.n4171 16.0005
R7647 AVSS.n4171 AVSS.n4170 16.0005
R7648 AVSS.n4153 AVSS.n4152 16.0005
R7649 AVSS.n4156 AVSS.n4153 16.0005
R7650 AVSS.n4157 AVSS.n4156 16.0005
R7651 AVSS.n4160 AVSS.n4157 16.0005
R7652 AVSS.n4161 AVSS.n4160 16.0005
R7653 AVSS.n4165 AVSS.n4164 16.0005
R7654 AVSS.n4168 AVSS.n4165 16.0005
R7655 AVSS.n4203 AVSS.n4115 16.0005
R7656 AVSS.n4137 AVSS.n4115 16.0005
R7657 AVSS.n4140 AVSS.n4137 16.0005
R7658 AVSS.n4141 AVSS.n4140 16.0005
R7659 AVSS.n4144 AVSS.n4141 16.0005
R7660 AVSS.n4145 AVSS.n4144 16.0005
R7661 AVSS.n4148 AVSS.n4145 16.0005
R7662 AVSS.n4149 AVSS.n4148 16.0005
R7663 AVSS.n4061 AVSS.n3997 16.0005
R7664 AVSS.n4056 AVSS.n3997 16.0005
R7665 AVSS.n4056 AVSS.n4055 16.0005
R7666 AVSS.n4055 AVSS.n3999 16.0005
R7667 AVSS.n4050 AVSS.n3999 16.0005
R7668 AVSS.n4050 AVSS.n4049 16.0005
R7669 AVSS.n4049 AVSS.n4048 16.0005
R7670 AVSS.n4048 AVSS.n4001 16.0005
R7671 AVSS.n4042 AVSS.n4041 16.0005
R7672 AVSS.n4041 AVSS.n4040 16.0005
R7673 AVSS.n4040 AVSS.n4003 16.0005
R7674 AVSS.n4034 AVSS.n4003 16.0005
R7675 AVSS.n4034 AVSS.n4033 16.0005
R7676 AVSS.n4033 AVSS.n4032 16.0005
R7677 AVSS.n4032 AVSS.n4005 16.0005
R7678 AVSS.n4027 AVSS.n4005 16.0005
R7679 AVSS.n4012 AVSS.n3990 16.0005
R7680 AVSS.n4013 AVSS.n4012 16.0005
R7681 AVSS.n4013 AVSS.n4009 16.0005
R7682 AVSS.n4019 AVSS.n4009 16.0005
R7683 AVSS.n4020 AVSS.n4019 16.0005
R7684 AVSS.n4021 AVSS.n4007 16.0005
R7685 AVSS.n4026 AVSS.n4007 16.0005
R7686 AVSS.n4064 AVSS.n4063 16.0005
R7687 AVSS.n4064 AVSS.n3995 16.0005
R7688 AVSS.n4070 AVSS.n3995 16.0005
R7689 AVSS.n4071 AVSS.n4070 16.0005
R7690 AVSS.n4072 AVSS.n4071 16.0005
R7691 AVSS.n4072 AVSS.n3993 16.0005
R7692 AVSS.n3993 AVSS.n3991 16.0005
R7693 AVSS.n4079 AVSS.n3991 16.0005
R7694 AVSS.n3850 AVSS.n3786 16.0005
R7695 AVSS.n3845 AVSS.n3786 16.0005
R7696 AVSS.n3845 AVSS.n3844 16.0005
R7697 AVSS.n3844 AVSS.n3788 16.0005
R7698 AVSS.n3839 AVSS.n3788 16.0005
R7699 AVSS.n3839 AVSS.n3838 16.0005
R7700 AVSS.n3838 AVSS.n3837 16.0005
R7701 AVSS.n3837 AVSS.n3790 16.0005
R7702 AVSS.n3831 AVSS.n3830 16.0005
R7703 AVSS.n3830 AVSS.n3829 16.0005
R7704 AVSS.n3829 AVSS.n3792 16.0005
R7705 AVSS.n3823 AVSS.n3792 16.0005
R7706 AVSS.n3823 AVSS.n3822 16.0005
R7707 AVSS.n3822 AVSS.n3821 16.0005
R7708 AVSS.n3821 AVSS.n3794 16.0005
R7709 AVSS.n3816 AVSS.n3794 16.0005
R7710 AVSS.n3801 AVSS.n3779 16.0005
R7711 AVSS.n3802 AVSS.n3801 16.0005
R7712 AVSS.n3802 AVSS.n3798 16.0005
R7713 AVSS.n3808 AVSS.n3798 16.0005
R7714 AVSS.n3809 AVSS.n3808 16.0005
R7715 AVSS.n3810 AVSS.n3796 16.0005
R7716 AVSS.n3815 AVSS.n3796 16.0005
R7717 AVSS.n3853 AVSS.n3852 16.0005
R7718 AVSS.n3853 AVSS.n3784 16.0005
R7719 AVSS.n3859 AVSS.n3784 16.0005
R7720 AVSS.n3860 AVSS.n3859 16.0005
R7721 AVSS.n3861 AVSS.n3860 16.0005
R7722 AVSS.n3861 AVSS.n3782 16.0005
R7723 AVSS.n3782 AVSS.n3780 16.0005
R7724 AVSS.n3868 AVSS.n3780 16.0005
R7725 AVSS.n3442 AVSS.n3420 16.0005
R7726 AVSS.n3443 AVSS.n3442 16.0005
R7727 AVSS.n3443 AVSS.n3439 16.0005
R7728 AVSS.n3449 AVSS.n3439 16.0005
R7729 AVSS.n3450 AVSS.n3449 16.0005
R7730 AVSS.n3451 AVSS.n3437 16.0005
R7731 AVSS.n3456 AVSS.n3437 16.0005
R7732 AVSS.n3472 AVSS.n3471 16.0005
R7733 AVSS.n3471 AVSS.n3470 16.0005
R7734 AVSS.n3470 AVSS.n3433 16.0005
R7735 AVSS.n3464 AVSS.n3433 16.0005
R7736 AVSS.n3464 AVSS.n3463 16.0005
R7737 AVSS.n3463 AVSS.n3462 16.0005
R7738 AVSS.n3462 AVSS.n3435 16.0005
R7739 AVSS.n3457 AVSS.n3435 16.0005
R7740 AVSS.n3491 AVSS.n3427 16.0005
R7741 AVSS.n3486 AVSS.n3427 16.0005
R7742 AVSS.n3486 AVSS.n3485 16.0005
R7743 AVSS.n3485 AVSS.n3429 16.0005
R7744 AVSS.n3480 AVSS.n3429 16.0005
R7745 AVSS.n3480 AVSS.n3479 16.0005
R7746 AVSS.n3479 AVSS.n3478 16.0005
R7747 AVSS.n3478 AVSS.n3431 16.0005
R7748 AVSS.n3493 AVSS.n3492 16.0005
R7749 AVSS.n3493 AVSS.n3425 16.0005
R7750 AVSS.n3499 AVSS.n3425 16.0005
R7751 AVSS.n3500 AVSS.n3499 16.0005
R7752 AVSS.n3501 AVSS.n3500 16.0005
R7753 AVSS.n3501 AVSS.n3423 16.0005
R7754 AVSS.n3423 AVSS.n3421 16.0005
R7755 AVSS.n3508 AVSS.n3421 16.0005
R7756 AVSS.n5810 AVSS.n5797 16.0005
R7757 AVSS.n5810 AVSS.n5809 16.0005
R7758 AVSS.n5809 AVSS.n5808 16.0005
R7759 AVSS.n5808 AVSS.n5805 16.0005
R7760 AVSS.n5805 AVSS.n5804 16.0005
R7761 AVSS.n5804 AVSS.n5801 16.0005
R7762 AVSS.n5801 AVSS.n5800 16.0005
R7763 AVSS.n5800 AVSS.n5727 16.0005
R7764 AVSS.n5796 AVSS.n5794 16.0005
R7765 AVSS.n5794 AVSS.n5791 16.0005
R7766 AVSS.n5791 AVSS.n5790 16.0005
R7767 AVSS.n5790 AVSS.n5787 16.0005
R7768 AVSS.n5787 AVSS.n5786 16.0005
R7769 AVSS.n5786 AVSS.n5783 16.0005
R7770 AVSS.n5783 AVSS.n5782 16.0005
R7771 AVSS.n5782 AVSS.n5779 16.0005
R7772 AVSS.n5778 AVSS.n5775 16.0005
R7773 AVSS.n5775 AVSS.n5774 16.0005
R7774 AVSS.n5774 AVSS.n5771 16.0005
R7775 AVSS.n5771 AVSS.n5770 16.0005
R7776 AVSS.n5770 AVSS.n5767 16.0005
R7777 AVSS.n5766 AVSS.n5763 16.0005
R7778 AVSS.n5763 AVSS.n5762 16.0005
R7779 AVSS.n5816 AVSS.n5728 16.0005
R7780 AVSS.n5748 AVSS.n5728 16.0005
R7781 AVSS.n5750 AVSS.n5748 16.0005
R7782 AVSS.n5751 AVSS.n5750 16.0005
R7783 AVSS.n5754 AVSS.n5751 16.0005
R7784 AVSS.n5755 AVSS.n5754 16.0005
R7785 AVSS.n5758 AVSS.n5755 16.0005
R7786 AVSS.n5759 AVSS.n5758 16.0005
R7787 AVSS.n5538 AVSS.n5525 16.0005
R7788 AVSS.n5538 AVSS.n5537 16.0005
R7789 AVSS.n5537 AVSS.n5536 16.0005
R7790 AVSS.n5536 AVSS.n5533 16.0005
R7791 AVSS.n5533 AVSS.n5532 16.0005
R7792 AVSS.n5532 AVSS.n5529 16.0005
R7793 AVSS.n5529 AVSS.n5528 16.0005
R7794 AVSS.n5528 AVSS.n5455 16.0005
R7795 AVSS.n5524 AVSS.n5522 16.0005
R7796 AVSS.n5522 AVSS.n5519 16.0005
R7797 AVSS.n5519 AVSS.n5518 16.0005
R7798 AVSS.n5518 AVSS.n5515 16.0005
R7799 AVSS.n5515 AVSS.n5514 16.0005
R7800 AVSS.n5514 AVSS.n5511 16.0005
R7801 AVSS.n5511 AVSS.n5510 16.0005
R7802 AVSS.n5510 AVSS.n5507 16.0005
R7803 AVSS.n5506 AVSS.n5503 16.0005
R7804 AVSS.n5503 AVSS.n5502 16.0005
R7805 AVSS.n5502 AVSS.n5499 16.0005
R7806 AVSS.n5499 AVSS.n5498 16.0005
R7807 AVSS.n5498 AVSS.n5495 16.0005
R7808 AVSS.n5494 AVSS.n5491 16.0005
R7809 AVSS.n5491 AVSS.n5490 16.0005
R7810 AVSS.n5544 AVSS.n5456 16.0005
R7811 AVSS.n5476 AVSS.n5456 16.0005
R7812 AVSS.n5478 AVSS.n5476 16.0005
R7813 AVSS.n5479 AVSS.n5478 16.0005
R7814 AVSS.n5482 AVSS.n5479 16.0005
R7815 AVSS.n5483 AVSS.n5482 16.0005
R7816 AVSS.n5486 AVSS.n5483 16.0005
R7817 AVSS.n5487 AVSS.n5486 16.0005
R7818 AVSS.n5335 AVSS.n5334 16.0005
R7819 AVSS.n5334 AVSS.n5333 16.0005
R7820 AVSS.n5333 AVSS.n5318 16.0005
R7821 AVSS.n5328 AVSS.n5318 16.0005
R7822 AVSS.n5328 AVSS.n5327 16.0005
R7823 AVSS.n5326 AVSS.n5321 16.0005
R7824 AVSS.n5321 AVSS.n5301 16.0005
R7825 AVSS.n5351 AVSS.n5312 16.0005
R7826 AVSS.n5351 AVSS.n5350 16.0005
R7827 AVSS.n5350 AVSS.n5349 16.0005
R7828 AVSS.n5349 AVSS.n5314 16.0005
R7829 AVSS.n5343 AVSS.n5314 16.0005
R7830 AVSS.n5343 AVSS.n5342 16.0005
R7831 AVSS.n5342 AVSS.n5341 16.0005
R7832 AVSS.n5341 AVSS.n5316 16.0005
R7833 AVSS.n5358 AVSS.n5357 16.0005
R7834 AVSS.n5359 AVSS.n5358 16.0005
R7835 AVSS.n5359 AVSS.n5310 16.0005
R7836 AVSS.n5365 AVSS.n5310 16.0005
R7837 AVSS.n5366 AVSS.n5365 16.0005
R7838 AVSS.n5367 AVSS.n5366 16.0005
R7839 AVSS.n5367 AVSS.n5308 16.0005
R7840 AVSS.n5373 AVSS.n5308 16.0005
R7841 AVSS.n5376 AVSS.n5375 16.0005
R7842 AVSS.n5376 AVSS.n5306 16.0005
R7843 AVSS.n5382 AVSS.n5306 16.0005
R7844 AVSS.n5383 AVSS.n5382 16.0005
R7845 AVSS.n5384 AVSS.n5383 16.0005
R7846 AVSS.n5384 AVSS.n5304 16.0005
R7847 AVSS.n5304 AVSS.n5302 16.0005
R7848 AVSS.n5391 AVSS.n5302 16.0005
R7849 AVSS.n5136 AVSS.n5135 16.0005
R7850 AVSS.n5135 AVSS.n5134 16.0005
R7851 AVSS.n5134 AVSS.n5119 16.0005
R7852 AVSS.n5129 AVSS.n5119 16.0005
R7853 AVSS.n5129 AVSS.n5128 16.0005
R7854 AVSS.n5127 AVSS.n5122 16.0005
R7855 AVSS.n5122 AVSS.n5102 16.0005
R7856 AVSS.n5152 AVSS.n5113 16.0005
R7857 AVSS.n5152 AVSS.n5151 16.0005
R7858 AVSS.n5151 AVSS.n5150 16.0005
R7859 AVSS.n5150 AVSS.n5115 16.0005
R7860 AVSS.n5144 AVSS.n5115 16.0005
R7861 AVSS.n5144 AVSS.n5143 16.0005
R7862 AVSS.n5143 AVSS.n5142 16.0005
R7863 AVSS.n5142 AVSS.n5117 16.0005
R7864 AVSS.n5159 AVSS.n5158 16.0005
R7865 AVSS.n5160 AVSS.n5159 16.0005
R7866 AVSS.n5160 AVSS.n5111 16.0005
R7867 AVSS.n5166 AVSS.n5111 16.0005
R7868 AVSS.n5167 AVSS.n5166 16.0005
R7869 AVSS.n5168 AVSS.n5167 16.0005
R7870 AVSS.n5168 AVSS.n5109 16.0005
R7871 AVSS.n5174 AVSS.n5109 16.0005
R7872 AVSS.n5177 AVSS.n5176 16.0005
R7873 AVSS.n5177 AVSS.n5107 16.0005
R7874 AVSS.n5183 AVSS.n5107 16.0005
R7875 AVSS.n5184 AVSS.n5183 16.0005
R7876 AVSS.n5185 AVSS.n5184 16.0005
R7877 AVSS.n5185 AVSS.n5105 16.0005
R7878 AVSS.n5105 AVSS.n5103 16.0005
R7879 AVSS.n5192 AVSS.n5103 16.0005
R7880 AVSS.n500 AVSS.n498 16.0005
R7881 AVSS.n498 AVSS.n495 16.0005
R7882 AVSS.n495 AVSS.n494 16.0005
R7883 AVSS.n494 AVSS.n491 16.0005
R7884 AVSS.n491 AVSS.n490 16.0005
R7885 AVSS.n487 AVSS.n486 16.0005
R7886 AVSS.n486 AVSS.n462 16.0005
R7887 AVSS.n516 AVSS.n514 16.0005
R7888 AVSS.n514 AVSS.n513 16.0005
R7889 AVSS.n513 AVSS.n511 16.0005
R7890 AVSS.n511 AVSS.n508 16.0005
R7891 AVSS.n508 AVSS.n507 16.0005
R7892 AVSS.n507 AVSS.n504 16.0005
R7893 AVSS.n504 AVSS.n503 16.0005
R7894 AVSS.n503 AVSS.n501 16.0005
R7895 AVSS.n520 AVSS.n517 16.0005
R7896 AVSS.n521 AVSS.n520 16.0005
R7897 AVSS.n524 AVSS.n521 16.0005
R7898 AVSS.n525 AVSS.n524 16.0005
R7899 AVSS.n528 AVSS.n525 16.0005
R7900 AVSS.n529 AVSS.n528 16.0005
R7901 AVSS.n532 AVSS.n529 16.0005
R7902 AVSS.n533 AVSS.n532 16.0005
R7903 AVSS.n545 AVSS.n544 16.0005
R7904 AVSS.n544 AVSS.n543 16.0005
R7905 AVSS.n543 AVSS.n541 16.0005
R7906 AVSS.n541 AVSS.n538 16.0005
R7907 AVSS.n538 AVSS.n537 16.0005
R7908 AVSS.n537 AVSS.n534 16.0005
R7909 AVSS.n534 AVSS.n463 16.0005
R7910 AVSS.n550 AVSS.n463 16.0005
R7911 AVSS.n1443 AVSS.n1390 16.0005
R7912 AVSS.n1446 AVSS.n1443 16.0005
R7913 AVSS.n1447 AVSS.n1446 16.0005
R7914 AVSS.n1450 AVSS.n1447 16.0005
R7915 AVSS.n1451 AVSS.n1450 16.0005
R7916 AVSS.n1455 AVSS.n1454 16.0005
R7917 AVSS.n1458 AVSS.n1455 16.0005
R7918 AVSS.n1425 AVSS.n1423 16.0005
R7919 AVSS.n1423 AVSS.n1422 16.0005
R7920 AVSS.n1422 AVSS.n1420 16.0005
R7921 AVSS.n1420 AVSS.n1417 16.0005
R7922 AVSS.n1417 AVSS.n1416 16.0005
R7923 AVSS.n1416 AVSS.n1413 16.0005
R7924 AVSS.n1413 AVSS.n1391 16.0005
R7925 AVSS.n1479 AVSS.n1391 16.0005
R7926 AVSS.n1429 AVSS.n1426 16.0005
R7927 AVSS.n1430 AVSS.n1429 16.0005
R7928 AVSS.n1433 AVSS.n1430 16.0005
R7929 AVSS.n1434 AVSS.n1433 16.0005
R7930 AVSS.n1437 AVSS.n1434 16.0005
R7931 AVSS.n1438 AVSS.n1437 16.0005
R7932 AVSS.n1441 AVSS.n1438 16.0005
R7933 AVSS.n1442 AVSS.n1441 16.0005
R7934 AVSS.n1475 AVSS.n1474 16.0005
R7935 AVSS.n1474 AVSS.n1473 16.0005
R7936 AVSS.n1473 AVSS.n1471 16.0005
R7937 AVSS.n1471 AVSS.n1468 16.0005
R7938 AVSS.n1468 AVSS.n1467 16.0005
R7939 AVSS.n1467 AVSS.n1464 16.0005
R7940 AVSS.n1464 AVSS.n1463 16.0005
R7941 AVSS.n1463 AVSS.n1460 16.0005
R7942 AVSS.n4863 AVSS.n4810 16.0005
R7943 AVSS.n4866 AVSS.n4863 16.0005
R7944 AVSS.n4867 AVSS.n4866 16.0005
R7945 AVSS.n4870 AVSS.n4867 16.0005
R7946 AVSS.n4871 AVSS.n4870 16.0005
R7947 AVSS.n4875 AVSS.n4874 16.0005
R7948 AVSS.n4878 AVSS.n4875 16.0005
R7949 AVSS.n4845 AVSS.n4843 16.0005
R7950 AVSS.n4843 AVSS.n4842 16.0005
R7951 AVSS.n4842 AVSS.n4840 16.0005
R7952 AVSS.n4840 AVSS.n4837 16.0005
R7953 AVSS.n4837 AVSS.n4836 16.0005
R7954 AVSS.n4836 AVSS.n4833 16.0005
R7955 AVSS.n4833 AVSS.n4811 16.0005
R7956 AVSS.n4899 AVSS.n4811 16.0005
R7957 AVSS.n4849 AVSS.n4846 16.0005
R7958 AVSS.n4850 AVSS.n4849 16.0005
R7959 AVSS.n4853 AVSS.n4850 16.0005
R7960 AVSS.n4854 AVSS.n4853 16.0005
R7961 AVSS.n4857 AVSS.n4854 16.0005
R7962 AVSS.n4858 AVSS.n4857 16.0005
R7963 AVSS.n4861 AVSS.n4858 16.0005
R7964 AVSS.n4862 AVSS.n4861 16.0005
R7965 AVSS.n4895 AVSS.n4894 16.0005
R7966 AVSS.n4894 AVSS.n4893 16.0005
R7967 AVSS.n4893 AVSS.n4891 16.0005
R7968 AVSS.n4891 AVSS.n4888 16.0005
R7969 AVSS.n4888 AVSS.n4887 16.0005
R7970 AVSS.n4887 AVSS.n4884 16.0005
R7971 AVSS.n4884 AVSS.n4883 16.0005
R7972 AVSS.n4883 AVSS.n4880 16.0005
R7973 AVSS.n3145 AVSS.n3123 16.0005
R7974 AVSS.n3148 AVSS.n3145 16.0005
R7975 AVSS.n3149 AVSS.n3148 16.0005
R7976 AVSS.n3152 AVSS.n3149 16.0005
R7977 AVSS.n3153 AVSS.n3152 16.0005
R7978 AVSS.n3156 AVSS.n3153 16.0005
R7979 AVSS.n3158 AVSS.n3156 16.0005
R7980 AVSS.n3159 AVSS.n3158 16.0005
R7981 AVSS.n3213 AVSS.n3124 16.0005
R7982 AVSS.n3162 AVSS.n3124 16.0005
R7983 AVSS.n3163 AVSS.n3162 16.0005
R7984 AVSS.n3166 AVSS.n3163 16.0005
R7985 AVSS.n3167 AVSS.n3166 16.0005
R7986 AVSS.n3170 AVSS.n3167 16.0005
R7987 AVSS.n3171 AVSS.n3170 16.0005
R7988 AVSS.n3174 AVSS.n3171 16.0005
R7989 AVSS.n3178 AVSS.n3175 16.0005
R7990 AVSS.n3179 AVSS.n3178 16.0005
R7991 AVSS.n3182 AVSS.n3179 16.0005
R7992 AVSS.n3183 AVSS.n3182 16.0005
R7993 AVSS.n3186 AVSS.n3183 16.0005
R7994 AVSS.n3190 AVSS.n3187 16.0005
R7995 AVSS.n3191 AVSS.n3190 16.0005
R7996 AVSS.n3208 AVSS.n3207 16.0005
R7997 AVSS.n3207 AVSS.n3206 16.0005
R7998 AVSS.n3206 AVSS.n3203 16.0005
R7999 AVSS.n3203 AVSS.n3202 16.0005
R8000 AVSS.n3202 AVSS.n3199 16.0005
R8001 AVSS.n3199 AVSS.n3198 16.0005
R8002 AVSS.n3198 AVSS.n3195 16.0005
R8003 AVSS.n3195 AVSS.n3194 16.0005
R8004 AVSS.n1221 AVSS.n1199 16.0005
R8005 AVSS.n1224 AVSS.n1221 16.0005
R8006 AVSS.n1225 AVSS.n1224 16.0005
R8007 AVSS.n1228 AVSS.n1225 16.0005
R8008 AVSS.n1229 AVSS.n1228 16.0005
R8009 AVSS.n1232 AVSS.n1229 16.0005
R8010 AVSS.n1234 AVSS.n1232 16.0005
R8011 AVSS.n1235 AVSS.n1234 16.0005
R8012 AVSS.n1289 AVSS.n1200 16.0005
R8013 AVSS.n1238 AVSS.n1200 16.0005
R8014 AVSS.n1239 AVSS.n1238 16.0005
R8015 AVSS.n1242 AVSS.n1239 16.0005
R8016 AVSS.n1243 AVSS.n1242 16.0005
R8017 AVSS.n1246 AVSS.n1243 16.0005
R8018 AVSS.n1247 AVSS.n1246 16.0005
R8019 AVSS.n1250 AVSS.n1247 16.0005
R8020 AVSS.n1254 AVSS.n1251 16.0005
R8021 AVSS.n1255 AVSS.n1254 16.0005
R8022 AVSS.n1258 AVSS.n1255 16.0005
R8023 AVSS.n1259 AVSS.n1258 16.0005
R8024 AVSS.n1262 AVSS.n1259 16.0005
R8025 AVSS.n1266 AVSS.n1263 16.0005
R8026 AVSS.n1267 AVSS.n1266 16.0005
R8027 AVSS.n1284 AVSS.n1283 16.0005
R8028 AVSS.n1283 AVSS.n1282 16.0005
R8029 AVSS.n1282 AVSS.n1279 16.0005
R8030 AVSS.n1279 AVSS.n1278 16.0005
R8031 AVSS.n1278 AVSS.n1275 16.0005
R8032 AVSS.n1275 AVSS.n1274 16.0005
R8033 AVSS.n1274 AVSS.n1271 16.0005
R8034 AVSS.n1271 AVSS.n1270 16.0005
R8035 AVSS.n4608 AVSS.n4595 16.0005
R8036 AVSS.n4608 AVSS.n4607 16.0005
R8037 AVSS.n4607 AVSS.n4606 16.0005
R8038 AVSS.n4606 AVSS.n4603 16.0005
R8039 AVSS.n4603 AVSS.n4602 16.0005
R8040 AVSS.n4602 AVSS.n4599 16.0005
R8041 AVSS.n4599 AVSS.n4598 16.0005
R8042 AVSS.n4598 AVSS.n4524 16.0005
R8043 AVSS.n4593 AVSS.n4591 16.0005
R8044 AVSS.n4591 AVSS.n4588 16.0005
R8045 AVSS.n4588 AVSS.n4587 16.0005
R8046 AVSS.n4587 AVSS.n4584 16.0005
R8047 AVSS.n4584 AVSS.n4583 16.0005
R8048 AVSS.n4583 AVSS.n4580 16.0005
R8049 AVSS.n4580 AVSS.n4579 16.0005
R8050 AVSS.n4579 AVSS.n4576 16.0005
R8051 AVSS.n4575 AVSS.n4572 16.0005
R8052 AVSS.n4572 AVSS.n4571 16.0005
R8053 AVSS.n4571 AVSS.n4568 16.0005
R8054 AVSS.n4568 AVSS.n4567 16.0005
R8055 AVSS.n4567 AVSS.n4564 16.0005
R8056 AVSS.n4563 AVSS.n4560 16.0005
R8057 AVSS.n4560 AVSS.n4559 16.0005
R8058 AVSS.n4614 AVSS.n4525 16.0005
R8059 AVSS.n4545 AVSS.n4525 16.0005
R8060 AVSS.n4547 AVSS.n4545 16.0005
R8061 AVSS.n4548 AVSS.n4547 16.0005
R8062 AVSS.n4551 AVSS.n4548 16.0005
R8063 AVSS.n4552 AVSS.n4551 16.0005
R8064 AVSS.n4555 AVSS.n4552 16.0005
R8065 AVSS.n4556 AVSS.n4555 16.0005
R8066 AVSS.n2706 AVSS.n2684 16.0005
R8067 AVSS.n2709 AVSS.n2706 16.0005
R8068 AVSS.n2710 AVSS.n2709 16.0005
R8069 AVSS.n2713 AVSS.n2710 16.0005
R8070 AVSS.n2714 AVSS.n2713 16.0005
R8071 AVSS.n2768 AVSS.n2714 16.0005
R8072 AVSS.n2768 AVSS.n2767 16.0005
R8073 AVSS.n2767 AVSS.n2766 16.0005
R8074 AVSS.n2764 AVSS.n2761 16.0005
R8075 AVSS.n2761 AVSS.n2760 16.0005
R8076 AVSS.n2760 AVSS.n2757 16.0005
R8077 AVSS.n2757 AVSS.n2756 16.0005
R8078 AVSS.n2756 AVSS.n2753 16.0005
R8079 AVSS.n2753 AVSS.n2752 16.0005
R8080 AVSS.n2752 AVSS.n2749 16.0005
R8081 AVSS.n2749 AVSS.n2748 16.0005
R8082 AVSS.n2732 AVSS.n2729 16.0005
R8083 AVSS.n2733 AVSS.n2732 16.0005
R8084 AVSS.n2736 AVSS.n2733 16.0005
R8085 AVSS.n2737 AVSS.n2736 16.0005
R8086 AVSS.n2740 AVSS.n2737 16.0005
R8087 AVSS.n2744 AVSS.n2741 16.0005
R8088 AVSS.n2745 AVSS.n2744 16.0005
R8089 AVSS.n2773 AVSS.n2685 16.0005
R8090 AVSS.n2716 AVSS.n2685 16.0005
R8091 AVSS.n2717 AVSS.n2716 16.0005
R8092 AVSS.n2720 AVSS.n2717 16.0005
R8093 AVSS.n2721 AVSS.n2720 16.0005
R8094 AVSS.n2724 AVSS.n2721 16.0005
R8095 AVSS.n2725 AVSS.n2724 16.0005
R8096 AVSS.n2728 AVSS.n2725 16.0005
R8097 AVSS.n2663 AVSS.n2599 16.0005
R8098 AVSS.n2658 AVSS.n2599 16.0005
R8099 AVSS.n2658 AVSS.n2657 16.0005
R8100 AVSS.n2657 AVSS.n2601 16.0005
R8101 AVSS.n2652 AVSS.n2601 16.0005
R8102 AVSS.n2652 AVSS.n2651 16.0005
R8103 AVSS.n2651 AVSS.n2650 16.0005
R8104 AVSS.n2650 AVSS.n2603 16.0005
R8105 AVSS.n2644 AVSS.n2643 16.0005
R8106 AVSS.n2643 AVSS.n2642 16.0005
R8107 AVSS.n2642 AVSS.n2605 16.0005
R8108 AVSS.n2636 AVSS.n2605 16.0005
R8109 AVSS.n2636 AVSS.n2635 16.0005
R8110 AVSS.n2635 AVSS.n2634 16.0005
R8111 AVSS.n2634 AVSS.n2607 16.0005
R8112 AVSS.n2629 AVSS.n2607 16.0005
R8113 AVSS.n2614 AVSS.n2592 16.0005
R8114 AVSS.n2615 AVSS.n2614 16.0005
R8115 AVSS.n2615 AVSS.n2611 16.0005
R8116 AVSS.n2621 AVSS.n2611 16.0005
R8117 AVSS.n2622 AVSS.n2621 16.0005
R8118 AVSS.n2623 AVSS.n2609 16.0005
R8119 AVSS.n2628 AVSS.n2609 16.0005
R8120 AVSS.n2666 AVSS.n2665 16.0005
R8121 AVSS.n2666 AVSS.n2597 16.0005
R8122 AVSS.n2672 AVSS.n2597 16.0005
R8123 AVSS.n2673 AVSS.n2672 16.0005
R8124 AVSS.n2674 AVSS.n2673 16.0005
R8125 AVSS.n2674 AVSS.n2595 16.0005
R8126 AVSS.n2595 AVSS.n2593 16.0005
R8127 AVSS.n2681 AVSS.n2593 16.0005
R8128 AVSS.n1647 AVSS.n1625 16.0005
R8129 AVSS.n1648 AVSS.n1647 16.0005
R8130 AVSS.n1648 AVSS.n1644 16.0005
R8131 AVSS.n1654 AVSS.n1644 16.0005
R8132 AVSS.n1655 AVSS.n1654 16.0005
R8133 AVSS.n1656 AVSS.n1642 16.0005
R8134 AVSS.n1661 AVSS.n1642 16.0005
R8135 AVSS.n1677 AVSS.n1676 16.0005
R8136 AVSS.n1676 AVSS.n1675 16.0005
R8137 AVSS.n1675 AVSS.n1638 16.0005
R8138 AVSS.n1669 AVSS.n1638 16.0005
R8139 AVSS.n1669 AVSS.n1668 16.0005
R8140 AVSS.n1668 AVSS.n1667 16.0005
R8141 AVSS.n1667 AVSS.n1640 16.0005
R8142 AVSS.n1662 AVSS.n1640 16.0005
R8143 AVSS.n1696 AVSS.n1632 16.0005
R8144 AVSS.n1691 AVSS.n1632 16.0005
R8145 AVSS.n1691 AVSS.n1690 16.0005
R8146 AVSS.n1690 AVSS.n1634 16.0005
R8147 AVSS.n1685 AVSS.n1634 16.0005
R8148 AVSS.n1685 AVSS.n1684 16.0005
R8149 AVSS.n1684 AVSS.n1683 16.0005
R8150 AVSS.n1683 AVSS.n1636 16.0005
R8151 AVSS.n1698 AVSS.n1697 16.0005
R8152 AVSS.n1698 AVSS.n1630 16.0005
R8153 AVSS.n1704 AVSS.n1630 16.0005
R8154 AVSS.n1705 AVSS.n1704 16.0005
R8155 AVSS.n1706 AVSS.n1705 16.0005
R8156 AVSS.n1706 AVSS.n1628 16.0005
R8157 AVSS.n1628 AVSS.n1626 16.0005
R8158 AVSS.n1713 AVSS.n1626 16.0005
R8159 AVSS.n1790 AVSS.n1750 16.0005
R8160 AVSS.n1791 AVSS.n1790 16.0005
R8161 AVSS.n1794 AVSS.n1791 16.0005
R8162 AVSS.n1795 AVSS.n1794 16.0005
R8163 AVSS.n1798 AVSS.n1795 16.0005
R8164 AVSS.n1802 AVSS.n1799 16.0005
R8165 AVSS.n1803 AVSS.n1802 16.0005
R8166 AVSS.n2030 AVSS.n1977 16.0005
R8167 AVSS.n2033 AVSS.n2030 16.0005
R8168 AVSS.n2034 AVSS.n2033 16.0005
R8169 AVSS.n2037 AVSS.n2034 16.0005
R8170 AVSS.n2038 AVSS.n2037 16.0005
R8171 AVSS.n2042 AVSS.n2041 16.0005
R8172 AVSS.n2045 AVSS.n2042 16.0005
R8173 AVSS.n2012 AVSS.n2010 16.0005
R8174 AVSS.n2010 AVSS.n2009 16.0005
R8175 AVSS.n2009 AVSS.n2007 16.0005
R8176 AVSS.n2007 AVSS.n2004 16.0005
R8177 AVSS.n2004 AVSS.n2003 16.0005
R8178 AVSS.n2003 AVSS.n2000 16.0005
R8179 AVSS.n2000 AVSS.n1978 16.0005
R8180 AVSS.n2066 AVSS.n1978 16.0005
R8181 AVSS.n2016 AVSS.n2013 16.0005
R8182 AVSS.n2017 AVSS.n2016 16.0005
R8183 AVSS.n2020 AVSS.n2017 16.0005
R8184 AVSS.n2021 AVSS.n2020 16.0005
R8185 AVSS.n2024 AVSS.n2021 16.0005
R8186 AVSS.n2025 AVSS.n2024 16.0005
R8187 AVSS.n2028 AVSS.n2025 16.0005
R8188 AVSS.n2029 AVSS.n2028 16.0005
R8189 AVSS.n2062 AVSS.n2061 16.0005
R8190 AVSS.n2061 AVSS.n2060 16.0005
R8191 AVSS.n2060 AVSS.n2058 16.0005
R8192 AVSS.n2058 AVSS.n2055 16.0005
R8193 AVSS.n2055 AVSS.n2054 16.0005
R8194 AVSS.n2054 AVSS.n2051 16.0005
R8195 AVSS.n2051 AVSS.n2050 16.0005
R8196 AVSS.n2050 AVSS.n2047 16.0005
R8197 AVSS.n762 AVSS.n740 16.0005
R8198 AVSS.n765 AVSS.n762 16.0005
R8199 AVSS.n766 AVSS.n765 16.0005
R8200 AVSS.n769 AVSS.n766 16.0005
R8201 AVSS.n770 AVSS.n769 16.0005
R8202 AVSS.n773 AVSS.n770 16.0005
R8203 AVSS.n775 AVSS.n773 16.0005
R8204 AVSS.n776 AVSS.n775 16.0005
R8205 AVSS.n830 AVSS.n741 16.0005
R8206 AVSS.n779 AVSS.n741 16.0005
R8207 AVSS.n780 AVSS.n779 16.0005
R8208 AVSS.n783 AVSS.n780 16.0005
R8209 AVSS.n784 AVSS.n783 16.0005
R8210 AVSS.n787 AVSS.n784 16.0005
R8211 AVSS.n788 AVSS.n787 16.0005
R8212 AVSS.n791 AVSS.n788 16.0005
R8213 AVSS.n795 AVSS.n792 16.0005
R8214 AVSS.n796 AVSS.n795 16.0005
R8215 AVSS.n799 AVSS.n796 16.0005
R8216 AVSS.n800 AVSS.n799 16.0005
R8217 AVSS.n803 AVSS.n800 16.0005
R8218 AVSS.n807 AVSS.n804 16.0005
R8219 AVSS.n808 AVSS.n807 16.0005
R8220 AVSS.n825 AVSS.n824 16.0005
R8221 AVSS.n824 AVSS.n823 16.0005
R8222 AVSS.n823 AVSS.n820 16.0005
R8223 AVSS.n820 AVSS.n819 16.0005
R8224 AVSS.n819 AVSS.n816 16.0005
R8225 AVSS.n816 AVSS.n815 16.0005
R8226 AVSS.n815 AVSS.n812 16.0005
R8227 AVSS.n812 AVSS.n811 16.0005
R8228 AVSS.n1058 AVSS.n1045 16.0005
R8229 AVSS.n1058 AVSS.n1057 16.0005
R8230 AVSS.n1057 AVSS.n1056 16.0005
R8231 AVSS.n1056 AVSS.n1053 16.0005
R8232 AVSS.n1053 AVSS.n1052 16.0005
R8233 AVSS.n1052 AVSS.n1049 16.0005
R8234 AVSS.n1049 AVSS.n1048 16.0005
R8235 AVSS.n1048 AVSS.n975 16.0005
R8236 AVSS.n1044 AVSS.n1042 16.0005
R8237 AVSS.n1042 AVSS.n1039 16.0005
R8238 AVSS.n1039 AVSS.n1038 16.0005
R8239 AVSS.n1038 AVSS.n1035 16.0005
R8240 AVSS.n1035 AVSS.n1034 16.0005
R8241 AVSS.n1034 AVSS.n1031 16.0005
R8242 AVSS.n1031 AVSS.n1030 16.0005
R8243 AVSS.n1030 AVSS.n1027 16.0005
R8244 AVSS.n1026 AVSS.n1023 16.0005
R8245 AVSS.n1023 AVSS.n1022 16.0005
R8246 AVSS.n1022 AVSS.n1019 16.0005
R8247 AVSS.n1019 AVSS.n1018 16.0005
R8248 AVSS.n1018 AVSS.n1015 16.0005
R8249 AVSS.n1014 AVSS.n1011 16.0005
R8250 AVSS.n1011 AVSS.n1010 16.0005
R8251 AVSS.n1064 AVSS.n976 16.0005
R8252 AVSS.n996 AVSS.n976 16.0005
R8253 AVSS.n998 AVSS.n996 16.0005
R8254 AVSS.n999 AVSS.n998 16.0005
R8255 AVSS.n1002 AVSS.n999 16.0005
R8256 AVSS.n1003 AVSS.n1002 16.0005
R8257 AVSS.n1006 AVSS.n1003 16.0005
R8258 AVSS.n1007 AVSS.n1006 16.0005
R8259 AVSS.n2468 AVSS.n2467 16.0005
R8260 AVSS.n2467 AVSS.n2466 16.0005
R8261 AVSS.n2466 AVSS.n2430 16.0005
R8262 AVSS.n2461 AVSS.n2430 16.0005
R8263 AVSS.n2461 AVSS.n2460 16.0005
R8264 AVSS.n2459 AVSS.n2433 16.0005
R8265 AVSS.n2454 AVSS.n2433 16.0005
R8266 AVSS.n2484 AVSS.n2424 16.0005
R8267 AVSS.n2484 AVSS.n2483 16.0005
R8268 AVSS.n2483 AVSS.n2482 16.0005
R8269 AVSS.n2482 AVSS.n2426 16.0005
R8270 AVSS.n2476 AVSS.n2426 16.0005
R8271 AVSS.n2476 AVSS.n2475 16.0005
R8272 AVSS.n2475 AVSS.n2474 16.0005
R8273 AVSS.n2474 AVSS.n2428 16.0005
R8274 AVSS.n2491 AVSS.n2490 16.0005
R8275 AVSS.n2492 AVSS.n2491 16.0005
R8276 AVSS.n2492 AVSS.n2422 16.0005
R8277 AVSS.n2498 AVSS.n2422 16.0005
R8278 AVSS.n2499 AVSS.n2498 16.0005
R8279 AVSS.n2500 AVSS.n2499 16.0005
R8280 AVSS.n2500 AVSS.n2420 16.0005
R8281 AVSS.n2420 AVSS.n2417 16.0005
R8282 AVSS.n2507 AVSS.n2418 16.0005
R8283 AVSS.n2438 AVSS.n2418 16.0005
R8284 AVSS.n2443 AVSS.n2438 16.0005
R8285 AVSS.n2444 AVSS.n2443 16.0005
R8286 AVSS.n2445 AVSS.n2444 16.0005
R8287 AVSS.n2445 AVSS.n2436 16.0005
R8288 AVSS.n2451 AVSS.n2436 16.0005
R8289 AVSS.n2452 AVSS.n2451 16.0005
R8290 AVSS.n1924 AVSS.n1922 16.0005
R8291 AVSS.n1922 AVSS.n1919 16.0005
R8292 AVSS.n1919 AVSS.n1918 16.0005
R8293 AVSS.n1918 AVSS.n1915 16.0005
R8294 AVSS.n1915 AVSS.n1914 16.0005
R8295 AVSS.n1911 AVSS.n1910 16.0005
R8296 AVSS.n1910 AVSS.n1886 16.0005
R8297 AVSS.n1940 AVSS.n1938 16.0005
R8298 AVSS.n1938 AVSS.n1937 16.0005
R8299 AVSS.n1937 AVSS.n1935 16.0005
R8300 AVSS.n1935 AVSS.n1932 16.0005
R8301 AVSS.n1932 AVSS.n1931 16.0005
R8302 AVSS.n1931 AVSS.n1928 16.0005
R8303 AVSS.n1928 AVSS.n1927 16.0005
R8304 AVSS.n1927 AVSS.n1925 16.0005
R8305 AVSS.n1944 AVSS.n1941 16.0005
R8306 AVSS.n1945 AVSS.n1944 16.0005
R8307 AVSS.n1948 AVSS.n1945 16.0005
R8308 AVSS.n1949 AVSS.n1948 16.0005
R8309 AVSS.n1952 AVSS.n1949 16.0005
R8310 AVSS.n1953 AVSS.n1952 16.0005
R8311 AVSS.n1956 AVSS.n1953 16.0005
R8312 AVSS.n1957 AVSS.n1956 16.0005
R8313 AVSS.n1969 AVSS.n1968 16.0005
R8314 AVSS.n1968 AVSS.n1967 16.0005
R8315 AVSS.n1967 AVSS.n1965 16.0005
R8316 AVSS.n1965 AVSS.n1962 16.0005
R8317 AVSS.n1962 AVSS.n1961 16.0005
R8318 AVSS.n1961 AVSS.n1958 16.0005
R8319 AVSS.n1958 AVSS.n1887 16.0005
R8320 AVSS.n1974 AVSS.n1887 16.0005
R8321 AVSS.n1785 AVSS.n1783 16.0005
R8322 AVSS.n1783 AVSS.n1780 16.0005
R8323 AVSS.n1780 AVSS.n1779 16.0005
R8324 AVSS.n1779 AVSS.n1776 16.0005
R8325 AVSS.n1776 AVSS.n1775 16.0005
R8326 AVSS.n1775 AVSS.n1772 16.0005
R8327 AVSS.n1772 AVSS.n1751 16.0005
R8328 AVSS.n2559 AVSS.n1751 16.0005
R8329 AVSS.n2554 AVSS.n1787 16.0005
R8330 AVSS.n2554 AVSS.n2553 16.0005
R8331 AVSS.n2553 AVSS.n2552 16.0005
R8332 AVSS.n2552 AVSS.n2549 16.0005
R8333 AVSS.n2549 AVSS.n2548 16.0005
R8334 AVSS.n2548 AVSS.n2545 16.0005
R8335 AVSS.n2545 AVSS.n2544 16.0005
R8336 AVSS.n2544 AVSS.n2541 16.0005
R8337 AVSS.n1822 AVSS.n1819 16.0005
R8338 AVSS.n1819 AVSS.n1818 16.0005
R8339 AVSS.n1818 AVSS.n1815 16.0005
R8340 AVSS.n1815 AVSS.n1814 16.0005
R8341 AVSS.n1814 AVSS.n1811 16.0005
R8342 AVSS.n1811 AVSS.n1810 16.0005
R8343 AVSS.n1810 AVSS.n1807 16.0005
R8344 AVSS.n1807 AVSS.n1806 16.0005
R8345 AVSS.n3342 AVSS.n3340 16.0005
R8346 AVSS.n3340 AVSS.n3337 16.0005
R8347 AVSS.n3337 AVSS.n3336 16.0005
R8348 AVSS.n3336 AVSS.n3333 16.0005
R8349 AVSS.n3333 AVSS.n3332 16.0005
R8350 AVSS.n3329 AVSS.n3328 16.0005
R8351 AVSS.n3328 AVSS.n3304 16.0005
R8352 AVSS.n3359 AVSS.n3357 16.0005
R8353 AVSS.n3357 AVSS.n3356 16.0005
R8354 AVSS.n3356 AVSS.n3354 16.0005
R8355 AVSS.n3354 AVSS.n3351 16.0005
R8356 AVSS.n3351 AVSS.n3350 16.0005
R8357 AVSS.n3350 AVSS.n3347 16.0005
R8358 AVSS.n3347 AVSS.n3346 16.0005
R8359 AVSS.n3346 AVSS.n3344 16.0005
R8360 AVSS.n3363 AVSS.n3360 16.0005
R8361 AVSS.n3364 AVSS.n3363 16.0005
R8362 AVSS.n3367 AVSS.n3364 16.0005
R8363 AVSS.n3368 AVSS.n3367 16.0005
R8364 AVSS.n3371 AVSS.n3368 16.0005
R8365 AVSS.n3372 AVSS.n3371 16.0005
R8366 AVSS.n3375 AVSS.n3372 16.0005
R8367 AVSS.n3376 AVSS.n3375 16.0005
R8368 AVSS.n3388 AVSS.n3387 16.0005
R8369 AVSS.n3387 AVSS.n3386 16.0005
R8370 AVSS.n3386 AVSS.n3384 16.0005
R8371 AVSS.n3384 AVSS.n3381 16.0005
R8372 AVSS.n3381 AVSS.n3380 16.0005
R8373 AVSS.n3380 AVSS.n3377 16.0005
R8374 AVSS.n3377 AVSS.n3305 16.0005
R8375 AVSS.n3393 AVSS.n3305 16.0005
R8376 AVSS.n6038 AVSS.n5935 14.2369
R8377 AVSS.n6029 AVSS.n6004 14.0847
R8378 AVSS.n4149 AVSS.n4136 13.5116
R8379 AVSS.n4080 AVSS.n4079 13.5116
R8380 AVSS.n3869 AVSS.n3868 13.5116
R8381 AVSS.n3509 AVSS.n3508 13.5116
R8382 AVSS.n5392 AVSS.n5301 13.5116
R8383 AVSS.n5193 AVSS.n5102 13.5116
R8384 AVSS.n551 AVSS.n462 13.5116
R8385 AVSS.n1459 AVSS.n1458 13.5116
R8386 AVSS.n1480 AVSS.n1479 13.5116
R8387 AVSS.n4879 AVSS.n4878 13.5116
R8388 AVSS.n4900 AVSS.n4899 13.5116
R8389 AVSS.n2682 AVSS.n2681 13.5116
R8390 AVSS.n1714 AVSS.n1713 13.5116
R8391 AVSS.n1803 AVSS.n1788 13.5116
R8392 AVSS.n2046 AVSS.n2045 13.5116
R8393 AVSS.n2067 AVSS.n2066 13.5116
R8394 AVSS.n2454 AVSS.n2453 13.5116
R8395 AVSS.n1975 AVSS.n1886 13.5116
R8396 AVSS.n2560 AVSS.n2559 13.5116
R8397 AVSS.n3394 AVSS.n3304 13.5116
R8398 AVSS.n3344 AVSS.n3343 13.5116
R8399 AVSS.n113 AVSS 12.9783
R8400 AVSS.n4164 AVSS 12.9783
R8401 AVSS.n4021 AVSS 12.9783
R8402 AVSS.n3810 AVSS 12.9783
R8403 AVSS.n3451 AVSS 12.9783
R8404 AVSS AVSS.n5766 12.9783
R8405 AVSS AVSS.n5494 12.9783
R8406 AVSS AVSS.n5326 12.9783
R8407 AVSS AVSS.n5127 12.9783
R8408 AVSS.n487 AVSS 12.9783
R8409 AVSS.n1454 AVSS 12.9783
R8410 AVSS.n4874 AVSS 12.9783
R8411 AVSS.n3187 AVSS 12.9783
R8412 AVSS.n1263 AVSS 12.9783
R8413 AVSS AVSS.n4563 12.9783
R8414 AVSS.n2741 AVSS 12.9783
R8415 AVSS.n2623 AVSS 12.9783
R8416 AVSS.n1656 AVSS 12.9783
R8417 AVSS.n1799 AVSS 12.9783
R8418 AVSS.n2041 AVSS 12.9783
R8419 AVSS.n804 AVSS 12.9783
R8420 AVSS AVSS.n1014 12.9783
R8421 AVSS AVSS.n2459 12.9783
R8422 AVSS.n1911 AVSS 12.9783
R8423 AVSS.n3329 AVSS 12.9783
R8424 AVSS.n4983 AVSS.n46 12.2888
R8425 AVSS.n4669 AVSS.n50 12.2888
R8426 AVSS.n2191 AVSS.n1595 12.2265
R8427 AVSS.n4723 AVSS.n4722 12.2265
R8428 AVSS.n1196 AVSS.n1195 11.6369
R8429 AVSS.n1195 AVSS.n1166 11.6369
R8430 AVSS.n1189 AVSS.n1166 11.6369
R8431 AVSS.n1189 AVSS.n1188 11.6369
R8432 AVSS.n1188 AVSS.n1187 11.6369
R8433 AVSS.n1187 AVSS.n1184 11.6369
R8434 AVSS.n1184 AVSS.n1183 11.6369
R8435 AVSS.n1183 AVSS.n1180 11.6369
R8436 AVSS.n1180 AVSS.n1179 11.6369
R8437 AVSS.n1179 AVSS.n1176 11.6369
R8438 AVSS.n1176 AVSS.n1175 11.6369
R8439 AVSS.n1300 AVSS.n1164 11.6369
R8440 AVSS.n1301 AVSS.n1300 11.6369
R8441 AVSS.n1302 AVSS.n1301 11.6369
R8442 AVSS.n1302 AVSS.n1162 11.6369
R8443 AVSS.n1308 AVSS.n1162 11.6369
R8444 AVSS.n1309 AVSS.n1308 11.6369
R8445 AVSS.n1310 AVSS.n1309 11.6369
R8446 AVSS.n1310 AVSS.n1160 11.6369
R8447 AVSS.n1315 AVSS.n1160 11.6369
R8448 AVSS.n1316 AVSS.n1315 11.6369
R8449 AVSS.n1316 AVSS.n1158 11.6369
R8450 AVSS.n1323 AVSS.n1322 11.6369
R8451 AVSS.n1324 AVSS.n1323 11.6369
R8452 AVSS.n1324 AVSS.n1154 11.6369
R8453 AVSS.n1331 AVSS.n1154 11.6369
R8454 AVSS.n1332 AVSS.n1331 11.6369
R8455 AVSS.n1333 AVSS.n1332 11.6369
R8456 AVSS.n1338 AVSS.n1152 11.6369
R8457 AVSS.n1339 AVSS.n1338 11.6369
R8458 AVSS.n1341 AVSS.n1339 11.6369
R8459 AVSS.n1341 AVSS.n1340 11.6369
R8460 AVSS.n1366 AVSS.n1365 11.6369
R8461 AVSS.n1365 AVSS.n1364 11.6369
R8462 AVSS.n1364 AVSS.n1361 11.6369
R8463 AVSS.n1361 AVSS.n1360 11.6369
R8464 AVSS.n1360 AVSS.n1357 11.6369
R8465 AVSS.n1357 AVSS.n1356 11.6369
R8466 AVSS.n1356 AVSS.n1353 11.6369
R8467 AVSS.n1353 AVSS.n1352 11.6369
R8468 AVSS.n1352 AVSS.n1349 11.6369
R8469 AVSS.n1349 AVSS.n1348 11.6369
R8470 AVSS.n1348 AVSS.n1148 11.6369
R8471 AVSS.n4624 AVSS.n4623 11.6369
R8472 AVSS.n4630 AVSS.n4623 11.6369
R8473 AVSS.n4631 AVSS.n4630 11.6369
R8474 AVSS.n4632 AVSS.n4631 11.6369
R8475 AVSS.n4632 AVSS.n4621 11.6369
R8476 AVSS.n4638 AVSS.n4621 11.6369
R8477 AVSS.n4639 AVSS.n4638 11.6369
R8478 AVSS.n4640 AVSS.n4639 11.6369
R8479 AVSS.n4640 AVSS.n4619 11.6369
R8480 AVSS.n4619 AVSS.n4617 11.6369
R8481 AVSS.n4647 AVSS.n4617 11.6369
R8482 AVSS.n4980 AVSS.n1069 11.6369
R8483 AVSS.n1072 AVSS.n1069 11.6369
R8484 AVSS.n4973 AVSS.n1072 11.6369
R8485 AVSS.n4973 AVSS.n4972 11.6369
R8486 AVSS.n4972 AVSS.n4971 11.6369
R8487 AVSS.n4971 AVSS.n1074 11.6369
R8488 AVSS.n4966 AVSS.n1074 11.6369
R8489 AVSS.n4966 AVSS.n4965 11.6369
R8490 AVSS.n4965 AVSS.n4964 11.6369
R8491 AVSS.n4964 AVSS.n1077 11.6369
R8492 AVSS.n4959 AVSS.n1077 11.6369
R8493 AVSS.n4958 AVSS.n4957 11.6369
R8494 AVSS.n4957 AVSS.n1080 11.6369
R8495 AVSS.n4952 AVSS.n1080 11.6369
R8496 AVSS.n4952 AVSS.n4951 11.6369
R8497 AVSS.n4951 AVSS.n4950 11.6369
R8498 AVSS.n4950 AVSS.n1084 11.6369
R8499 AVSS.n4945 AVSS.n4944 11.6369
R8500 AVSS.n4944 AVSS.n4943 11.6369
R8501 AVSS.n4943 AVSS.n1087 11.6369
R8502 AVSS.n4938 AVSS.n1087 11.6369
R8503 AVSS.n4666 AVSS.n4664 11.6369
R8504 AVSS.n4664 AVSS.n4661 11.6369
R8505 AVSS.n4661 AVSS.n4660 11.6369
R8506 AVSS.n4660 AVSS.n4657 11.6369
R8507 AVSS.n4657 AVSS.n4656 11.6369
R8508 AVSS.n4656 AVSS.n4653 11.6369
R8509 AVSS.n4653 AVSS.n4652 11.6369
R8510 AVSS.n4652 AVSS.n4649 11.6369
R8511 AVSS.n4649 AVSS.n1090 11.6369
R8512 AVSS.n4936 AVSS.n1090 11.6369
R8513 AVSS.n4937 AVSS.n4936 11.6369
R8514 AVSS.n2114 AVSS.n2088 11.6369
R8515 AVSS.n2120 AVSS.n2088 11.6369
R8516 AVSS.n2121 AVSS.n2120 11.6369
R8517 AVSS.n2122 AVSS.n2121 11.6369
R8518 AVSS.n2122 AVSS.n2086 11.6369
R8519 AVSS.n2128 AVSS.n2086 11.6369
R8520 AVSS.n2129 AVSS.n2128 11.6369
R8521 AVSS.n2130 AVSS.n2129 11.6369
R8522 AVSS.n2130 AVSS.n2084 11.6369
R8523 AVSS.n2084 AVSS.n2082 11.6369
R8524 AVSS.n2137 AVSS.n2082 11.6369
R8525 AVSS.n2113 AVSS.n2112 11.6369
R8526 AVSS.n2112 AVSS.n2090 11.6369
R8527 AVSS.n2091 AVSS.n2090 11.6369
R8528 AVSS.n2105 AVSS.n2091 11.6369
R8529 AVSS.n2105 AVSS.n2104 11.6369
R8530 AVSS.n2104 AVSS.n2103 11.6369
R8531 AVSS.n2103 AVSS.n2093 11.6369
R8532 AVSS.n2098 AVSS.n2093 11.6369
R8533 AVSS.n2098 AVSS.n2097 11.6369
R8534 AVSS.n2097 AVSS.n2069 11.6369
R8535 AVSS.n2188 AVSS.n2070 11.6369
R8536 AVSS.n2181 AVSS.n2072 11.6369
R8537 AVSS.n2181 AVSS.n2180 11.6369
R8538 AVSS.n2180 AVSS.n2179 11.6369
R8539 AVSS.n2179 AVSS.n2075 11.6369
R8540 AVSS.n2174 AVSS.n2075 11.6369
R8541 AVSS.n2174 AVSS.n2173 11.6369
R8542 AVSS.n2172 AVSS.n2078 11.6369
R8543 AVSS.n2167 AVSS.n2078 11.6369
R8544 AVSS.n2167 AVSS.n2166 11.6369
R8545 AVSS.n2166 AVSS.n2165 11.6369
R8546 AVSS.n2140 AVSS.n2138 11.6369
R8547 AVSS.n2141 AVSS.n2140 11.6369
R8548 AVSS.n2144 AVSS.n2141 11.6369
R8549 AVSS.n2145 AVSS.n2144 11.6369
R8550 AVSS.n2148 AVSS.n2145 11.6369
R8551 AVSS.n2149 AVSS.n2148 11.6369
R8552 AVSS.n2152 AVSS.n2149 11.6369
R8553 AVSS.n2153 AVSS.n2152 11.6369
R8554 AVSS.n2156 AVSS.n2153 11.6369
R8555 AVSS.n2157 AVSS.n2156 11.6369
R8556 AVSS.n2161 AVSS.n2160 11.6369
R8557 AVSS.n5570 AVSS.n5276 11.6369
R8558 AVSS.n5576 AVSS.n5276 11.6369
R8559 AVSS.n5577 AVSS.n5576 11.6369
R8560 AVSS.n5578 AVSS.n5577 11.6369
R8561 AVSS.n5578 AVSS.n5272 11.6369
R8562 AVSS.n5584 AVSS.n5272 11.6369
R8563 AVSS.n5585 AVSS.n5584 11.6369
R8564 AVSS.n5586 AVSS.n5585 11.6369
R8565 AVSS.n5586 AVSS.n5268 11.6369
R8566 AVSS.n5592 AVSS.n5268 11.6369
R8567 AVSS.n5593 AVSS.n5592 11.6369
R8568 AVSS.n5614 AVSS.n5593 11.6369
R8569 AVSS.n5613 AVSS.n5612 11.6369
R8570 AVSS.n5612 AVSS.n5609 11.6369
R8571 AVSS.n5609 AVSS.n5608 11.6369
R8572 AVSS.n5608 AVSS.n5605 11.6369
R8573 AVSS.n5605 AVSS.n5604 11.6369
R8574 AVSS.n5604 AVSS.n5601 11.6369
R8575 AVSS.n5600 AVSS.n5597 11.6369
R8576 AVSS.n5597 AVSS.n5596 11.6369
R8577 AVSS.n5596 AVSS.n5594 11.6369
R8578 AVSS.n5594 AVSS.n5258 11.6369
R8579 AVSS.n5871 AVSS.n5870 11.6369
R8580 AVSS.n5870 AVSS.n5869 11.6369
R8581 AVSS.n5869 AVSS.n5866 11.6369
R8582 AVSS.n5866 AVSS.n5865 11.6369
R8583 AVSS.n5865 AVSS.n5862 11.6369
R8584 AVSS.n5862 AVSS.n5861 11.6369
R8585 AVSS.n5861 AVSS.n5858 11.6369
R8586 AVSS.n5858 AVSS.n5857 11.6369
R8587 AVSS.n5857 AVSS.n5854 11.6369
R8588 AVSS.n5854 AVSS.n5853 11.6369
R8589 AVSS.n5853 AVSS.n5850 11.6369
R8590 AVSS.n5850 AVSS.n5849 11.6369
R8591 AVSS.n5569 AVSS.n5568 11.6369
R8592 AVSS.n5568 AVSS.n5448 11.6369
R8593 AVSS.n5562 AVSS.n5448 11.6369
R8594 AVSS.n5562 AVSS.n5561 11.6369
R8595 AVSS.n5561 AVSS.n5560 11.6369
R8596 AVSS.n5560 AVSS.n5557 11.6369
R8597 AVSS.n5557 AVSS.n5556 11.6369
R8598 AVSS.n5556 AVSS.n5553 11.6369
R8599 AVSS.n5553 AVSS.n5552 11.6369
R8600 AVSS.n5552 AVSS.n5549 11.6369
R8601 AVSS.n6277 AVSS.n6276 11.6369
R8602 AVSS.n6276 AVSS.n12 11.6369
R8603 AVSS.n6270 AVSS.n12 11.6369
R8604 AVSS.n6270 AVSS.n6269 11.6369
R8605 AVSS.n6269 AVSS.n6268 11.6369
R8606 AVSS.n6268 AVSS.n17 11.6369
R8607 AVSS.n5286 AVSS.n17 11.6369
R8608 AVSS.n5287 AVSS.n5286 11.6369
R8609 AVSS.n5287 AVSS.n5282 11.6369
R8610 AVSS.n5293 AVSS.n5282 11.6369
R8611 AVSS.n5294 AVSS.n5293 11.6369
R8612 AVSS.n5443 AVSS.n5294 11.6369
R8613 AVSS.n5442 AVSS.n5441 11.6369
R8614 AVSS.n5441 AVSS.n5295 11.6369
R8615 AVSS.n5435 AVSS.n5295 11.6369
R8616 AVSS.n5435 AVSS.n5434 11.6369
R8617 AVSS.n5434 AVSS.n5433 11.6369
R8618 AVSS.n5433 AVSS.n5297 11.6369
R8619 AVSS.n5427 AVSS.n5426 11.6369
R8620 AVSS.n5426 AVSS.n5425 11.6369
R8621 AVSS.n5425 AVSS.n5299 11.6369
R8622 AVSS.n5397 AVSS.n3 11.6369
R8623 AVSS.n5398 AVSS.n5397 11.6369
R8624 AVSS.n5401 AVSS.n5398 11.6369
R8625 AVSS.n5402 AVSS.n5401 11.6369
R8626 AVSS.n5405 AVSS.n5402 11.6369
R8627 AVSS.n5406 AVSS.n5405 11.6369
R8628 AVSS.n5409 AVSS.n5406 11.6369
R8629 AVSS.n5410 AVSS.n5409 11.6369
R8630 AVSS.n5413 AVSS.n5410 11.6369
R8631 AVSS.n5414 AVSS.n5413 11.6369
R8632 AVSS.n5417 AVSS.n5414 11.6369
R8633 AVSS.n5418 AVSS.n5417 11.6369
R8634 AVSS.n6278 AVSS.n10 11.6369
R8635 AVSS.n6284 AVSS.n10 11.6369
R8636 AVSS.n6285 AVSS.n6284 11.6369
R8637 AVSS.n6286 AVSS.n6285 11.6369
R8638 AVSS.n6286 AVSS.n8 11.6369
R8639 AVSS.n6292 AVSS.n8 11.6369
R8640 AVSS.n6293 AVSS.n6292 11.6369
R8641 AVSS.n6294 AVSS.n6293 11.6369
R8642 AVSS.n6294 AVSS.n6 11.6369
R8643 AVSS.n6 AVSS.n2 11.6369
R8644 AVSS.n5076 AVSS.n5075 11.6369
R8645 AVSS.n5075 AVSS.n429 11.6369
R8646 AVSS.n5069 AVSS.n429 11.6369
R8647 AVSS.n5069 AVSS.n5068 11.6369
R8648 AVSS.n5068 AVSS.n5067 11.6369
R8649 AVSS.n5067 AVSS.n434 11.6369
R8650 AVSS.n445 AVSS.n434 11.6369
R8651 AVSS.n445 AVSS.n444 11.6369
R8652 AVSS.n444 AVSS.n443 11.6369
R8653 AVSS.n443 AVSS.n438 11.6369
R8654 AVSS.n438 AVSS.n419 11.6369
R8655 AVSS.n5217 AVSS.n419 11.6369
R8656 AVSS.n5216 AVSS.n5215 11.6369
R8657 AVSS.n5215 AVSS.n5212 11.6369
R8658 AVSS.n5212 AVSS.n5211 11.6369
R8659 AVSS.n5211 AVSS.n5208 11.6369
R8660 AVSS.n5208 AVSS.n5207 11.6369
R8661 AVSS.n5207 AVSS.n5204 11.6369
R8662 AVSS.n5203 AVSS.n5200 11.6369
R8663 AVSS.n5200 AVSS.n5199 11.6369
R8664 AVSS.n5199 AVSS.n5197 11.6369
R8665 AVSS.n5247 AVSS.n5246 11.6369
R8666 AVSS.n5246 AVSS.n5245 11.6369
R8667 AVSS.n5245 AVSS.n5242 11.6369
R8668 AVSS.n5242 AVSS.n5241 11.6369
R8669 AVSS.n5241 AVSS.n5238 11.6369
R8670 AVSS.n5238 AVSS.n5237 11.6369
R8671 AVSS.n5237 AVSS.n5234 11.6369
R8672 AVSS.n5234 AVSS.n5233 11.6369
R8673 AVSS.n5233 AVSS.n5230 11.6369
R8674 AVSS.n5230 AVSS.n5229 11.6369
R8675 AVSS.n5229 AVSS.n5226 11.6369
R8676 AVSS.n5226 AVSS.n5225 11.6369
R8677 AVSS.n5092 AVSS.n5091 11.6369
R8678 AVSS.n5091 AVSS.n5090 11.6369
R8679 AVSS.n5090 AVSS.n5088 11.6369
R8680 AVSS.n5088 AVSS.n5085 11.6369
R8681 AVSS.n5085 AVSS.n5084 11.6369
R8682 AVSS.n5084 AVSS.n5081 11.6369
R8683 AVSS.n5081 AVSS.n5080 11.6369
R8684 AVSS.n5080 AVSS.n5077 11.6369
R8685 AVSS.n5077 AVSS.n421 11.6369
R8686 AVSS.n5098 AVSS.n421 11.6369
R8687 AVSS.n5923 AVSS.n5922 11.6369
R8688 AVSS.n5922 AVSS.n5921 11.6369
R8689 AVSS.n5921 AVSS.n303 11.6369
R8690 AVSS.n5915 AVSS.n303 11.6369
R8691 AVSS.n5915 AVSS.n5914 11.6369
R8692 AVSS.n5914 AVSS.n5913 11.6369
R8693 AVSS.n5913 AVSS.n307 11.6369
R8694 AVSS.n5907 AVSS.n307 11.6369
R8695 AVSS.n5907 AVSS.n5906 11.6369
R8696 AVSS.n5906 AVSS.n5905 11.6369
R8697 AVSS.n5905 AVSS.n311 11.6369
R8698 AVSS.n5899 AVSS.n311 11.6369
R8699 AVSS.n358 AVSS.n302 11.6369
R8700 AVSS.n359 AVSS.n358 11.6369
R8701 AVSS.n360 AVSS.n359 11.6369
R8702 AVSS.n360 AVSS.n352 11.6369
R8703 AVSS.n366 AVSS.n352 11.6369
R8704 AVSS.n367 AVSS.n366 11.6369
R8705 AVSS.n368 AVSS.n367 11.6369
R8706 AVSS.n368 AVSS.n348 11.6369
R8707 AVSS.n374 AVSS.n348 11.6369
R8708 AVSS.n375 AVSS.n374 11.6369
R8709 AVSS.n396 AVSS.n375 11.6369
R8710 AVSS.n395 AVSS.n394 11.6369
R8711 AVSS.n394 AVSS.n392 11.6369
R8712 AVSS.n392 AVSS.n389 11.6369
R8713 AVSS.n389 AVSS.n388 11.6369
R8714 AVSS.n388 AVSS.n385 11.6369
R8715 AVSS.n385 AVSS.n384 11.6369
R8716 AVSS.n384 AVSS.n381 11.6369
R8717 AVSS.n381 AVSS.n380 11.6369
R8718 AVSS.n380 AVSS.n377 11.6369
R8719 AVSS.n377 AVSS.n376 11.6369
R8720 AVSS.n5877 AVSS.n5876 11.6369
R8721 AVSS.n5898 AVSS.n5897 11.6369
R8722 AVSS.n5897 AVSS.n315 11.6369
R8723 AVSS.n5892 AVSS.n315 11.6369
R8724 AVSS.n5892 AVSS.n5891 11.6369
R8725 AVSS.n5891 AVSS.n5890 11.6369
R8726 AVSS.n5890 AVSS.n319 11.6369
R8727 AVSS.n5885 AVSS.n5884 11.6369
R8728 AVSS.n5884 AVSS.n5883 11.6369
R8729 AVSS.n5883 AVSS.n322 11.6369
R8730 AVSS.n5840 AVSS.n5839 11.6369
R8731 AVSS.n5839 AVSS.n5838 11.6369
R8732 AVSS.n5838 AVSS.n5836 11.6369
R8733 AVSS.n5836 AVSS.n5833 11.6369
R8734 AVSS.n5833 AVSS.n5832 11.6369
R8735 AVSS.n5832 AVSS.n5829 11.6369
R8736 AVSS.n5829 AVSS.n5828 11.6369
R8737 AVSS.n5828 AVSS.n5825 11.6369
R8738 AVSS.n5825 AVSS.n5824 11.6369
R8739 AVSS.n5824 AVSS.n5821 11.6369
R8740 AVSS.n5652 AVSS.n5625 11.6369
R8741 AVSS.n5654 AVSS.n5652 11.6369
R8742 AVSS.n5654 AVSS.n5653 11.6369
R8743 AVSS.n5653 AVSS.n5648 11.6369
R8744 AVSS.n5661 AVSS.n5648 11.6369
R8745 AVSS.n5662 AVSS.n5661 11.6369
R8746 AVSS.n5663 AVSS.n5662 11.6369
R8747 AVSS.n5663 AVSS.n5645 11.6369
R8748 AVSS.n5669 AVSS.n5645 11.6369
R8749 AVSS.n5670 AVSS.n5669 11.6369
R8750 AVSS.n5671 AVSS.n5670 11.6369
R8751 AVSS.n5671 AVSS.n5641 11.6369
R8752 AVSS.n5678 AVSS.n5677 11.6369
R8753 AVSS.n5679 AVSS.n5678 11.6369
R8754 AVSS.n5679 AVSS.n5637 11.6369
R8755 AVSS.n5686 AVSS.n5637 11.6369
R8756 AVSS.n5687 AVSS.n5686 11.6369
R8757 AVSS.n5688 AVSS.n5687 11.6369
R8758 AVSS.n5694 AVSS.n5634 11.6369
R8759 AVSS.n5695 AVSS.n5694 11.6369
R8760 AVSS.n5697 AVSS.n5695 11.6369
R8761 AVSS.n5697 AVSS.n5696 11.6369
R8762 AVSS.n5724 AVSS.n5721 11.6369
R8763 AVSS.n5721 AVSS.n5720 11.6369
R8764 AVSS.n5720 AVSS.n5717 11.6369
R8765 AVSS.n5717 AVSS.n5716 11.6369
R8766 AVSS.n5716 AVSS.n5713 11.6369
R8767 AVSS.n5713 AVSS.n5712 11.6369
R8768 AVSS.n5712 AVSS.n5709 11.6369
R8769 AVSS.n5709 AVSS.n5708 11.6369
R8770 AVSS.n5708 AVSS.n5705 11.6369
R8771 AVSS.n5705 AVSS.n5704 11.6369
R8772 AVSS.n5704 AVSS.n5630 11.6369
R8773 AVSS.n838 AVSS.n835 11.6369
R8774 AVSS.n839 AVSS.n838 11.6369
R8775 AVSS.n842 AVSS.n839 11.6369
R8776 AVSS.n843 AVSS.n842 11.6369
R8777 AVSS.n846 AVSS.n843 11.6369
R8778 AVSS.n847 AVSS.n846 11.6369
R8779 AVSS.n850 AVSS.n847 11.6369
R8780 AVSS.n851 AVSS.n850 11.6369
R8781 AVSS.n854 AVSS.n851 11.6369
R8782 AVSS.n855 AVSS.n854 11.6369
R8783 AVSS.n856 AVSS.n855 11.6369
R8784 AVSS.n862 AVSS.n680 11.6369
R8785 AVSS.n863 AVSS.n862 11.6369
R8786 AVSS.n865 AVSS.n863 11.6369
R8787 AVSS.n865 AVSS.n864 11.6369
R8788 AVSS.n864 AVSS.n676 11.6369
R8789 AVSS.n873 AVSS.n676 11.6369
R8790 AVSS.n875 AVSS.n874 11.6369
R8791 AVSS.n875 AVSS.n672 11.6369
R8792 AVSS.n881 AVSS.n672 11.6369
R8793 AVSS.n882 AVSS.n881 11.6369
R8794 AVSS.n736 AVSS.n733 11.6369
R8795 AVSS.n733 AVSS.n732 11.6369
R8796 AVSS.n732 AVSS.n729 11.6369
R8797 AVSS.n729 AVSS.n728 11.6369
R8798 AVSS.n728 AVSS.n725 11.6369
R8799 AVSS.n725 AVSS.n724 11.6369
R8800 AVSS.n724 AVSS.n721 11.6369
R8801 AVSS.n721 AVSS.n720 11.6369
R8802 AVSS.n720 AVSS.n717 11.6369
R8803 AVSS.n717 AVSS.n671 11.6369
R8804 AVSS.n883 AVSS.n671 11.6369
R8805 AVSS.n694 AVSS.n693 11.6369
R8806 AVSS.n695 AVSS.n694 11.6369
R8807 AVSS.n695 AVSS.n688 11.6369
R8808 AVSS.n701 AVSS.n688 11.6369
R8809 AVSS.n702 AVSS.n701 11.6369
R8810 AVSS.n703 AVSS.n702 11.6369
R8811 AVSS.n703 AVSS.n686 11.6369
R8812 AVSS.n709 AVSS.n686 11.6369
R8813 AVSS.n710 AVSS.n709 11.6369
R8814 AVSS.n711 AVSS.n710 11.6369
R8815 AVSS.n711 AVSS.n684 11.6369
R8816 AVSS.n2277 AVSS.n2276 11.6369
R8817 AVSS.n2276 AVSS.n2274 11.6369
R8818 AVSS.n2274 AVSS.n2271 11.6369
R8819 AVSS.n2271 AVSS.n2270 11.6369
R8820 AVSS.n2270 AVSS.n2267 11.6369
R8821 AVSS.n2267 AVSS.n2266 11.6369
R8822 AVSS.n2266 AVSS.n2263 11.6369
R8823 AVSS.n2263 AVSS.n2262 11.6369
R8824 AVSS.n2262 AVSS.n2259 11.6369
R8825 AVSS.n2259 AVSS.n2258 11.6369
R8826 AVSS.n2258 AVSS.n2255 11.6369
R8827 AVSS.n2255 AVSS.n2254 11.6369
R8828 AVSS.n2249 AVSS.n2201 11.6369
R8829 AVSS.n2249 AVSS.n2248 11.6369
R8830 AVSS.n2248 AVSS.n2247 11.6369
R8831 AVSS.n2247 AVSS.n2203 11.6369
R8832 AVSS.n2242 AVSS.n2203 11.6369
R8833 AVSS.n2242 AVSS.n2241 11.6369
R8834 AVSS.n2240 AVSS.n2206 11.6369
R8835 AVSS.n2235 AVSS.n2206 11.6369
R8836 AVSS.n2235 AVSS.n2234 11.6369
R8837 AVSS.n2234 AVSS.n2233 11.6369
R8838 AVSS.n2209 AVSS.n974 11.6369
R8839 AVSS.n2212 AVSS.n2209 11.6369
R8840 AVSS.n2213 AVSS.n2212 11.6369
R8841 AVSS.n2216 AVSS.n2213 11.6369
R8842 AVSS.n2217 AVSS.n2216 11.6369
R8843 AVSS.n2220 AVSS.n2217 11.6369
R8844 AVSS.n2221 AVSS.n2220 11.6369
R8845 AVSS.n2224 AVSS.n2221 11.6369
R8846 AVSS.n2225 AVSS.n2224 11.6369
R8847 AVSS.n2228 AVSS.n2225 11.6369
R8848 AVSS.n2229 AVSS.n2228 11.6369
R8849 AVSS.n2278 AVSS.n2200 11.6369
R8850 AVSS.n2284 AVSS.n2200 11.6369
R8851 AVSS.n2285 AVSS.n2284 11.6369
R8852 AVSS.n2286 AVSS.n2285 11.6369
R8853 AVSS.n2286 AVSS.n2198 11.6369
R8854 AVSS.n2292 AVSS.n2198 11.6369
R8855 AVSS.n2293 AVSS.n2292 11.6369
R8856 AVSS.n2294 AVSS.n2293 11.6369
R8857 AVSS.n2294 AVSS.n2196 11.6369
R8858 AVSS.n2300 AVSS.n2196 11.6369
R8859 AVSS.n2366 AVSS.n2364 11.6369
R8860 AVSS.n2367 AVSS.n2366 11.6369
R8861 AVSS.n2370 AVSS.n2367 11.6369
R8862 AVSS.n2371 AVSS.n2370 11.6369
R8863 AVSS.n2374 AVSS.n2371 11.6369
R8864 AVSS.n2375 AVSS.n2374 11.6369
R8865 AVSS.n2378 AVSS.n2375 11.6369
R8866 AVSS.n2379 AVSS.n2378 11.6369
R8867 AVSS.n2382 AVSS.n2379 11.6369
R8868 AVSS.n2383 AVSS.n2382 11.6369
R8869 AVSS.n2386 AVSS.n2383 11.6369
R8870 AVSS.n2387 AVSS.n2386 11.6369
R8871 AVSS.n2392 AVSS.n2391 11.6369
R8872 AVSS.n2393 AVSS.n2392 11.6369
R8873 AVSS.n2393 AVSS.n2308 11.6369
R8874 AVSS.n2399 AVSS.n2308 11.6369
R8875 AVSS.n2400 AVSS.n2399 11.6369
R8876 AVSS.n2401 AVSS.n2400 11.6369
R8877 AVSS.n2406 AVSS.n2306 11.6369
R8878 AVSS.n2407 AVSS.n2406 11.6369
R8879 AVSS.n2407 AVSS.n2303 11.6369
R8880 AVSS.n2338 AVSS.n2337 11.6369
R8881 AVSS.n2337 AVSS.n2335 11.6369
R8882 AVSS.n2335 AVSS.n2332 11.6369
R8883 AVSS.n2332 AVSS.n2331 11.6369
R8884 AVSS.n2331 AVSS.n2328 11.6369
R8885 AVSS.n2328 AVSS.n2327 11.6369
R8886 AVSS.n2327 AVSS.n2324 11.6369
R8887 AVSS.n2324 AVSS.n2323 11.6369
R8888 AVSS.n2323 AVSS.n2320 11.6369
R8889 AVSS.n2320 AVSS.n2319 11.6369
R8890 AVSS.n2319 AVSS.n2316 11.6369
R8891 AVSS.n2316 AVSS.n2304 11.6369
R8892 AVSS.n2363 AVSS.n2310 11.6369
R8893 AVSS.n2358 AVSS.n2310 11.6369
R8894 AVSS.n2358 AVSS.n2357 11.6369
R8895 AVSS.n2357 AVSS.n2312 11.6369
R8896 AVSS.n2352 AVSS.n2312 11.6369
R8897 AVSS.n2352 AVSS.n2351 11.6369
R8898 AVSS.n2351 AVSS.n2350 11.6369
R8899 AVSS.n2350 AVSS.n2314 11.6369
R8900 AVSS.n2344 AVSS.n2314 11.6369
R8901 AVSS.n2344 AVSS.n2343 11.6369
R8902 AVSS.n1541 AVSS.n1539 11.6369
R8903 AVSS.n1542 AVSS.n1541 11.6369
R8904 AVSS.n1545 AVSS.n1542 11.6369
R8905 AVSS.n1546 AVSS.n1545 11.6369
R8906 AVSS.n1549 AVSS.n1546 11.6369
R8907 AVSS.n1550 AVSS.n1549 11.6369
R8908 AVSS.n1553 AVSS.n1550 11.6369
R8909 AVSS.n1554 AVSS.n1553 11.6369
R8910 AVSS.n1557 AVSS.n1554 11.6369
R8911 AVSS.n1558 AVSS.n1557 11.6369
R8912 AVSS.n1562 AVSS.n1561 11.6369
R8913 AVSS.n1538 AVSS.n1484 11.6369
R8914 AVSS.n1532 AVSS.n1484 11.6369
R8915 AVSS.n1532 AVSS.n1531 11.6369
R8916 AVSS.n1531 AVSS.n1530 11.6369
R8917 AVSS.n1530 AVSS.n1488 11.6369
R8918 AVSS.n1490 AVSS.n1488 11.6369
R8919 AVSS.n1493 AVSS.n1490 11.6369
R8920 AVSS.n1520 AVSS.n1493 11.6369
R8921 AVSS.n1520 AVSS.n1519 11.6369
R8922 AVSS.n1519 AVSS.n1518 11.6369
R8923 AVSS.n1518 AVSS.n1513 11.6369
R8924 AVSS.n1512 AVSS.n1511 11.6369
R8925 AVSS.n1511 AVSS.n1509 11.6369
R8926 AVSS.n1509 AVSS.n1506 11.6369
R8927 AVSS.n1506 AVSS.n1505 11.6369
R8928 AVSS.n1505 AVSS.n1502 11.6369
R8929 AVSS.n1502 AVSS.n1501 11.6369
R8930 AVSS.n1501 AVSS.n1498 11.6369
R8931 AVSS.n1498 AVSS.n1497 11.6369
R8932 AVSS.n1497 AVSS.n1494 11.6369
R8933 AVSS.n1494 AVSS.n1383 11.6369
R8934 AVSS.n1592 AVSS.n1589 11.6369
R8935 AVSS.n1567 AVSS.n1566 11.6369
R8936 AVSS.n1568 AVSS.n1567 11.6369
R8937 AVSS.n1568 AVSS.n1388 11.6369
R8938 AVSS.n1574 AVSS.n1388 11.6369
R8939 AVSS.n1575 AVSS.n1574 11.6369
R8940 AVSS.n1576 AVSS.n1575 11.6369
R8941 AVSS.n1582 AVSS.n1386 11.6369
R8942 AVSS.n1583 AVSS.n1582 11.6369
R8943 AVSS.n1584 AVSS.n1583 11.6369
R8944 AVSS.n1584 AVSS.n1384 11.6369
R8945 AVSS.n920 AVSS.n919 11.6369
R8946 AVSS.n919 AVSS.n916 11.6369
R8947 AVSS.n916 AVSS.n915 11.6369
R8948 AVSS.n915 AVSS.n912 11.6369
R8949 AVSS.n912 AVSS.n911 11.6369
R8950 AVSS.n911 AVSS.n908 11.6369
R8951 AVSS.n908 AVSS.n907 11.6369
R8952 AVSS.n907 AVSS.n904 11.6369
R8953 AVSS.n904 AVSS.n903 11.6369
R8954 AVSS.n903 AVSS.n900 11.6369
R8955 AVSS.n900 AVSS.n635 11.6369
R8956 AVSS.n5014 AVSS.n635 11.6369
R8957 AVSS.n921 AVSS.n898 11.6369
R8958 AVSS.n927 AVSS.n898 11.6369
R8959 AVSS.n928 AVSS.n927 11.6369
R8960 AVSS.n929 AVSS.n928 11.6369
R8961 AVSS.n929 AVSS.n896 11.6369
R8962 AVSS.n935 AVSS.n896 11.6369
R8963 AVSS.n936 AVSS.n935 11.6369
R8964 AVSS.n937 AVSS.n936 11.6369
R8965 AVSS.n937 AVSS.n894 11.6369
R8966 AVSS.n943 AVSS.n894 11.6369
R8967 AVSS.n944 AVSS.n943 11.6369
R8968 AVSS.n963 AVSS.n962 11.6369
R8969 AVSS.n962 AVSS.n961 11.6369
R8970 AVSS.n961 AVSS.n958 11.6369
R8971 AVSS.n958 AVSS.n957 11.6369
R8972 AVSS.n957 AVSS.n954 11.6369
R8973 AVSS.n954 AVSS.n953 11.6369
R8974 AVSS.n953 AVSS.n950 11.6369
R8975 AVSS.n950 AVSS.n949 11.6369
R8976 AVSS.n949 AVSS.n946 11.6369
R8977 AVSS.n946 AVSS.n945 11.6369
R8978 AVSS.n4992 AVSS.n4991 11.6369
R8979 AVSS.n5013 AVSS.n5012 11.6369
R8980 AVSS.n5012 AVSS.n636 11.6369
R8981 AVSS.n5007 AVSS.n636 11.6369
R8982 AVSS.n5007 AVSS.n5006 11.6369
R8983 AVSS.n5006 AVSS.n5005 11.6369
R8984 AVSS.n5005 AVSS.n639 11.6369
R8985 AVSS.n5000 AVSS.n4999 11.6369
R8986 AVSS.n4999 AVSS.n4998 11.6369
R8987 AVSS.n4998 AVSS.n642 11.6369
R8988 AVSS.n3224 AVSS.n3090 11.6369
R8989 AVSS.n3225 AVSS.n3224 11.6369
R8990 AVSS.n3226 AVSS.n3225 11.6369
R8991 AVSS.n3226 AVSS.n3088 11.6369
R8992 AVSS.n3232 AVSS.n3088 11.6369
R8993 AVSS.n3233 AVSS.n3232 11.6369
R8994 AVSS.n3234 AVSS.n3233 11.6369
R8995 AVSS.n3234 AVSS.n3086 11.6369
R8996 AVSS.n3239 AVSS.n3086 11.6369
R8997 AVSS.n3240 AVSS.n3239 11.6369
R8998 AVSS.n3240 AVSS.n3084 11.6369
R8999 AVSS.n3247 AVSS.n3246 11.6369
R9000 AVSS.n3248 AVSS.n3247 11.6369
R9001 AVSS.n3248 AVSS.n3080 11.6369
R9002 AVSS.n3255 AVSS.n3080 11.6369
R9003 AVSS.n3256 AVSS.n3255 11.6369
R9004 AVSS.n3257 AVSS.n3256 11.6369
R9005 AVSS.n3263 AVSS.n3077 11.6369
R9006 AVSS.n3264 AVSS.n3263 11.6369
R9007 AVSS.n3266 AVSS.n3264 11.6369
R9008 AVSS.n3266 AVSS.n3265 11.6369
R9009 AVSS.n3291 AVSS.n3290 11.6369
R9010 AVSS.n3290 AVSS.n3289 11.6369
R9011 AVSS.n3289 AVSS.n3286 11.6369
R9012 AVSS.n3286 AVSS.n3285 11.6369
R9013 AVSS.n3285 AVSS.n3282 11.6369
R9014 AVSS.n3282 AVSS.n3281 11.6369
R9015 AVSS.n3281 AVSS.n3278 11.6369
R9016 AVSS.n3278 AVSS.n3277 11.6369
R9017 AVSS.n3277 AVSS.n3274 11.6369
R9018 AVSS.n3274 AVSS.n3273 11.6369
R9019 AVSS.n3273 AVSS.n3073 11.6369
R9020 AVSS.n3121 AVSS.n3120 11.6369
R9021 AVSS.n3120 AVSS.n3092 11.6369
R9022 AVSS.n3114 AVSS.n3092 11.6369
R9023 AVSS.n3114 AVSS.n3113 11.6369
R9024 AVSS.n3113 AVSS.n3112 11.6369
R9025 AVSS.n3112 AVSS.n3094 11.6369
R9026 AVSS.n3106 AVSS.n3094 11.6369
R9027 AVSS.n3106 AVSS.n3105 11.6369
R9028 AVSS.n3105 AVSS.n3104 11.6369
R9029 AVSS.n3104 AVSS.n3096 11.6369
R9030 AVSS.n3098 AVSS.n3096 11.6369
R9031 AVSS.n4523 AVSS.n4522 11.6369
R9032 AVSS.n4522 AVSS.n2781 11.6369
R9033 AVSS.n4517 AVSS.n2781 11.6369
R9034 AVSS.n4517 AVSS.n4516 11.6369
R9035 AVSS.n4516 AVSS.n4515 11.6369
R9036 AVSS.n4515 AVSS.n2784 11.6369
R9037 AVSS.n4510 AVSS.n2784 11.6369
R9038 AVSS.n4510 AVSS.n4509 11.6369
R9039 AVSS.n4509 AVSS.n4508 11.6369
R9040 AVSS.n4508 AVSS.n2787 11.6369
R9041 AVSS.n4503 AVSS.n2787 11.6369
R9042 AVSS.n4502 AVSS.n4501 11.6369
R9043 AVSS.n4501 AVSS.n2790 11.6369
R9044 AVSS.n2882 AVSS.n2790 11.6369
R9045 AVSS.n2885 AVSS.n2882 11.6369
R9046 AVSS.n2886 AVSS.n2885 11.6369
R9047 AVSS.n2889 AVSS.n2886 11.6369
R9048 AVSS.n2893 AVSS.n2890 11.6369
R9049 AVSS.n2894 AVSS.n2893 11.6369
R9050 AVSS.n2897 AVSS.n2894 11.6369
R9051 AVSS.n2898 AVSS.n2897 11.6369
R9052 AVSS.n2862 AVSS.n2860 11.6369
R9053 AVSS.n2863 AVSS.n2862 11.6369
R9054 AVSS.n2866 AVSS.n2863 11.6369
R9055 AVSS.n2867 AVSS.n2866 11.6369
R9056 AVSS.n2870 AVSS.n2867 11.6369
R9057 AVSS.n2871 AVSS.n2870 11.6369
R9058 AVSS.n2874 AVSS.n2871 11.6369
R9059 AVSS.n2875 AVSS.n2874 11.6369
R9060 AVSS.n2878 AVSS.n2875 11.6369
R9061 AVSS.n2880 AVSS.n2878 11.6369
R9062 AVSS.n2881 AVSS.n2880 11.6369
R9063 AVSS.n2899 AVSS.n2881 11.6369
R9064 AVSS.n4677 AVSS.n2777 11.6369
R9065 AVSS.n2843 AVSS.n2777 11.6369
R9066 AVSS.n2844 AVSS.n2843 11.6369
R9067 AVSS.n2844 AVSS.n2840 11.6369
R9068 AVSS.n2850 AVSS.n2840 11.6369
R9069 AVSS.n2851 AVSS.n2850 11.6369
R9070 AVSS.n2852 AVSS.n2851 11.6369
R9071 AVSS.n2852 AVSS.n2838 11.6369
R9072 AVSS.n2838 AVSS.n2837 11.6369
R9073 AVSS.n2859 AVSS.n2837 11.6369
R9074 AVSS.n4704 AVSS.n4703 11.6369
R9075 AVSS.n4703 AVSS.n4702 11.6369
R9076 AVSS.n4702 AVSS.n1728 11.6369
R9077 AVSS.n4697 AVSS.n1728 11.6369
R9078 AVSS.n4697 AVSS.n4696 11.6369
R9079 AVSS.n4696 AVSS.n4695 11.6369
R9080 AVSS.n4695 AVSS.n1731 11.6369
R9081 AVSS.n4690 AVSS.n1731 11.6369
R9082 AVSS.n4690 AVSS.n4689 11.6369
R9083 AVSS.n4689 AVSS.n4688 11.6369
R9084 AVSS.n4688 AVSS.n1734 11.6369
R9085 AVSS.n4683 AVSS.n1734 11.6369
R9086 AVSS.n3020 AVSS.n1737 11.6369
R9087 AVSS.n3020 AVSS.n3017 11.6369
R9088 AVSS.n3026 AVSS.n3017 11.6369
R9089 AVSS.n3027 AVSS.n3026 11.6369
R9090 AVSS.n3028 AVSS.n3027 11.6369
R9091 AVSS.n3034 AVSS.n3015 11.6369
R9092 AVSS.n3035 AVSS.n3034 11.6369
R9093 AVSS.n3036 AVSS.n3035 11.6369
R9094 AVSS.n3036 AVSS.n3013 11.6369
R9095 AVSS.n3063 AVSS.n3062 11.6369
R9096 AVSS.n3062 AVSS.n3061 11.6369
R9097 AVSS.n3061 AVSS.n3058 11.6369
R9098 AVSS.n3058 AVSS.n3057 11.6369
R9099 AVSS.n3057 AVSS.n3054 11.6369
R9100 AVSS.n3054 AVSS.n3053 11.6369
R9101 AVSS.n3053 AVSS.n3050 11.6369
R9102 AVSS.n3050 AVSS.n3049 11.6369
R9103 AVSS.n3049 AVSS.n3046 11.6369
R9104 AVSS.n3046 AVSS.n3045 11.6369
R9105 AVSS.n3045 AVSS.n3042 11.6369
R9106 AVSS.n3042 AVSS.n3041 11.6369
R9107 AVSS.n4709 AVSS.n1724 11.6369
R9108 AVSS.n2996 AVSS.n1724 11.6369
R9109 AVSS.n2997 AVSS.n2996 11.6369
R9110 AVSS.n2997 AVSS.n2993 11.6369
R9111 AVSS.n3003 AVSS.n2993 11.6369
R9112 AVSS.n3004 AVSS.n3003 11.6369
R9113 AVSS.n3005 AVSS.n3004 11.6369
R9114 AVSS.n3005 AVSS.n2991 11.6369
R9115 AVSS.n3011 AVSS.n2991 11.6369
R9116 AVSS.n3012 AVSS.n3011 11.6369
R9117 AVSS.n2811 AVSS.n1721 11.6369
R9118 AVSS.n2812 AVSS.n2811 11.6369
R9119 AVSS.n2815 AVSS.n2812 11.6369
R9120 AVSS.n2816 AVSS.n2815 11.6369
R9121 AVSS.n2819 AVSS.n2816 11.6369
R9122 AVSS.n2823 AVSS.n2820 11.6369
R9123 AVSS.n2825 AVSS.n2823 11.6369
R9124 AVSS.n2826 AVSS.n2825 11.6369
R9125 AVSS.n4473 AVSS.n2826 11.6369
R9126 AVSS.n2965 AVSS.n2963 11.6369
R9127 AVSS.n2966 AVSS.n2965 11.6369
R9128 AVSS.n2969 AVSS.n2966 11.6369
R9129 AVSS.n2970 AVSS.n2969 11.6369
R9130 AVSS.n2973 AVSS.n2970 11.6369
R9131 AVSS.n2974 AVSS.n2973 11.6369
R9132 AVSS.n2977 AVSS.n2974 11.6369
R9133 AVSS.n2978 AVSS.n2977 11.6369
R9134 AVSS.n2979 AVSS.n2978 11.6369
R9135 AVSS.n2979 AVSS.n2827 11.6369
R9136 AVSS.n4471 AVSS.n2827 11.6369
R9137 AVSS.n4472 AVSS.n4471 11.6369
R9138 AVSS.n2942 AVSS.n2941 11.6369
R9139 AVSS.n2943 AVSS.n2942 11.6369
R9140 AVSS.n2943 AVSS.n2912 11.6369
R9141 AVSS.n2949 AVSS.n2912 11.6369
R9142 AVSS.n2950 AVSS.n2949 11.6369
R9143 AVSS.n2951 AVSS.n2950 11.6369
R9144 AVSS.n2951 AVSS.n2910 11.6369
R9145 AVSS.n2956 AVSS.n2910 11.6369
R9146 AVSS.n2957 AVSS.n2956 11.6369
R9147 AVSS.n2957 AVSS.n2908 11.6369
R9148 AVSS.n2962 AVSS.n2908 11.6369
R9149 AVSS.n2915 AVSS.n2914 11.6369
R9150 AVSS.n2934 AVSS.n2915 11.6369
R9151 AVSS.n2934 AVSS.n2933 11.6369
R9152 AVSS.n2933 AVSS.n2932 11.6369
R9153 AVSS.n2932 AVSS.n2917 11.6369
R9154 AVSS.n2927 AVSS.n2917 11.6369
R9155 AVSS.n2927 AVSS.n2926 11.6369
R9156 AVSS.n2926 AVSS.n2925 11.6369
R9157 AVSS.n2925 AVSS.n2920 11.6369
R9158 AVSS.n2920 AVSS.n1716 11.6369
R9159 AVSS.n4719 AVSS.n1717 11.6369
R9160 AVSS.n4757 AVSS.n4756 11.6369
R9161 AVSS.n4756 AVSS.n4755 11.6369
R9162 AVSS.n4755 AVSS.n4735 11.6369
R9163 AVSS.n4750 AVSS.n4735 11.6369
R9164 AVSS.n4750 AVSS.n4749 11.6369
R9165 AVSS.n4749 AVSS.n4748 11.6369
R9166 AVSS.n4748 AVSS.n4738 11.6369
R9167 AVSS.n4743 AVSS.n4738 11.6369
R9168 AVSS.n4743 AVSS.n4742 11.6369
R9169 AVSS.n4742 AVSS.n1381 11.6369
R9170 AVSS.n4904 AVSS.n1379 11.6369
R9171 AVSS.n4763 AVSS.n4733 11.6369
R9172 AVSS.n4764 AVSS.n4763 11.6369
R9173 AVSS.n4766 AVSS.n4764 11.6369
R9174 AVSS.n4766 AVSS.n4765 11.6369
R9175 AVSS.n4765 AVSS.n4730 11.6369
R9176 AVSS.n4730 AVSS.n4728 11.6369
R9177 AVSS.n4776 AVSS.n4728 11.6369
R9178 AVSS.n4777 AVSS.n4776 11.6369
R9179 AVSS.n4779 AVSS.n4777 11.6369
R9180 AVSS.n4779 AVSS.n4778 11.6369
R9181 AVSS.n4778 AVSS.n4724 11.6369
R9182 AVSS.n4787 AVSS.n4786 11.6369
R9183 AVSS.n4790 AVSS.n4787 11.6369
R9184 AVSS.n4791 AVSS.n4790 11.6369
R9185 AVSS.n4794 AVSS.n4791 11.6369
R9186 AVSS.n4795 AVSS.n4794 11.6369
R9187 AVSS.n4798 AVSS.n4795 11.6369
R9188 AVSS.n4799 AVSS.n4798 11.6369
R9189 AVSS.n4802 AVSS.n4799 11.6369
R9190 AVSS.n4803 AVSS.n4802 11.6369
R9191 AVSS.n4806 AVSS.n4803 11.6369
R9192 AVSS.n4931 AVSS.n1371 11.6369
R9193 AVSS.n4910 AVSS.n4909 11.6369
R9194 AVSS.n4913 AVSS.n4910 11.6369
R9195 AVSS.n4914 AVSS.n4913 11.6369
R9196 AVSS.n4917 AVSS.n4914 11.6369
R9197 AVSS.n4918 AVSS.n4917 11.6369
R9198 AVSS.n4921 AVSS.n4918 11.6369
R9199 AVSS.n4923 AVSS.n4922 11.6369
R9200 AVSS.n4923 AVSS.n1372 11.6369
R9201 AVSS.n4929 AVSS.n1372 11.6369
R9202 AVSS.n4930 AVSS.n4929 11.6369
R9203 AVSS.n1885 AVSS.n1854 11.6369
R9204 AVSS.n1879 AVSS.n1854 11.6369
R9205 AVSS.n1879 AVSS.n1878 11.6369
R9206 AVSS.n1878 AVSS.n1877 11.6369
R9207 AVSS.n1877 AVSS.n1856 11.6369
R9208 AVSS.n1871 AVSS.n1856 11.6369
R9209 AVSS.n1871 AVSS.n1870 11.6369
R9210 AVSS.n1870 AVSS.n1869 11.6369
R9211 AVSS.n1869 AVSS.n1858 11.6369
R9212 AVSS.n1863 AVSS.n1862 11.6369
R9213 AVSS.n2566 AVSS.n2563 11.6369
R9214 AVSS.n2567 AVSS.n2566 11.6369
R9215 AVSS.n2570 AVSS.n2567 11.6369
R9216 AVSS.n2571 AVSS.n2570 11.6369
R9217 AVSS.n2574 AVSS.n2571 11.6369
R9218 AVSS.n2577 AVSS.n2576 11.6369
R9219 AVSS.n2579 AVSS.n2577 11.6369
R9220 AVSS.n2579 AVSS.n2578 11.6369
R9221 AVSS.n1843 AVSS.n1840 11.6369
R9222 AVSS.n1840 AVSS.n1839 11.6369
R9223 AVSS.n1839 AVSS.n1836 11.6369
R9224 AVSS.n1836 AVSS.n1835 11.6369
R9225 AVSS.n1835 AVSS.n1832 11.6369
R9226 AVSS.n1832 AVSS.n1831 11.6369
R9227 AVSS.n1831 AVSS.n1828 11.6369
R9228 AVSS.n1828 AVSS.n1827 11.6369
R9229 AVSS.n1827 AVSS.n1739 11.6369
R9230 AVSS.n2588 AVSS.n2586 11.6369
R9231 AVSS.n2520 AVSS.n1852 11.6369
R9232 AVSS.n2521 AVSS.n2520 11.6369
R9233 AVSS.n2522 AVSS.n2521 11.6369
R9234 AVSS.n2522 AVSS.n1850 11.6369
R9235 AVSS.n2528 AVSS.n1850 11.6369
R9236 AVSS.n2529 AVSS.n2528 11.6369
R9237 AVSS.n2530 AVSS.n2529 11.6369
R9238 AVSS.n2530 AVSS.n1848 11.6369
R9239 AVSS.n1848 AVSS.n1824 11.6369
R9240 AVSS.n6188 AVSS.n159 11.6369
R9241 AVSS.n6182 AVSS.n159 11.6369
R9242 AVSS.n6182 AVSS.n6181 11.6369
R9243 AVSS.n6181 AVSS.n6180 11.6369
R9244 AVSS.n6180 AVSS.n164 11.6369
R9245 AVSS.n6174 AVSS.n164 11.6369
R9246 AVSS.n6173 AVSS.n6172 11.6369
R9247 AVSS.n6172 AVSS.n171 11.6369
R9248 AVSS.n6166 AVSS.n171 11.6369
R9249 AVSS.n6166 AVSS.n6165 11.6369
R9250 AVSS.n6141 AVSS.n6140 11.6369
R9251 AVSS.n6142 AVSS.n6141 11.6369
R9252 AVSS.n6142 AVSS.n181 11.6369
R9253 AVSS.n6148 AVSS.n181 11.6369
R9254 AVSS.n6149 AVSS.n6148 11.6369
R9255 AVSS.n6150 AVSS.n6149 11.6369
R9256 AVSS.n6150 AVSS.n179 11.6369
R9257 AVSS.n6156 AVSS.n179 11.6369
R9258 AVSS.n6157 AVSS.n6156 11.6369
R9259 AVSS.n6158 AVSS.n6157 11.6369
R9260 AVSS.n6158 AVSS.n175 11.6369
R9261 AVSS.n6164 AVSS.n175 11.6369
R9262 AVSS.n260 AVSS.n233 11.6369
R9263 AVSS.n252 AVSS.n233 11.6369
R9264 AVSS.n252 AVSS.n251 11.6369
R9265 AVSS.n251 AVSS.n250 11.6369
R9266 AVSS.n250 AVSS.n235 11.6369
R9267 AVSS.n244 AVSS.n235 11.6369
R9268 AVSS.n244 AVSS.n243 11.6369
R9269 AVSS.n243 AVSS.n242 11.6369
R9270 AVSS.n242 AVSS.n237 11.6369
R9271 AVSS.n237 AVSS.n185 11.6369
R9272 AVSS.n6209 AVSS.n149 11.6369
R9273 AVSS.n6204 AVSS.n149 11.6369
R9274 AVSS.n6204 AVSS.n6203 11.6369
R9275 AVSS.n6203 AVSS.n6202 11.6369
R9276 AVSS.n6202 AVSS.n153 11.6369
R9277 AVSS.n6197 AVSS.n153 11.6369
R9278 AVSS.n6197 AVSS.n6196 11.6369
R9279 AVSS.n6196 AVSS.n6195 11.6369
R9280 AVSS.n6195 AVSS.n156 11.6369
R9281 AVSS.n6190 AVSS.n156 11.6369
R9282 AVSS.n6190 AVSS.n6189 11.6369
R9283 AVSS.n4291 AVSS.n4290 11.6369
R9284 AVSS.n4290 AVSS.n4289 11.6369
R9285 AVSS.n4289 AVSS.n3893 11.6369
R9286 AVSS.n4284 AVSS.n3893 11.6369
R9287 AVSS.n4284 AVSS.n4283 11.6369
R9288 AVSS.n4283 AVSS.n4282 11.6369
R9289 AVSS.n4282 AVSS.n3896 11.6369
R9290 AVSS.n4277 AVSS.n3896 11.6369
R9291 AVSS.n4277 AVSS.n4276 11.6369
R9292 AVSS.n4276 AVSS.n4275 11.6369
R9293 AVSS.n4275 AVSS.n3899 11.6369
R9294 AVSS.n4270 AVSS.n3899 11.6369
R9295 AVSS.n3989 AVSS.n3902 11.6369
R9296 AVSS.n3983 AVSS.n3902 11.6369
R9297 AVSS.n3983 AVSS.n3982 11.6369
R9298 AVSS.n3982 AVSS.n3981 11.6369
R9299 AVSS.n3981 AVSS.n3904 11.6369
R9300 AVSS.n3975 AVSS.n3974 11.6369
R9301 AVSS.n3974 AVSS.n3973 11.6369
R9302 AVSS.n3973 AVSS.n3906 11.6369
R9303 AVSS.n3967 AVSS.n3906 11.6369
R9304 AVSS.n3943 AVSS.n3942 11.6369
R9305 AVSS.n3943 AVSS.n3916 11.6369
R9306 AVSS.n3949 AVSS.n3916 11.6369
R9307 AVSS.n3950 AVSS.n3949 11.6369
R9308 AVSS.n3951 AVSS.n3950 11.6369
R9309 AVSS.n3951 AVSS.n3912 11.6369
R9310 AVSS.n3957 AVSS.n3912 11.6369
R9311 AVSS.n3958 AVSS.n3957 11.6369
R9312 AVSS.n3959 AVSS.n3958 11.6369
R9313 AVSS.n3959 AVSS.n3908 11.6369
R9314 AVSS.n3965 AVSS.n3908 11.6369
R9315 AVSS.n3966 AVSS.n3965 11.6369
R9316 AVSS.n4296 AVSS.n3890 11.6369
R9317 AVSS.n3925 AVSS.n3890 11.6369
R9318 AVSS.n3926 AVSS.n3925 11.6369
R9319 AVSS.n3926 AVSS.n3922 11.6369
R9320 AVSS.n3932 AVSS.n3922 11.6369
R9321 AVSS.n3933 AVSS.n3932 11.6369
R9322 AVSS.n3934 AVSS.n3933 11.6369
R9323 AVSS.n3934 AVSS.n3920 11.6369
R9324 AVSS.n3920 AVSS.n3919 11.6369
R9325 AVSS.n3941 AVSS.n3919 11.6369
R9326 AVSS.n4324 AVSS.n4323 11.6369
R9327 AVSS.n4323 AVSS.n4322 11.6369
R9328 AVSS.n4322 AVSS.n3682 11.6369
R9329 AVSS.n4317 AVSS.n3682 11.6369
R9330 AVSS.n4317 AVSS.n4316 11.6369
R9331 AVSS.n4316 AVSS.n4315 11.6369
R9332 AVSS.n4315 AVSS.n3685 11.6369
R9333 AVSS.n4310 AVSS.n3685 11.6369
R9334 AVSS.n4310 AVSS.n4309 11.6369
R9335 AVSS.n4309 AVSS.n4308 11.6369
R9336 AVSS.n4308 AVSS.n3688 11.6369
R9337 AVSS.n4303 AVSS.n3688 11.6369
R9338 AVSS.n3778 AVSS.n3691 11.6369
R9339 AVSS.n3772 AVSS.n3691 11.6369
R9340 AVSS.n3772 AVSS.n3771 11.6369
R9341 AVSS.n3771 AVSS.n3770 11.6369
R9342 AVSS.n3770 AVSS.n3693 11.6369
R9343 AVSS.n3764 AVSS.n3763 11.6369
R9344 AVSS.n3763 AVSS.n3762 11.6369
R9345 AVSS.n3762 AVSS.n3695 11.6369
R9346 AVSS.n3756 AVSS.n3695 11.6369
R9347 AVSS.n3732 AVSS.n3731 11.6369
R9348 AVSS.n3732 AVSS.n3705 11.6369
R9349 AVSS.n3738 AVSS.n3705 11.6369
R9350 AVSS.n3739 AVSS.n3738 11.6369
R9351 AVSS.n3740 AVSS.n3739 11.6369
R9352 AVSS.n3740 AVSS.n3701 11.6369
R9353 AVSS.n3746 AVSS.n3701 11.6369
R9354 AVSS.n3747 AVSS.n3746 11.6369
R9355 AVSS.n3748 AVSS.n3747 11.6369
R9356 AVSS.n3748 AVSS.n3697 11.6369
R9357 AVSS.n3754 AVSS.n3697 11.6369
R9358 AVSS.n3755 AVSS.n3754 11.6369
R9359 AVSS.n4329 AVSS.n3679 11.6369
R9360 AVSS.n3714 AVSS.n3679 11.6369
R9361 AVSS.n3715 AVSS.n3714 11.6369
R9362 AVSS.n3715 AVSS.n3711 11.6369
R9363 AVSS.n3721 AVSS.n3711 11.6369
R9364 AVSS.n3722 AVSS.n3721 11.6369
R9365 AVSS.n3723 AVSS.n3722 11.6369
R9366 AVSS.n3723 AVSS.n3709 11.6369
R9367 AVSS.n3709 AVSS.n3708 11.6369
R9368 AVSS.n3730 AVSS.n3708 11.6369
R9369 AVSS.n3640 AVSS.n3515 11.6369
R9370 AVSS.n3635 AVSS.n3515 11.6369
R9371 AVSS.n3635 AVSS.n3634 11.6369
R9372 AVSS.n3634 AVSS.n3633 11.6369
R9373 AVSS.n3633 AVSS.n3517 11.6369
R9374 AVSS.n3627 AVSS.n3626 11.6369
R9375 AVSS.n3626 AVSS.n3625 11.6369
R9376 AVSS.n3625 AVSS.n3519 11.6369
R9377 AVSS.n3619 AVSS.n3519 11.6369
R9378 AVSS.n3593 AVSS.n3577 11.6369
R9379 AVSS.n3587 AVSS.n3577 11.6369
R9380 AVSS.n3587 AVSS.n3586 11.6369
R9381 AVSS.n3586 AVSS.n3585 11.6369
R9382 AVSS.n3585 AVSS.n3581 11.6369
R9383 AVSS.n3581 AVSS.n3525 11.6369
R9384 AVSS.n3609 AVSS.n3525 11.6369
R9385 AVSS.n3610 AVSS.n3609 11.6369
R9386 AVSS.n3611 AVSS.n3610 11.6369
R9387 AVSS.n3611 AVSS.n3521 11.6369
R9388 AVSS.n3617 AVSS.n3521 11.6369
R9389 AVSS.n3618 AVSS.n3617 11.6369
R9390 AVSS.n3564 AVSS.n3563 11.6369
R9391 AVSS.n3565 AVSS.n3564 11.6369
R9392 AVSS.n3565 AVSS.n3532 11.6369
R9393 AVSS.n3571 AVSS.n3532 11.6369
R9394 AVSS.n3572 AVSS.n3571 11.6369
R9395 AVSS.n3603 AVSS.n3572 11.6369
R9396 AVSS.n3603 AVSS.n3602 11.6369
R9397 AVSS.n3602 AVSS.n3601 11.6369
R9398 AVSS.n3601 AVSS.n3573 11.6369
R9399 AVSS.n3595 AVSS.n3573 11.6369
R9400 AVSS.n3595 AVSS.n3594 11.6369
R9401 AVSS.n3537 AVSS.n3536 11.6369
R9402 AVSS.n3556 AVSS.n3537 11.6369
R9403 AVSS.n3556 AVSS.n3555 11.6369
R9404 AVSS.n3555 AVSS.n3554 11.6369
R9405 AVSS.n3554 AVSS.n3539 11.6369
R9406 AVSS.n3549 AVSS.n3539 11.6369
R9407 AVSS.n3549 AVSS.n3548 11.6369
R9408 AVSS.n3548 AVSS.n3547 11.6369
R9409 AVSS.n3547 AVSS.n3542 11.6369
R9410 AVSS.n3542 AVSS.n3511 11.6369
R9411 AVSS.n4340 AVSS.n3512 11.6369
R9412 AVSS.n4258 AVSS.n4257 11.6369
R9413 AVSS.n4257 AVSS.n4231 11.6369
R9414 AVSS.n4252 AVSS.n4231 11.6369
R9415 AVSS.n4252 AVSS.n4251 11.6369
R9416 AVSS.n4251 AVSS.n4250 11.6369
R9417 AVSS.n4250 AVSS.n4233 11.6369
R9418 AVSS.n4244 AVSS.n4233 11.6369
R9419 AVSS.n4244 AVSS.n4243 11.6369
R9420 AVSS.n4243 AVSS.n4242 11.6369
R9421 AVSS.n4242 AVSS.n4235 11.6369
R9422 AVSS.n4236 AVSS.n4235 11.6369
R9423 AVSS.n4236 AVSS.n230 11.6369
R9424 AVSS.n4263 AVSS.n4207 11.6369
R9425 AVSS.n4226 AVSS.n4207 11.6369
R9426 AVSS.n4226 AVSS.n4225 11.6369
R9427 AVSS.n4225 AVSS.n4224 11.6369
R9428 AVSS.n4224 AVSS.n4209 11.6369
R9429 AVSS.n4218 AVSS.n4209 11.6369
R9430 AVSS.n4218 AVSS.n4217 11.6369
R9431 AVSS.n4217 AVSS.n4216 11.6369
R9432 AVSS.n4216 AVSS.n4211 11.6369
R9433 AVSS.n4211 AVSS.n213 11.6369
R9434 AVSS.n6135 AVSS.n6134 11.6369
R9435 AVSS.n6134 AVSS.n6133 11.6369
R9436 AVSS.n6133 AVSS.n214 11.6369
R9437 AVSS.n6127 AVSS.n214 11.6369
R9438 AVSS.n6127 AVSS.n6126 11.6369
R9439 AVSS.n6126 AVSS.n6125 11.6369
R9440 AVSS.n6125 AVSS.n218 11.6369
R9441 AVSS.n6119 AVSS.n218 11.6369
R9442 AVSS.n6119 AVSS.n6118 11.6369
R9443 AVSS.n6118 AVSS.n6117 11.6369
R9444 AVSS.n6117 AVSS.n222 11.6369
R9445 AVSS.n6111 AVSS.n222 11.6369
R9446 AVSS.n6093 AVSS.n228 11.6369
R9447 AVSS.n6094 AVSS.n6093 11.6369
R9448 AVSS.n6095 AVSS.n6094 11.6369
R9449 AVSS.n6095 AVSS.n226 11.6369
R9450 AVSS.n6101 AVSS.n226 11.6369
R9451 AVSS.n6103 AVSS.n6102 11.6369
R9452 AVSS.n6103 AVSS.n224 11.6369
R9453 AVSS.n6109 AVSS.n224 11.6369
R9454 AVSS.n6110 AVSS.n6109 11.6369
R9455 AVSS.n4363 AVSS.n4360 11.6369
R9456 AVSS.n4387 AVSS.n4363 11.6369
R9457 AVSS.n4387 AVSS.n4386 11.6369
R9458 AVSS.n4386 AVSS.n4385 11.6369
R9459 AVSS.n4385 AVSS.n4364 11.6369
R9460 AVSS.n4366 AVSS.n4364 11.6369
R9461 AVSS.n4369 AVSS.n4366 11.6369
R9462 AVSS.n4375 AVSS.n4369 11.6369
R9463 AVSS.n4375 AVSS.n4374 11.6369
R9464 AVSS.n4374 AVSS.n4373 11.6369
R9465 AVSS.n4373 AVSS.n3302 11.6369
R9466 AVSS.n4396 AVSS.n4358 11.6369
R9467 AVSS.n4397 AVSS.n4396 11.6369
R9468 AVSS.n4398 AVSS.n4397 11.6369
R9469 AVSS.n4398 AVSS.n4356 11.6369
R9470 AVSS.n4404 AVSS.n4356 11.6369
R9471 AVSS.n4405 AVSS.n4404 11.6369
R9472 AVSS.n4406 AVSS.n4405 11.6369
R9473 AVSS.n4406 AVSS.n4354 11.6369
R9474 AVSS.n4412 AVSS.n4354 11.6369
R9475 AVSS.n4413 AVSS.n4412 11.6369
R9476 AVSS.n4415 AVSS.n4352 11.6369
R9477 AVSS.n4422 AVSS.n4421 11.6369
R9478 AVSS.n4423 AVSS.n4422 11.6369
R9479 AVSS.n4423 AVSS.n4350 11.6369
R9480 AVSS.n4429 AVSS.n4350 11.6369
R9481 AVSS.n4430 AVSS.n4429 11.6369
R9482 AVSS.n4431 AVSS.n4430 11.6369
R9483 AVSS.n4437 AVSS.n4348 11.6369
R9484 AVSS.n4438 AVSS.n4437 11.6369
R9485 AVSS.n4439 AVSS.n4438 11.6369
R9486 AVSS.n4439 AVSS.n4346 11.6369
R9487 AVSS.n4466 AVSS.n4465 11.6369
R9488 AVSS.n4465 AVSS.n4464 11.6369
R9489 AVSS.n4464 AVSS.n4461 11.6369
R9490 AVSS.n4461 AVSS.n4460 11.6369
R9491 AVSS.n4460 AVSS.n4457 11.6369
R9492 AVSS.n4457 AVSS.n4456 11.6369
R9493 AVSS.n4456 AVSS.n4453 11.6369
R9494 AVSS.n4453 AVSS.n4452 11.6369
R9495 AVSS.n4452 AVSS.n4449 11.6369
R9496 AVSS.n4449 AVSS.n4448 11.6369
R9497 AVSS.n4445 AVSS.n4444 11.6369
R9498 AVSS.n6051 AVSS.n5930 10.6369
R9499 AVSS.n6020 AVSS.n5930 10.6369
R9500 AVSS.n5931 AVSS.n5929 10.6369
R9501 AVSS.n6014 AVSS.n5929 10.6369
R9502 AVSS.n6029 AVSS.n6028 10.4516
R9503 AVSS AVSS.n1152 10.3439
R9504 AVSS.n4945 AVSS 10.3439
R9505 AVSS AVSS.n2172 10.3439
R9506 AVSS AVSS.n5600 10.3439
R9507 AVSS.n5427 AVSS 10.3439
R9508 AVSS AVSS.n5203 10.3439
R9509 AVSS.n5885 AVSS 10.3439
R9510 AVSS AVSS.n5634 10.3439
R9511 AVSS.n874 AVSS 10.3439
R9512 AVSS AVSS.n2240 10.3439
R9513 AVSS AVSS.n2306 10.3439
R9514 AVSS AVSS.n1386 10.3439
R9515 AVSS.n5000 AVSS 10.3439
R9516 AVSS AVSS.n3077 10.3439
R9517 AVSS.n2890 AVSS 10.3439
R9518 AVSS AVSS.n3015 10.3439
R9519 AVSS.n2820 AVSS 10.3439
R9520 AVSS.n4922 AVSS 10.3439
R9521 AVSS.n2576 AVSS 10.3439
R9522 AVSS AVSS.n6173 10.3439
R9523 AVSS.n3975 AVSS 10.3439
R9524 AVSS.n3764 AVSS 10.3439
R9525 AVSS.n3627 AVSS 10.3439
R9526 AVSS.n6102 AVSS 10.3439
R9527 AVSS AVSS.n4348 10.3439
R9528 AVSS.n5392 AVSS.n5391 10.1338
R9529 AVSS.n5193 AVSS.n5192 10.1338
R9530 AVSS.n551 AVSS.n550 10.1338
R9531 AVSS.n1460 AVSS.n1459 10.1338
R9532 AVSS.n4880 AVSS.n4879 10.1338
R9533 AVSS.n2047 AVSS.n2046 10.1338
R9534 AVSS.n2453 AVSS.n2452 10.1338
R9535 AVSS.n1975 AVSS.n1974 10.1338
R9536 AVSS.n1806 AVSS.n1788 10.1338
R9537 AVSS.n3394 AVSS.n3393 10.1338
R9538 AVSS.n6063 AVSS.n6062 10.1119
R9539 AVSS.n1322 AVSS.n1158 10.0853
R9540 AVSS.n4959 AVSS.n4958 10.0853
R9541 AVSS.n2072 AVSS.n2070 10.0853
R9542 AVSS.n5614 AVSS.n5613 10.0853
R9543 AVSS.n5443 AVSS.n5442 10.0853
R9544 AVSS.n5217 AVSS.n5216 10.0853
R9545 AVSS.n5899 AVSS.n5898 10.0853
R9546 AVSS.n5677 AVSS.n5641 10.0853
R9547 AVSS.n856 AVSS.n680 10.0853
R9548 AVSS.n2254 AVSS.n2201 10.0853
R9549 AVSS.n2391 AVSS.n2387 10.0853
R9550 AVSS.n1566 AVSS.n1562 10.0853
R9551 AVSS.n5014 AVSS.n5013 10.0853
R9552 AVSS.n3246 AVSS.n3084 10.0853
R9553 AVSS.n4503 AVSS.n4502 10.0853
R9554 AVSS.n4683 AVSS.n4682 10.0853
R9555 AVSS.n4714 AVSS.n1717 10.0853
R9556 AVSS.n4909 AVSS.n1379 10.0853
R9557 AVSS.n1862 AVSS.n1747 10.0853
R9558 AVSS.n6189 AVSS.n6188 10.0853
R9559 AVSS.n4270 AVSS.n4269 10.0853
R9560 AVSS.n4303 AVSS.n4302 10.0853
R9561 AVSS.n4335 AVSS.n3512 10.0853
R9562 AVSS.n6087 AVSS.n230 10.0853
R9563 AVSS.n4421 AVSS.n4352 10.0853
R9564 AVSS.n146 AVSS.n56 9.95606
R9565 AVSS.n4204 AVSS.n4114 9.95606
R9566 AVSS.n4062 AVSS.n4061 9.95606
R9567 AVSS.n3851 AVSS.n3850 9.95606
R9568 AVSS.n3214 AVSS.n3123 9.95606
R9569 AVSS.n1290 AVSS.n1199 9.95606
R9570 AVSS.n4595 AVSS.n4594 9.95606
R9571 AVSS.n2774 AVSS.n2684 9.95606
R9572 AVSS.n2664 AVSS.n2663 9.95606
R9573 AVSS.n831 AVSS.n740 9.95606
R9574 AVSS.n1787 AVSS.n1786 9.95606
R9575 AVSS.n1340 AVSS.n1148 9.56818
R9576 AVSS.n4938 AVSS.n4937 9.56818
R9577 AVSS.n2165 AVSS.n2161 9.56818
R9578 AVSS.n5849 AVSS.n5258 9.56818
R9579 AVSS.n5419 AVSS.n5418 9.56818
R9580 AVSS.n5225 AVSS.n409 9.56818
R9581 AVSS.n5878 AVSS.n5877 9.56818
R9582 AVSS.n5696 AVSS.n5630 9.56818
R9583 AVSS.n883 AVSS.n882 9.56818
R9584 AVSS.n2233 AVSS.n2229 9.56818
R9585 AVSS.n2413 AVSS.n2304 9.56818
R9586 AVSS.n1589 AVSS.n1384 9.56818
R9587 AVSS.n4993 AVSS.n4992 9.56818
R9588 AVSS.n3265 AVSS.n3073 9.56818
R9589 AVSS.n2899 AVSS.n2898 9.56818
R9590 AVSS.n3041 AVSS.n3013 9.56818
R9591 AVSS.n4473 AVSS.n4472 9.56818
R9592 AVSS.n4931 AVSS.n4930 9.56818
R9593 AVSS.n2586 AVSS.n2585 9.56818
R9594 AVSS.n6165 AVSS.n6164 9.56818
R9595 AVSS.n3967 AVSS.n3966 9.56818
R9596 AVSS.n3756 AVSS.n3755 9.56818
R9597 AVSS.n3619 AVSS.n3618 9.56818
R9598 AVSS.n6111 AVSS.n6110 9.56818
R9599 AVSS.n4444 AVSS.n4346 9.56818
R9600 AVSS.n2562 AVSS.n2561 9.52371
R9601 AVSS.n1740 AVSS.n1738 9.52371
R9602 AVSS.n2513 AVSS.n1749 9.52223
R9603 AVSS.n2539 AVSS.n2538 9.52223
R9604 AVSS.n3510 AVSS.n3509 9.47828
R9605 AVSS.n3666 AVSS.n3663 9.33749
R9606 AVSS.n553 AVSS.n551 9.30178
R9607 AVSS.n589 AVSS.n575 9.3005
R9608 AVSS.n575 AVSS.n573 9.3005
R9609 AVSS.n587 AVSS.n575 9.3005
R9610 AVSS.n584 AVSS.n44 9.3005
R9611 AVSS.n589 AVSS.n44 9.3005
R9612 AVSS.n573 AVSS.n44 9.3005
R9613 AVSS.n587 AVSS.n44 9.3005
R9614 AVSS.n584 AVSS.n45 9.3005
R9615 AVSS.n589 AVSS.n45 9.3005
R9616 AVSS.n573 AVSS.n45 9.3005
R9617 AVSS.n587 AVSS.n45 9.3005
R9618 AVSS.n589 AVSS.n576 9.3005
R9619 AVSS.n576 AVSS.n573 9.3005
R9620 AVSS.n587 AVSS.n576 9.3005
R9621 AVSS.n589 AVSS.n574 9.3005
R9622 AVSS.n574 AVSS.n573 9.3005
R9623 AVSS.n580 AVSS.n574 9.3005
R9624 AVSS.n587 AVSS.n574 9.3005
R9625 AVSS.n589 AVSS.n588 9.3005
R9626 AVSS.n588 AVSS.n573 9.3005
R9627 AVSS.n588 AVSS.n580 9.3005
R9628 AVSS.n588 AVSS.n587 9.3005
R9629 AVSS.n1110 AVSS.n1096 9.3005
R9630 AVSS.n1096 AVSS.n1094 9.3005
R9631 AVSS.n1108 AVSS.n1096 9.3005
R9632 AVSS.n1105 AVSS.n48 9.3005
R9633 AVSS.n1110 AVSS.n48 9.3005
R9634 AVSS.n1094 AVSS.n48 9.3005
R9635 AVSS.n1108 AVSS.n48 9.3005
R9636 AVSS.n1105 AVSS.n49 9.3005
R9637 AVSS.n1110 AVSS.n49 9.3005
R9638 AVSS.n1094 AVSS.n49 9.3005
R9639 AVSS.n1108 AVSS.n49 9.3005
R9640 AVSS.n1110 AVSS.n1097 9.3005
R9641 AVSS.n1097 AVSS.n1094 9.3005
R9642 AVSS.n1108 AVSS.n1097 9.3005
R9643 AVSS.n1110 AVSS.n1095 9.3005
R9644 AVSS.n1095 AVSS.n1094 9.3005
R9645 AVSS.n1101 AVSS.n1095 9.3005
R9646 AVSS.n1108 AVSS.n1095 9.3005
R9647 AVSS.n1110 AVSS.n1109 9.3005
R9648 AVSS.n1109 AVSS.n1094 9.3005
R9649 AVSS.n1109 AVSS.n1101 9.3005
R9650 AVSS.n1109 AVSS.n1108 9.3005
R9651 AVSS.n777 AVSS.n739 9.3005
R9652 AVSS.n832 AVSS.n831 9.3005
R9653 AVSS.n5726 AVSS.n5725 9.3005
R9654 AVSS.n834 AVSS.n833 9.3005
R9655 AVSS.n738 AVSS.n737 9.3005
R9656 AVSS.n2193 AVSS.n1975 9.3005
R9657 AVSS.n2453 AVSS.n2416 9.3005
R9658 AVSS.n2509 AVSS.n2508 9.3005
R9659 AVSS.n1066 AVSS.n1065 9.3005
R9660 AVSS.n2194 AVSS.n645 9.3005
R9661 AVSS.n2342 AVSS.n2195 9.3005
R9662 AVSS.n2415 AVSS.n2414 9.3005
R9663 AVSS.n2302 AVSS.n2301 9.3005
R9664 AVSS.n2046 AVSS.n1976 9.3005
R9665 AVSS.n2068 AVSS.n2067 9.3005
R9666 AVSS.n2081 AVSS.n1624 9.3005
R9667 AVSS.n2190 AVSS.n2189 9.3005
R9668 AVSS.n2192 AVSS.n646 9.3005
R9669 AVSS.n4721 AVSS.n4720 9.3005
R9670 AVSS.n1861 AVSS.n1748 9.3005
R9671 AVSS.n2511 AVSS.n2510 9.3005
R9672 AVSS.n1844 AVSS.n1823 9.3005
R9673 AVSS.n1786 AVSS.n1749 9.3005
R9674 AVSS.n2561 AVSS.n2560 9.3005
R9675 AVSS.n1788 AVSS.n1738 9.3005
R9676 AVSS.n2540 AVSS.n2539 9.3005
R9677 AVSS.n2590 AVSS.n2589 9.3005
R9678 AVSS.n1715 AVSS.n1714 9.3005
R9679 AVSS.n2664 AVSS.n1722 9.3005
R9680 AVSS.n2683 AVSS.n2682 9.3005
R9681 AVSS.n2775 AVSS.n2774 9.3005
R9682 AVSS.n4713 AVSS.n4712 9.3005
R9683 AVSS.n4711 AVSS.n4710 9.3005
R9684 AVSS.n4681 AVSS.n4680 9.3005
R9685 AVSS.n4679 AVSS.n4678 9.3005
R9686 AVSS.n4616 AVSS.n4615 9.3005
R9687 AVSS.n4594 AVSS.n1067 9.3005
R9688 AVSS.n4668 AVSS.n4667 9.3005
R9689 AVSS.n4982 AVSS.n4981 9.3005
R9690 AVSS.n4671 AVSS.n4670 9.3005
R9691 AVSS.n4985 AVSS.n4984 9.3005
R9692 AVSS.n1236 AVSS.n1198 9.3005
R9693 AVSS.n1291 AVSS.n1290 9.3005
R9694 AVSS.n1197 AVSS.n1147 9.3005
R9695 AVSS.n1293 AVSS.n1292 9.3005
R9696 AVSS.n3160 AVSS.n3122 9.3005
R9697 AVSS.n3215 AVSS.n3214 9.3005
R9698 AVSS.n3072 AVSS.n55 9.3005
R9699 AVSS.n3217 AVSS.n3216 9.3005
R9700 AVSS.n4495 AVSS.n4481 9.3005
R9701 AVSS.n4481 AVSS.n4479 9.3005
R9702 AVSS.n4493 AVSS.n4481 9.3005
R9703 AVSS.n4490 AVSS.n52 9.3005
R9704 AVSS.n4495 AVSS.n52 9.3005
R9705 AVSS.n4479 AVSS.n52 9.3005
R9706 AVSS.n4493 AVSS.n52 9.3005
R9707 AVSS.n4490 AVSS.n53 9.3005
R9708 AVSS.n4495 AVSS.n53 9.3005
R9709 AVSS.n4479 AVSS.n53 9.3005
R9710 AVSS.n4493 AVSS.n53 9.3005
R9711 AVSS.n4495 AVSS.n4482 9.3005
R9712 AVSS.n4482 AVSS.n4479 9.3005
R9713 AVSS.n4493 AVSS.n4482 9.3005
R9714 AVSS.n4495 AVSS.n4480 9.3005
R9715 AVSS.n4480 AVSS.n4479 9.3005
R9716 AVSS.n4486 AVSS.n4480 9.3005
R9717 AVSS.n4493 AVSS.n4480 9.3005
R9718 AVSS.n4495 AVSS.n4494 9.3005
R9719 AVSS.n4494 AVSS.n4479 9.3005
R9720 AVSS.n4494 AVSS.n4486 9.3005
R9721 AVSS.n4494 AVSS.n4493 9.3005
R9722 AVSS.n6211 AVSS.n6210 9.3005
R9723 AVSS.n3395 AVSS.n3394 9.3005
R9724 AVSS.n3343 AVSS.n3303 9.3005
R9725 AVSS.n4345 AVSS.n4344 9.3005
R9726 AVSS.n4414 AVSS.n1623 9.3005
R9727 AVSS.n4879 AVSS.n4809 9.3005
R9728 AVSS.n4901 AVSS.n4900 9.3005
R9729 AVSS.n4808 AVSS.n4807 9.3005
R9730 AVSS.n4903 AVSS.n4902 9.3005
R9731 AVSS.n1459 AVSS.n1382 9.3005
R9732 AVSS.n1481 AVSS.n1480 9.3005
R9733 AVSS.n1594 AVSS.n1593 9.3005
R9734 AVSS.n1483 AVSS.n1482 9.3005
R9735 AVSS.n4342 AVSS.n4341 9.3005
R9736 AVSS.n554 AVSS.n326 9.3005
R9737 AVSS.n5194 AVSS.n5193 9.3005
R9738 AVSS.n5175 AVSS.n5101 9.3005
R9739 AVSS.n5393 AVSS.n5392 9.3005
R9740 AVSS.n5374 AVSS.n1 9.3005
R9741 AVSS.n5546 AVSS.n5545 9.3005
R9742 AVSS.n5818 AVSS.n5817 9.3005
R9743 AVSS.n552 AVSS.n325 9.3005
R9744 AVSS.n5100 AVSS.n5099 9.3005
R9745 AVSS.n5196 AVSS.n5195 9.3005
R9746 AVSS.n6303 AVSS.n6302 9.3005
R9747 AVSS.n5395 AVSS.n5394 9.3005
R9748 AVSS.n5548 AVSS.n5547 9.3005
R9749 AVSS.n5820 AVSS.n5819 9.3005
R9750 AVSS.n564 AVSS.n559 9.3005
R9751 AVSS.n564 AVSS.n557 9.3005
R9752 AVSS.n564 AVSS.n560 9.3005
R9753 AVSS.n5025 AVSS.n564 9.3005
R9754 AVSS.n566 AVSS.n559 9.3005
R9755 AVSS.n566 AVSS.n557 9.3005
R9756 AVSS.n566 AVSS.n560 9.3005
R9757 AVSS.n5025 AVSS.n566 9.3005
R9758 AVSS.n563 AVSS.n559 9.3005
R9759 AVSS.n563 AVSS.n557 9.3005
R9760 AVSS.n563 AVSS.n560 9.3005
R9761 AVSS.n5025 AVSS.n563 9.3005
R9762 AVSS.n5024 AVSS.n559 9.3005
R9763 AVSS.n5024 AVSS.n557 9.3005
R9764 AVSS.n5024 AVSS.n560 9.3005
R9765 AVSS.n5025 AVSS.n5024 9.3005
R9766 AVSS.n562 AVSS.n559 9.3005
R9767 AVSS.n562 AVSS.n557 9.3005
R9768 AVSS.n562 AVSS.n560 9.3005
R9769 AVSS.n562 AVSS.n556 9.3005
R9770 AVSS.n5025 AVSS.n562 9.3005
R9771 AVSS.n5026 AVSS.n559 9.3005
R9772 AVSS.n5026 AVSS.n557 9.3005
R9773 AVSS.n5026 AVSS.n560 9.3005
R9774 AVSS.n5026 AVSS.n556 9.3005
R9775 AVSS.n5026 AVSS.n5025 9.3005
R9776 AVSS.n1605 AVSS.n1599 9.3005
R9777 AVSS.n1605 AVSS.n1598 9.3005
R9778 AVSS.n1605 AVSS.n1600 9.3005
R9779 AVSS.n1620 AVSS.n1605 9.3005
R9780 AVSS.n1607 AVSS.n1599 9.3005
R9781 AVSS.n1607 AVSS.n1598 9.3005
R9782 AVSS.n1607 AVSS.n1600 9.3005
R9783 AVSS.n1620 AVSS.n1607 9.3005
R9784 AVSS.n1604 AVSS.n1599 9.3005
R9785 AVSS.n1604 AVSS.n1598 9.3005
R9786 AVSS.n1604 AVSS.n1600 9.3005
R9787 AVSS.n1620 AVSS.n1604 9.3005
R9788 AVSS.n1609 AVSS.n1599 9.3005
R9789 AVSS.n1609 AVSS.n1598 9.3005
R9790 AVSS.n1609 AVSS.n1600 9.3005
R9791 AVSS.n1620 AVSS.n1609 9.3005
R9792 AVSS.n1621 AVSS.n1599 9.3005
R9793 AVSS.n1621 AVSS.n1598 9.3005
R9794 AVSS.n1621 AVSS.n1600 9.3005
R9795 AVSS.n1621 AVSS.n1597 9.3005
R9796 AVSS.n1621 AVSS.n1620 9.3005
R9797 AVSS.n1619 AVSS.n1599 9.3005
R9798 AVSS.n1619 AVSS.n1598 9.3005
R9799 AVSS.n1619 AVSS.n1600 9.3005
R9800 AVSS.n1619 AVSS.n1597 9.3005
R9801 AVSS.n1620 AVSS.n1619 9.3005
R9802 AVSS.n3405 AVSS.n3399 9.3005
R9803 AVSS.n3405 AVSS.n3398 9.3005
R9804 AVSS.n3405 AVSS.n3402 9.3005
R9805 AVSS.n3417 AVSS.n3405 9.3005
R9806 AVSS.n3407 AVSS.n3399 9.3005
R9807 AVSS.n3407 AVSS.n3398 9.3005
R9808 AVSS.n3407 AVSS.n3402 9.3005
R9809 AVSS.n3417 AVSS.n3407 9.3005
R9810 AVSS.n3404 AVSS.n3399 9.3005
R9811 AVSS.n3404 AVSS.n3398 9.3005
R9812 AVSS.n3404 AVSS.n3402 9.3005
R9813 AVSS.n3417 AVSS.n3404 9.3005
R9814 AVSS.n3409 AVSS.n3399 9.3005
R9815 AVSS.n3409 AVSS.n3398 9.3005
R9816 AVSS.n3409 AVSS.n3402 9.3005
R9817 AVSS.n3417 AVSS.n3409 9.3005
R9818 AVSS.n3418 AVSS.n3399 9.3005
R9819 AVSS.n3418 AVSS.n3398 9.3005
R9820 AVSS.n3418 AVSS.n3402 9.3005
R9821 AVSS.n3418 AVSS.n3397 9.3005
R9822 AVSS.n3418 AVSS.n3417 9.3005
R9823 AVSS.n3416 AVSS.n3399 9.3005
R9824 AVSS.n3416 AVSS.n3398 9.3005
R9825 AVSS.n3416 AVSS.n3402 9.3005
R9826 AVSS.n3416 AVSS.n3397 9.3005
R9827 AVSS.n3417 AVSS.n3416 9.3005
R9828 AVSS.n3670 AVSS.n3669 9.3005
R9829 AVSS.n3660 AVSS.n3653 9.3005
R9830 AVSS.n3667 AVSS.n3660 9.3005
R9831 AVSS.n3667 AVSS.n3666 9.3005
R9832 AVSS.n3660 AVSS.n3658 9.3005
R9833 AVSS.n3666 AVSS.n3658 9.3005
R9834 AVSS.n3669 AVSS.n3656 9.3005
R9835 AVSS.n3666 AVSS.n3656 9.3005
R9836 AVSS.n3666 AVSS.n3662 9.3005
R9837 AVSS.n3665 AVSS.n3660 9.3005
R9838 AVSS.n3666 AVSS.n3665 9.3005
R9839 AVSS.n3673 AVSS.n3647 9.3005
R9840 AVSS.n3652 AVSS.n3642 9.3005
R9841 AVSS.n3673 AVSS.n3652 9.3005
R9842 AVSS.n3646 AVSS.n3643 9.3005
R9843 AVSS.n3673 AVSS.n3646 9.3005
R9844 AVSS.n3643 AVSS.n3641 9.3005
R9845 AVSS.n3673 AVSS.n3641 9.3005
R9846 AVSS.n3674 AVSS.n3643 9.3005
R9847 AVSS.n3674 AVSS.n3642 9.3005
R9848 AVSS.n3674 AVSS.n3673 9.3005
R9849 AVSS.n3672 AVSS.n3643 9.3005
R9850 AVSS.n3673 AVSS.n3672 9.3005
R9851 AVSS.n3851 AVSS.n3677 9.3005
R9852 AVSS.n3870 AVSS.n3869 9.3005
R9853 AVSS.n4062 AVSS.n3888 9.3005
R9854 AVSS.n4081 AVSS.n4080 9.3005
R9855 AVSS.n4205 AVSS.n4204 9.3005
R9856 AVSS.n4136 AVSS.n231 9.3005
R9857 AVSS.n147 AVSS.n146 9.3005
R9858 AVSS.n4334 AVSS.n4333 9.3005
R9859 AVSS.n4331 AVSS.n4330 9.3005
R9860 AVSS.n4301 AVSS.n4300 9.3005
R9861 AVSS.n4298 AVSS.n4297 9.3005
R9862 AVSS.n4268 AVSS.n4267 9.3005
R9863 AVSS.n4265 AVSS.n4264 9.3005
R9864 AVSS.n6086 AVSS.n6085 9.3005
R9865 AVSS.n262 AVSS.n261 9.3005
R9866 AVSS.n276 AVSS.n270 9.3005
R9867 AVSS.n276 AVSS.n273 9.3005
R9868 AVSS.n6080 AVSS.n276 9.3005
R9869 AVSS.n6077 AVSS.n270 9.3005
R9870 AVSS.n6077 AVSS.n273 9.3005
R9871 AVSS.n6077 AVSS.n265 9.3005
R9872 AVSS.n6080 AVSS.n6077 9.3005
R9873 AVSS.n275 AVSS.n270 9.3005
R9874 AVSS.n275 AVSS.n266 9.3005
R9875 AVSS.n275 AVSS.n273 9.3005
R9876 AVSS.n6080 AVSS.n275 9.3005
R9877 AVSS.n270 AVSS.n264 9.3005
R9878 AVSS.n266 AVSS.n264 9.3005
R9879 AVSS.n273 AVSS.n264 9.3005
R9880 AVSS.n6080 AVSS.n264 9.3005
R9881 AVSS.n6081 AVSS.n270 9.3005
R9882 AVSS.n6081 AVSS.n266 9.3005
R9883 AVSS.n6081 AVSS.n273 9.3005
R9884 AVSS.n6081 AVSS.n265 9.3005
R9885 AVSS.n6081 AVSS.n6080 9.3005
R9886 AVSS.n6079 AVSS.n270 9.3005
R9887 AVSS.n6079 AVSS.n266 9.3005
R9888 AVSS.n6079 AVSS.n273 9.3005
R9889 AVSS.n6080 AVSS.n6079 9.3005
R9890 AVSS.n6025 AVSS.n6006 9.10376
R9891 AVSS.n6010 AVSS.n6006 9.10376
R9892 AVSS.n5983 AVSS.n5982 8.86463
R9893 AVSS.n1294 AVSS.n1293 8.53383
R9894 AVSS.n1173 AVSS.n1147 8.53383
R9895 AVSS.n4981 AVSS.n1068 8.53383
R9896 AVSS.n4667 AVSS.n4648 8.53383
R9897 AVSS.n5725 AVSS.n5629 8.53383
R9898 AVSS.n834 AVSS.n683 8.53383
R9899 AVSS.n737 AVSS.n716 8.53383
R9900 AVSS.n4986 AVSS.n4985 8.53383
R9901 AVSS.n3218 AVSS.n3217 8.53383
R9902 AVSS.n3097 AVSS.n3072 8.53383
R9903 AVSS.n4672 AVSS.n4671 8.53383
R9904 AVSS.n2512 AVSS.n2511 8.53383
R9905 AVSS.n1845 AVSS.n1844 8.53383
R9906 AVSS.n6210 AVSS.n148 8.53383
R9907 AVSS.n6009 AVSS.n6005 7.86463
R9908 AVSS.n5817 AVSS.n5727 7.46717
R9909 AVSS.n5545 AVSS.n5455 7.46717
R9910 AVSS.n5374 AVSS.n5373 7.46717
R9911 AVSS.n5175 AVSS.n5174 7.46717
R9912 AVSS.n3160 AVSS.n3159 7.46717
R9913 AVSS.n1236 AVSS.n1235 7.46717
R9914 AVSS.n4615 AVSS.n4524 7.46717
R9915 AVSS.n777 AVSS.n776 7.46717
R9916 AVSS.n1065 AVSS.n975 7.46717
R9917 AVSS.n2508 AVSS.n2417 7.46717
R9918 AVSS.n2541 AVSS.n2540 7.46717
R9919 AVSS.n4341 AVSS.n3511 7.3702
R9920 AVSS.n2189 AVSS.n2069 7.2409
R9921 AVSS.n2157 AVSS.n2081 7.2409
R9922 AVSS.n376 AVSS.n326 7.2409
R9923 AVSS.n1558 AVSS.n1483 7.2409
R9924 AVSS.n1593 AVSS.n1383 7.2409
R9925 AVSS.n945 AVSS.n646 7.2409
R9926 AVSS.n4720 AVSS.n1716 7.2409
R9927 AVSS.n4903 AVSS.n1381 7.2409
R9928 AVSS.n4807 AVSS.n4806 7.2409
R9929 AVSS.n1861 AVSS.n1858 7.2409
R9930 AVSS.n2589 AVSS.n1739 7.2409
R9931 AVSS.n4414 AVSS.n4413 7.2409
R9932 AVSS.n4448 AVSS.n4345 7.2409
R9933 AVSS.n6023 AVSS.n6022 6.96479
R9934 AVSS.n6022 AVSS.n6021 6.96479
R9935 AVSS.n6015 AVSS.n6007 6.96479
R9936 AVSS.n6016 AVSS.n6015 6.96479
R9937 AVSS.n5960 AVSS.n5942 6.85408
R9938 AVSS.n6044 AVSS.n5934 6.85104
R9939 AVSS.n5548 AVSS.n5257 6.72373
R9940 AVSS.n5419 AVSS.n5395 6.72373
R9941 AVSS.n6302 AVSS.n6301 6.72373
R9942 AVSS.n5196 AVSS.n409 6.72373
R9943 AVSS.n5099 AVSS.n408 6.72373
R9944 AVSS.n5878 AVSS.n325 6.72373
R9945 AVSS.n5820 AVSS.n5626 6.72373
R9946 AVSS.n2301 AVSS.n973 6.72373
R9947 AVSS.n2414 AVSS.n2413 6.72373
R9948 AVSS.n2342 AVSS.n2341 6.72373
R9949 AVSS.n4993 AVSS.n645 6.72373
R9950 AVSS.n2585 AVSS.n1740 6.72373
R9951 AVSS.n2538 AVSS.n2537 6.72373
R9952 AVSS.n4678 AVSS.n2776 6.20656
R9953 AVSS.n4682 AVSS.n4681 6.20656
R9954 AVSS.n4710 AVSS.n1723 6.20656
R9955 AVSS.n4714 AVSS.n4713 6.20656
R9956 AVSS.n2562 AVSS.n1747 6.20656
R9957 AVSS.n2514 AVSS.n2513 6.20656
R9958 AVSS.n261 AVSS.n232 6.20656
R9959 AVSS.n4269 AVSS.n4268 6.20656
R9960 AVSS.n4297 AVSS.n3889 6.20656
R9961 AVSS.n4302 AVSS.n4301 6.20656
R9962 AVSS.n4330 AVSS.n3678 6.20656
R9963 AVSS.n4335 AVSS.n4334 6.20656
R9964 AVSS.n4264 AVSS.n4206 6.20656
R9965 AVSS.n6087 AVSS.n6086 6.20656
R9966 AVSS.n6027 AVSS.n6025 6.06843
R9967 AVSS.n6050 AVSS.n6047 5.4543
R9968 AVSS.n6050 AVSS.n6049 5.4543
R9969 AVSS.n6042 AVSS.n6041 5.4543
R9970 AVSS.n4678 AVSS.n4677 5.4308
R9971 AVSS.n4681 AVSS.n1737 5.4308
R9972 AVSS.n4710 AVSS.n4709 5.4308
R9973 AVSS.n4713 AVSS.n1721 5.4308
R9974 AVSS.n2563 AVSS.n2562 5.4308
R9975 AVSS.n2513 AVSS.n1852 5.4308
R9976 AVSS.n261 AVSS.n260 5.4308
R9977 AVSS.n4268 AVSS.n3989 5.4308
R9978 AVSS.n4297 AVSS.n4296 5.4308
R9979 AVSS.n4301 AVSS.n3778 5.4308
R9980 AVSS.n4330 AVSS.n4329 5.4308
R9981 AVSS.n4334 AVSS.n3640 5.4308
R9982 AVSS.n4264 AVSS.n4263 5.4308
R9983 AVSS.n6086 AVSS.n228 5.4308
R9984 AVSS.t27 AVSS.t22 5.04521
R9985 AVSS.n5549 AVSS.n5548 4.91363
R9986 AVSS.n5395 AVSS.n5299 4.91363
R9987 AVSS.n6302 AVSS.n2 4.91363
R9988 AVSS.n5197 AVSS.n5196 4.91363
R9989 AVSS.n5099 AVSS.n5098 4.91363
R9990 AVSS.n325 AVSS.n322 4.91363
R9991 AVSS.n5821 AVSS.n5820 4.91363
R9992 AVSS.n2301 AVSS.n2300 4.91363
R9993 AVSS.n2414 AVSS.n2303 4.91363
R9994 AVSS.n2343 AVSS.n2342 4.91363
R9995 AVSS.n645 AVSS.n642 4.91363
R9996 AVSS.n2578 AVSS.n1740 4.91363
R9997 AVSS.n2538 AVSS.n1824 4.91363
R9998 AVSS.n565 AVSS.n556 4.64589
R9999 AVSS.n5022 AVSS.n568 4.64589
R10000 AVSS.n567 AVSS.n556 4.64589
R10001 AVSS.n5023 AVSS.n5022 4.64589
R10002 AVSS.n5022 AVSS.n558 4.64589
R10003 AVSS.n1606 AVSS.n1597 4.64589
R10004 AVSS.n1617 AVSS.n1611 4.64589
R10005 AVSS.n1608 AVSS.n1597 4.64589
R10006 AVSS.n1617 AVSS.n1596 4.64589
R10007 AVSS.n1618 AVSS.n1617 4.64589
R10008 AVSS.n3406 AVSS.n3397 4.64589
R10009 AVSS.n3414 AVSS.n3410 4.64589
R10010 AVSS.n3408 AVSS.n3397 4.64589
R10011 AVSS.n3414 AVSS.n3396 4.64589
R10012 AVSS.n3415 AVSS.n3414 4.64589
R10013 AVSS.n6078 AVSS.n265 4.64429
R10014 AVSS.n278 AVSS.n266 4.64429
R10015 AVSS.n274 AVSS.n265 4.64429
R10016 AVSS.n580 AVSS.n578 4.64414
R10017 AVSS.n580 AVSS.n579 4.64414
R10018 AVSS.n584 AVSS.n582 4.64414
R10019 AVSS.n585 AVSS.n584 4.64414
R10020 AVSS.n1101 AVSS.n1099 4.64414
R10021 AVSS.n1101 AVSS.n1100 4.64414
R10022 AVSS.n1105 AVSS.n1103 4.64414
R10023 AVSS.n1106 AVSS.n1105 4.64414
R10024 AVSS.n4486 AVSS.n4484 4.64414
R10025 AVSS.n4486 AVSS.n4485 4.64414
R10026 AVSS.n4490 AVSS.n4488 4.64414
R10027 AVSS.n4491 AVSS.n4490 4.64414
R10028 AVSS.n3651 AVSS.n3643 4.64199
R10029 AVSS.n3671 AVSS.n3642 4.64199
R10030 AVSS.n3645 AVSS.n3642 4.64199
R10031 AVSS.n3669 AVSS.n3668 4.63919
R10032 AVSS.n3661 AVSS.n3660 4.63919
R10033 AVSS.n3669 AVSS.n3655 4.63919
R10034 AVSS.n5939 AVSS.n5937 4.53538
R10035 AVSS.n6013 AVSS.n5939 4.53538
R10036 AVSS.n5938 AVSS.n5936 4.53538
R10037 AVSS.n5999 AVSS.n5938 4.53538
R10038 AVSS.n2189 AVSS.n2188 4.39646
R10039 AVSS.n2160 AVSS.n2081 4.39646
R10040 AVSS.n5876 AVSS.n326 4.39646
R10041 AVSS.n1561 AVSS.n1483 4.39646
R10042 AVSS.n1593 AVSS.n1592 4.39646
R10043 AVSS.n4991 AVSS.n646 4.39646
R10044 AVSS.n4720 AVSS.n4719 4.39646
R10045 AVSS.n4904 AVSS.n4903 4.39646
R10046 AVSS.n4807 AVSS.n1371 4.39646
R10047 AVSS.n1863 AVSS.n1861 4.39646
R10048 AVSS.n2589 AVSS.n2588 4.39646
R10049 AVSS.n4415 AVSS.n4414 4.39646
R10050 AVSS.n4445 AVSS.n4345 4.39646
R10051 AVSS.n4341 AVSS.n4340 4.26717
R10052 AVSS.n6031 AVSS.n6030 4.14168
R10053 AVSS.n6037 AVSS.n6036 4.14168
R10054 AVSS.n5998 AVSS 4.03627
R10055 AVSS.n4152 AVSS.n4136 3.91161
R10056 AVSS.n4080 AVSS.n3990 3.91161
R10057 AVSS.n3869 AVSS.n3779 3.91161
R10058 AVSS.n3509 AVSS.n3420 3.91161
R10059 AVSS.n1480 AVSS.n1390 3.91161
R10060 AVSS.n4900 AVSS.n4810 3.91161
R10061 AVSS.n2682 AVSS.n2592 3.91161
R10062 AVSS.n1714 AVSS.n1625 3.91161
R10063 AVSS.n2560 AVSS.n1750 3.91161
R10064 AVSS.n2067 AVSS.n1977 3.91161
R10065 AVSS.n3343 AVSS.n3342 3.91161
R10066 AVSS.n5029 AVSS.n461 3.14302
R10067 AVSS.n6229 AVSS.n6228 3.14287
R10068 AVSS.n6241 AVSS.n6240 3.14018
R10069 AVSS.n5041 AVSS.n453 3.14006
R10070 AVSS.n5029 AVSS.n5028 3.11197
R10071 AVSS.n6229 AVSS.n6226 3.10645
R10072 AVSS.n1293 AVSS.n1164 3.10353
R10073 AVSS.n1366 AVSS.n1147 3.10353
R10074 AVSS.n4981 AVSS.n4980 3.10353
R10075 AVSS.n4667 AVSS.n4666 3.10353
R10076 AVSS.n5725 AVSS.n5724 3.10353
R10077 AVSS.n835 AVSS.n834 3.10353
R10078 AVSS.n737 AVSS.n736 3.10353
R10079 AVSS.n4985 AVSS.n974 3.10353
R10080 AVSS.n3217 AVSS.n3090 3.10353
R10081 AVSS.n3291 AVSS.n3072 3.10353
R10082 AVSS.n4671 AVSS.n4523 3.10353
R10083 AVSS.n2511 AVSS.n1885 3.10353
R10084 AVSS.n1844 AVSS.n1843 3.10353
R10085 AVSS.n6210 AVSS.n6209 3.10353
R10086 AVSS.n6231 AVSS.n6228 3.1005
R10087 AVSS.n6234 AVSS.n39 3.1005
R10088 AVSS.n40 AVSS.n35 3.1005
R10089 AVSS.n6239 AVSS.n32 3.1005
R10090 AVSS.n6242 AVSS.n6241 3.1005
R10091 AVSS.n6232 AVSS.n6231 3.1005
R10092 AVSS.n6234 AVSS.n6233 3.1005
R10093 AVSS.n35 AVSS.n34 3.1005
R10094 AVSS.n6240 AVSS.n6239 3.1005
R10095 AVSS.n5042 AVSS.n5041 3.1005
R10096 AVSS.n5039 AVSS.n452 3.1005
R10097 AVSS.n5037 AVSS.n457 3.1005
R10098 AVSS.n5033 AVSS.n458 3.1005
R10099 AVSS.n461 AVSS.n460 3.1005
R10100 AVSS.n5039 AVSS.n453 3.1005
R10101 AVSS.n5037 AVSS.n5036 3.1005
R10102 AVSS.n5034 AVSS.n5033 3.1005
R10103 AVSS.n460 AVSS.n459 3.1005
R10104 AVSS.n6216 AVSS.n51 3.06583
R10105 AVSS.n6214 AVSS.n51 3.06583
R10106 AVSS.n6220 AVSS.n47 3.06583
R10107 AVSS.n6218 AVSS.n47 3.06583
R10108 AVSS.n6224 AVSS.n43 3.06583
R10109 AVSS.n6222 AVSS.n43 3.06583
R10110 AVSS AVSS.n112 3.02272
R10111 AVSS.n4161 AVSS 3.02272
R10112 AVSS AVSS.n4020 3.02272
R10113 AVSS AVSS.n3809 3.02272
R10114 AVSS AVSS.n3450 3.02272
R10115 AVSS.n5767 AVSS 3.02272
R10116 AVSS.n5495 AVSS 3.02272
R10117 AVSS.n5327 AVSS 3.02272
R10118 AVSS.n5128 AVSS 3.02272
R10119 AVSS.n490 AVSS 3.02272
R10120 AVSS.n1451 AVSS 3.02272
R10121 AVSS.n4871 AVSS 3.02272
R10122 AVSS AVSS.n3186 3.02272
R10123 AVSS AVSS.n1262 3.02272
R10124 AVSS.n4564 AVSS 3.02272
R10125 AVSS AVSS.n2740 3.02272
R10126 AVSS AVSS.n2622 3.02272
R10127 AVSS AVSS.n1655 3.02272
R10128 AVSS AVSS.n1798 3.02272
R10129 AVSS.n2038 AVSS 3.02272
R10130 AVSS AVSS.n803 3.02272
R10131 AVSS.n1015 AVSS 3.02272
R10132 AVSS.n2460 AVSS 3.02272
R10133 AVSS.n1914 AVSS 3.02272
R10134 AVSS.n3332 AVSS 3.02272
R10135 AVSS.n6045 AVSS.n6044 2.85104
R10136 AVSS.n6043 AVSS.n6039 2.84833
R10137 AVSS.n5997 AVSS.n5996 2.54398
R10138 AVSS.n5998 AVSS.n5997 2.54398
R10139 AVSS.n5994 AVSS.n5993 2.54398
R10140 AVSS.n5993 AVSS.n5992 2.54398
R10141 AVSS.n3876 AVSS.n3875 2.36206
R10142 AVSS.n4087 AVSS.n4086 2.36206
R10143 AVSS.n4112 AVSS.n4111 2.36206
R10144 AVSS.n6255 AVSS.n6254 2.36206
R10145 AVSS.n5054 AVSS.n5053 2.36206
R10146 AVSS.n5045 AVSS.n5044 2.36206
R10147 AVSS.n6061 AVSS.n290 2.24235
R10148 AVSS.n5982 AVSS.n5977 2.24235
R10149 AVSS.n5955 AVSS.n5953 2.22061
R10150 AVSS.n5956 AVSS.n5955 2.22061
R10151 AVSS.n5956 AVSS.n5946 2.22061
R10152 AVSS.n5953 AVSS.n5946 2.22061
R10153 AVSS.n3886 AVSS.n3885 2.19742
R10154 AVSS.n4097 AVSS.n4096 2.19742
R10155 AVSS.n4102 AVSS.n263 2.19742
R10156 AVSS.n6245 AVSS.n6244 2.19742
R10157 AVSS.n6259 AVSS.n6257 2.19742
R10158 AVSS.n5058 AVSS.n5056 2.19742
R10159 AVSS.n6039 AVSS.n6038 2.19615
R10160 AVSS.n269 AVSS.n54 2.18373
R10161 AVSS.n6062 AVSS.n6061 2.17441
R10162 AVSS.n5974 AVSS.n5973 1.9842
R10163 AVSS.n5972 AVSS.n5970 1.9842
R10164 AVSS.n5975 AVSS.n5974 1.94072
R10165 AVSS.n5972 AVSS.n5971 1.94072
R10166 AVSS.n5954 AVSS.n5948 1.88285
R10167 AVSS.n294 AVSS.n292 1.84012
R10168 AVSS.n293 AVSS.n291 1.84012
R10169 AVSS.n285 AVSS.n279 1.78458
R10170 AVSS.n286 AVSS.n285 1.77229
R10171 AVSS.n6068 AVSS.n279 1.64097
R10172 AVSS.n4101 AVSS.n4100 1.5505
R10173 AVSS.n4106 AVSS.n4105 1.5505
R10174 AVSS.n4108 AVSS.n4107 1.5505
R10175 AVSS.n4110 AVSS.n4098 1.5505
R10176 AVSS.n4095 AVSS.n4082 1.5505
R10177 AVSS.n4093 AVSS.n4092 1.5505
R10178 AVSS.n4091 AVSS.n4090 1.5505
R10179 AVSS.n4088 AVSS.n4085 1.5505
R10180 AVSS.n3884 AVSS.n3871 1.5505
R10181 AVSS.n3882 AVSS.n3881 1.5505
R10182 AVSS.n3880 AVSS.n3879 1.5505
R10183 AVSS.n3877 AVSS.n3874 1.5505
R10184 AVSS.n5060 AVSS.n5059 1.5505
R10185 AVSS.n5062 AVSS.n5061 1.5505
R10186 AVSS.n5049 AVSS.n451 1.5505
R10187 AVSS.n5048 AVSS.n5047 1.5505
R10188 AVSS.n6261 AVSS.n6260 1.5505
R10189 AVSS.n6263 AVSS.n6262 1.5505
R10190 AVSS.n23 AVSS.n22 1.5505
R10191 AVSS.n5052 AVSS.n5050 1.5505
R10192 AVSS.n29 AVSS.n28 1.5505
R10193 AVSS.n6249 AVSS.n6248 1.5505
R10194 AVSS.n6251 AVSS.n6250 1.5505
R10195 AVSS.n6253 AVSS.n25 1.5505
R10196 AVSS.n6221 AVSS.n46 1.54998
R10197 AVSS.n6217 AVSS.n50 1.54998
R10198 AVSS.n6213 AVSS.n6212 1.54998
R10199 AVSS.n5987 AVSS.n5965 1.52394
R10200 AVSS.n5991 AVSS.n5965 1.52394
R10201 AVSS.n5990 AVSS.n5989 1.52394
R10202 AVSS.n5991 AVSS.n5990 1.52394
R10203 AVSS.n6075 AVSS.t68 1.50457
R10204 AVSS.n5546 AVSS.n31 1.45331
R10205 AVSS.n4723 AVSS.n1622 1.42498
R10206 AVSS.n1610 AVSS.n1595 1.42498
R10207 AVSS.n5027 AVSS.n555 1.42498
R10208 AVSS.n4343 AVSS.n3419 1.42498
R10209 AVSS.n4266 AVSS.n4113 1.42238
R10210 AVSS.n4299 AVSS.n3887 1.42238
R10211 AVSS.n6225 AVSS.n42 1.42238
R10212 AVSS.n4332 AVSS.n3676 1.42238
R10213 AVSS.n6084 AVSS.n6083 1.42238
R10214 AVSS.n5055 AVSS.n0 1.41977
R10215 AVSS.n6256 AVSS.n24 1.41977
R10216 AVSS.n6243 AVSS.n31 1.41977
R10217 AVSS.n5043 AVSS.n420 1.41977
R10218 AVSS.n2561 AVSS.n1749 1.3249
R10219 AVSS.n2539 AVSS.n1738 1.3249
R10220 AVSS.n1333 AVSS 1.29343
R10221 AVSS AVSS.n1084 1.29343
R10222 AVSS.n2173 AVSS 1.29343
R10223 AVSS.n5601 AVSS 1.29343
R10224 AVSS AVSS.n5297 1.29343
R10225 AVSS.n5204 AVSS 1.29343
R10226 AVSS AVSS.n319 1.29343
R10227 AVSS.n5688 AVSS 1.29343
R10228 AVSS AVSS.n873 1.29343
R10229 AVSS.n2241 AVSS 1.29343
R10230 AVSS.n2401 AVSS 1.29343
R10231 AVSS.n1576 AVSS 1.29343
R10232 AVSS AVSS.n639 1.29343
R10233 AVSS.n3257 AVSS 1.29343
R10234 AVSS AVSS.n2889 1.29343
R10235 AVSS.n3028 AVSS 1.29343
R10236 AVSS AVSS.n2819 1.29343
R10237 AVSS AVSS.n4921 1.29343
R10238 AVSS AVSS.n2574 1.29343
R10239 AVSS.n6174 AVSS 1.29343
R10240 AVSS AVSS.n3904 1.29343
R10241 AVSS AVSS.n3693 1.29343
R10242 AVSS AVSS.n3517 1.29343
R10243 AVSS AVSS.n6101 1.29343
R10244 AVSS.n4431 AVSS 1.29343
R10245 AVSS.n3878 AVSS.n3877 1.25468
R10246 AVSS.n4089 AVSS.n4088 1.25468
R10247 AVSS.n4110 AVSS.n4109 1.25468
R10248 AVSS.n3660 AVSS.n3654 1.25468
R10249 AVSS.n3400 AVSS.n3397 1.25468
R10250 AVSS.n1601 AVSS.n1597 1.25468
R10251 AVSS.n569 AVSS.n556 1.25468
R10252 AVSS.n5032 AVSS.n460 1.25468
R10253 AVSS.n580 AVSS.n577 1.25468
R10254 AVSS.n1101 AVSS.n1098 1.25468
R10255 AVSS.n4486 AVSS.n4483 1.25468
R10256 AVSS.n6239 AVSS.n6238 1.25468
R10257 AVSS.n6253 AVSS.n6252 1.25468
R10258 AVSS.n5052 AVSS.n5051 1.25468
R10259 AVSS.n5047 AVSS.n5046 1.25468
R10260 AVSS.n271 AVSS.n265 1.25468
R10261 AVSS.n6010 AVSS.n6009 1.23963
R10262 AVSS.n2561 AVSS.n1738 1.1999
R10263 AVSS.n2539 AVSS.n1749 1.1999
R10264 AVSS.n3885 AVSS.n3884 1.19225
R10265 AVSS.n4096 AVSS.n4095 1.19225
R10266 AVSS.n4102 AVSS.n4101 1.19225
R10267 AVSS.n3648 AVSS.n3642 1.19225
R10268 AVSS.n3413 AVSS.n3399 1.19225
R10269 AVSS.n1616 AVSS.n1599 1.19225
R10270 AVSS.n5021 AVSS.n559 1.19225
R10271 AVSS.n5040 AVSS.n5039 1.19225
R10272 AVSS.n584 AVSS.n583 1.19225
R10273 AVSS.n1105 AVSS.n1104 1.19225
R10274 AVSS.n4490 AVSS.n4489 1.19225
R10275 AVSS.n6231 AVSS.n6230 1.19225
R10276 AVSS.n6245 AVSS.n29 1.19225
R10277 AVSS.n6260 AVSS.n6259 1.19225
R10278 AVSS.n5059 AVSS.n5058 1.19225
R10279 AVSS.n270 AVSS.n269 1.19225
R10280 AVSS.n2509 AVSS.n2416 1.15935
R10281 AVSS.n2068 AVSS.n1976 1.15935
R10282 AVSS.n4616 AVSS.n1067 1.15935
R10283 AVSS.n2591 AVSS.n1722 1.15805
R10284 AVSS.n6027 AVSS.n6026 1.1418
R10285 AVSS.n832 AVSS.n739 1.1357
R10286 AVSS.n1291 AVSS.n1198 1.1357
R10287 AVSS.n3215 AVSS.n3122 1.1357
R10288 AVSS.n1481 AVSS.n1382 1.1357
R10289 AVSS.n4901 AVSS.n4809 1.1357
R10290 AVSS.n3395 AVSS.n3303 1.1357
R10291 AVSS.n5194 AVSS.n5101 1.1357
R10292 AVSS.n5393 AVSS.n1 1.1357
R10293 AVSS.n3870 AVSS.n3677 1.1357
R10294 AVSS.n4081 AVSS.n3888 1.1357
R10295 AVSS.n4205 AVSS.n231 1.1357
R10296 AVSS AVSS.n6063 1.07226
R10297 AVSS.n3879 AVSS.n3873 1.07024
R10298 AVSS.n4090 AVSS.n4084 1.07024
R10299 AVSS.n4108 AVSS.n4099 1.07024
R10300 AVSS.n3669 AVSS.n3644 1.07024
R10301 AVSS.n3402 AVSS.n3401 1.07024
R10302 AVSS.n1612 AVSS.n1600 1.07024
R10303 AVSS.n5017 AVSS.n560 1.07024
R10304 AVSS.n5033 AVSS.n456 1.07024
R10305 AVSS.n590 AVSS.n573 1.07024
R10306 AVSS.n1111 AVSS.n1094 1.07024
R10307 AVSS.n4496 AVSS.n4479 1.07024
R10308 AVSS.n6235 AVSS.n35 1.07024
R10309 AVSS.n6251 AVSS.n27 1.07024
R10310 AVSS.n6264 AVSS.n22 1.07024
R10311 AVSS.n5063 AVSS.n451 1.07024
R10312 AVSS.n273 AVSS.n272 1.07024
R10313 AVSS.n6046 AVSS.n6045 1.06028
R10314 AVSS.n6047 AVSS.n6046 1.06028
R10315 AVSS.n3877 AVSS.n3876 1.0237
R10316 AVSS.n4088 AVSS.n4087 1.0237
R10317 AVSS.n4111 AVSS.n4110 1.0237
R10318 AVSS.n3664 AVSS.n3660 1.0237
R10319 AVSS.n3403 AVSS.n3397 1.0237
R10320 AVSS.n1603 AVSS.n1597 1.0237
R10321 AVSS.n561 AVSS.n556 1.0237
R10322 AVSS.n5030 AVSS.n460 1.0237
R10323 AVSS.n586 AVSS.n580 1.0237
R10324 AVSS.n1107 AVSS.n1101 1.0237
R10325 AVSS.n4492 AVSS.n4486 1.0237
R10326 AVSS.n6239 AVSS.n33 1.0237
R10327 AVSS.n6254 AVSS.n6253 1.0237
R10328 AVSS.n5053 AVSS.n5052 1.0237
R10329 AVSS.n5047 AVSS.n5045 1.0237
R10330 AVSS.n277 AVSS.n265 1.0237
R10331 AVSS.n3884 AVSS.n3883 0.959578
R10332 AVSS.n4095 AVSS.n4094 0.959578
R10333 AVSS.n4104 AVSS.n4101 0.959578
R10334 AVSS.n3650 AVSS.n3642 0.959578
R10335 AVSS.n3411 AVSS.n3399 0.959578
R10336 AVSS.n1614 AVSS.n1599 0.959578
R10337 AVSS.n5019 AVSS.n559 0.959578
R10338 AVSS.n5039 AVSS.n5038 0.959578
R10339 AVSS.n584 AVSS.n581 0.959578
R10340 AVSS.n1105 AVSS.n1102 0.959578
R10341 AVSS.n4490 AVSS.n4487 0.959578
R10342 AVSS.n6231 AVSS.n6227 0.959578
R10343 AVSS.n6247 AVSS.n29 0.959578
R10344 AVSS.n6260 AVSS.n6258 0.959578
R10345 AVSS.n5059 AVSS.n5057 0.959578
R10346 AVSS.n270 AVSS.n267 0.959578
R10347 AVSS.n6003 AVSS.n6002 0.878527
R10348 AVSS.n6001 AVSS.n6000 0.878527
R10349 AVSS.n5955 AVSS.n5954 0.845955
R10350 AVSS.n5958 AVSS.n5946 0.845955
R10351 AVSS.n5952 AVSS.n5950 0.842891
R10352 AVSS.n5985 AVSS.n289 0.839004
R10353 AVSS.n3666 AVSS.n3664 0.812055
R10354 AVSS.n6080 AVSS.n277 0.812055
R10355 AVSS.n3417 AVSS.n3403 0.812055
R10356 AVSS.n1620 AVSS.n1603 0.812055
R10357 AVSS.n5025 AVSS.n561 0.812055
R10358 AVSS.n5030 AVSS.n5029 0.812055
R10359 AVSS.n587 AVSS.n586 0.812055
R10360 AVSS.n1108 AVSS.n1107 0.812055
R10361 AVSS.n4493 AVSS.n4492 0.812055
R10362 AVSS.n6241 AVSS.n33 0.812055
R10363 AVSS.n6049 AVSS.n6048 0.792006
R10364 AVSS.n6041 AVSS.n6040 0.792006
R10365 AVSS.n3882 AVSS.n3873 0.77514
R10366 AVSS.n4093 AVSS.n4084 0.77514
R10367 AVSS.n4105 AVSS.n4099 0.77514
R10368 AVSS.n3673 AVSS.n3644 0.77514
R10369 AVSS.n3401 AVSS.n3398 0.77514
R10370 AVSS.n1612 AVSS.n1598 0.77514
R10371 AVSS.n5017 AVSS.n557 0.77514
R10372 AVSS.n5037 AVSS.n456 0.77514
R10373 AVSS.n590 AVSS.n589 0.77514
R10374 AVSS.n1111 AVSS.n1110 0.77514
R10375 AVSS.n4496 AVSS.n4495 0.77514
R10376 AVSS.n6235 AVSS.n6234 0.77514
R10377 AVSS.n6248 AVSS.n27 0.77514
R10378 AVSS.n6264 AVSS.n6263 0.77514
R10379 AVSS.n5063 AVSS.n5062 0.77514
R10380 AVSS.n272 AVSS.n266 0.77514
R10381 AVSS.n5953 AVSS.n5945 0.715885
R10382 AVSS.n5957 AVSS.n5956 0.715885
R10383 AVSS.n6025 AVSS.n6024 0.715885
R10384 AVSS.n6011 AVSS.n6010 0.715885
R10385 AVSS.n6044 AVSS.n6043 0.710007
R10386 AVSS.n3648 AVSS.n3643 0.647417
R10387 AVSS.n3414 AVSS.n3413 0.647417
R10388 AVSS.n1617 AVSS.n1616 0.647417
R10389 AVSS.n5022 AVSS.n5021 0.647417
R10390 AVSS.n5041 AVSS.n5040 0.647417
R10391 AVSS.n583 AVSS.n43 0.647417
R10392 AVSS.n1104 AVSS.n47 0.647417
R10393 AVSS.n4489 AVSS.n51 0.647417
R10394 AVSS.n6230 AVSS.n6229 0.647417
R10395 AVSS.n6046 AVSS.n5933 0.6205
R10396 AVSS.n6052 AVSS.n5932 0.6205
R10397 AVSS.n3879 AVSS.n3878 0.590702
R10398 AVSS.n4090 AVSS.n4089 0.590702
R10399 AVSS.n4109 AVSS.n4108 0.590702
R10400 AVSS.n3669 AVSS.n3654 0.590702
R10401 AVSS.n3402 AVSS.n3400 0.590702
R10402 AVSS.n1601 AVSS.n1600 0.590702
R10403 AVSS.n569 AVSS.n560 0.590702
R10404 AVSS.n5033 AVSS.n5032 0.590702
R10405 AVSS.n577 AVSS.n573 0.590702
R10406 AVSS.n1098 AVSS.n1094 0.590702
R10407 AVSS.n4483 AVSS.n4479 0.590702
R10408 AVSS.n6238 AVSS.n35 0.590702
R10409 AVSS.n6252 AVSS.n6251 0.590702
R10410 AVSS.n5051 AVSS.n22 0.590702
R10411 AVSS.n5046 AVSS.n451 0.590702
R10412 AVSS.n273 AVSS.n271 0.590702
R10413 AVSS.n6004 AVSS.n6003 0.590174
R10414 AVSS.n6000 AVSS.n5934 0.590174
R10415 AVSS.n5956 AVSS.n5950 0.587457
R10416 AVSS.n3883 AVSS 0.572258
R10417 AVSS.n4094 AVSS 0.572258
R10418 AVSS AVSS.n4104 0.572258
R10419 AVSS AVSS.n3650 0.572258
R10420 AVSS.n3411 AVSS 0.572258
R10421 AVSS.n1614 AVSS 0.572258
R10422 AVSS.n5019 AVSS 0.572258
R10423 AVSS.n5038 AVSS 0.572258
R10424 AVSS.n581 AVSS 0.572258
R10425 AVSS.n1102 AVSS 0.572258
R10426 AVSS.n4487 AVSS 0.572258
R10427 AVSS.n6227 AVSS 0.572258
R10428 AVSS AVSS.n6247 0.572258
R10429 AVSS.n6258 AVSS 0.572258
R10430 AVSS.n5057 AVSS 0.572258
R10431 AVSS.n267 AVSS 0.572258
R10432 AVSS.n6028 AVSS.n6027 0.536293
R10433 AVSS.n6019 AVSS.n6018 0.504971
R10434 AVSS AVSS.n5952 0.492348
R10435 AVSS.n6213 AVSS.n54 0.488676
R10436 AVSS.n5982 AVSS.n5981 0.4655
R10437 AVSS.n6061 AVSS.n6060 0.4655
R10438 AVSS.n2510 AVSS.n2509 0.448417
R10439 AVSS.n2416 AVSS.n1748 0.448417
R10440 AVSS.n1823 AVSS.n1722 0.446929
R10441 AVSS.n2591 AVSS.n2590 0.445861
R10442 AVSS.n6225 AVSS.n6224 0.442488
R10443 AVSS.n6221 AVSS.n6220 0.442488
R10444 AVSS.n6217 AVSS.n6216 0.442488
R10445 AVSS.n6222 AVSS.n6221 0.430929
R10446 AVSS.n6218 AVSS.n6217 0.430929
R10447 AVSS.n6214 AVSS.n6213 0.430929
R10448 AVSS.n6043 AVSS.n6042 0.413543
R10449 AVSS.n6030 AVSS.n6029 0.404848
R10450 AVSS.n6038 AVSS.n6037 0.404848
R10451 AVSS.n6076 AVSS.n6075 0.40216
R10452 AVSS.n6028 AVSS.n6005 0.391804
R10453 AVSS.n6064 AVSS 0.376829
R10454 AVSS.n5974 AVSS.n5968 0.3725
R10455 AVSS.n5988 AVSS.n5972 0.3725
R10456 AVSS.n288 AVSS 0.358259
R10457 AVSS.n5043 AVSS.n5042 0.338559
R10458 AVSS.n6243 AVSS.n6242 0.332538
R10459 AVSS.n5056 AVSS.n5055 0.324904
R10460 AVSS.n6257 AVSS.n6256 0.324904
R10461 AVSS.n6244 AVSS.n6243 0.324904
R10462 AVSS.n6083 AVSS.n263 0.324883
R10463 AVSS.n4113 AVSS.n4097 0.324883
R10464 AVSS.n3887 AVSS.n3886 0.324883
R10465 AVSS.n5027 AVSS.n5026 0.324883
R10466 AVSS.n1619 AVSS.n1610 0.324883
R10467 AVSS.n3416 AVSS.n1622 0.324883
R10468 AVSS.n5044 AVSS.n5043 0.322035
R10469 AVSS.n5055 AVSS.n5054 0.322035
R10470 AVSS.n6256 AVSS.n6255 0.322035
R10471 AVSS.n4113 AVSS.n4112 0.322019
R10472 AVSS.n4086 AVSS.n3887 0.322019
R10473 AVSS.n3875 AVSS.n3676 0.322019
R10474 AVSS.n1610 AVSS.n562 0.322019
R10475 AVSS.n1622 AVSS.n1621 0.322019
R10476 AVSS.n3419 AVSS.n3418 0.322019
R10477 AVSS AVSS.n3882 0.314045
R10478 AVSS AVSS.n4093 0.314045
R10479 AVSS.n4105 AVSS 0.314045
R10480 AVSS.n3673 AVSS 0.314045
R10481 AVSS AVSS.n3398 0.314045
R10482 AVSS AVSS.n1598 0.314045
R10483 AVSS AVSS.n557 0.314045
R10484 AVSS AVSS.n5037 0.314045
R10485 AVSS.n589 AVSS 0.314045
R10486 AVSS.n1110 AVSS 0.314045
R10487 AVSS.n4495 AVSS 0.314045
R10488 AVSS.n6234 AVSS 0.314045
R10489 AVSS.n6248 AVSS 0.314045
R10490 AVSS.n6263 AVSS 0.314045
R10491 AVSS.n5062 AVSS 0.314045
R10492 AVSS AVSS.n266 0.314045
R10493 AVSS.n6002 AVSS.n6001 0.313186
R10494 AVSS.n5971 AVSS.n287 0.313
R10495 AVSS.n6226 AVSS.n6225 0.312199
R10496 AVSS.n5028 AVSS.n5027 0.312199
R10497 AVSS.n3663 AVSS.n3419 0.312199
R10498 AVSS.n3676 AVSS.n3675 0.312199
R10499 AVSS.n6083 AVSS.n6082 0.304186
R10500 AVSS.t84 AVSS.n188 0.290206
R10501 AVSS.t84 AVSS.n190 0.290206
R10502 AVSS.t84 AVSS.n192 0.290206
R10503 AVSS.t84 AVSS.n194 0.290206
R10504 AVSS.t76 AVSS.n2798 0.290206
R10505 AVSS.n1613 AVSS.t78 0.290206
R10506 AVSS.n5018 AVSS.t80 0.290206
R10507 AVSS.n455 AVSS.t104 0.290206
R10508 AVSS.t80 AVSS.n591 0.290206
R10509 AVSS.t78 AVSS.n1112 0.290206
R10510 AVSS.t76 AVSS.n4497 0.290206
R10511 AVSS.t106 AVSS.n6236 0.290206
R10512 AVSS.t92 AVSS.n30 0.290206
R10513 AVSS.t89 AVSS.n6265 0.290206
R10514 AVSS.t99 AVSS.n5064 0.290206
R10515 AVSS.t84 AVSS.n196 0.290206
R10516 AVSS.n280 AVSS.t66 0.283033
R10517 AVSS.n289 AVSS.n288 0.269897
R10518 AVSS.n2195 AVSS.n2194 0.259615
R10519 AVSS.n2415 AVSS.n2302 0.259615
R10520 AVSS.n4712 AVSS.n4711 0.259615
R10521 AVSS.n4680 AVSS.n4679 0.259615
R10522 AVSS.n6063 AVSS.n287 0.220609
R10523 AVSS.n283 AVSS.n282 0.205635
R10524 AVSS.n286 AVSS.n284 0.205635
R10525 AVSS.n281 AVSS.n280 0.204796
R10526 AVSS.n2194 AVSS.n2193 0.195812
R10527 AVSS.n2416 AVSS.n2415 0.195812
R10528 AVSS.n1976 AVSS.n1624 0.195812
R10529 AVSS.n4712 AVSS.n1715 0.195812
R10530 AVSS.n4680 AVSS.n2683 0.195812
R10531 AVSS.n4668 AVSS.n4616 0.195812
R10532 AVSS.n2509 AVSS.n2195 0.19451
R10533 AVSS.n2302 AVSS.n1066 0.19451
R10534 AVSS.n2190 AVSS.n2068 0.19451
R10535 AVSS.n4711 AVSS.n1722 0.19451
R10536 AVSS.n4679 AVSS.n2775 0.19451
R10537 AVSS.n4982 AVSS.n1067 0.19451
R10538 AVSS.n739 AVSS.n738 0.191827
R10539 AVSS.n1198 AVSS.n1197 0.191827
R10540 AVSS.n3122 AVSS.n55 0.191827
R10541 AVSS.n1594 AVSS.n1382 0.191827
R10542 AVSS.n4809 AVSS.n4808 0.191827
R10543 AVSS.n4344 AVSS.n3395 0.191827
R10544 AVSS.n5195 AVSS.n5194 0.191827
R10545 AVSS.n5394 AVSS.n5393 0.191827
R10546 AVSS.n4333 AVSS.n3510 0.191827
R10547 AVSS.n4300 AVSS.n3870 0.191827
R10548 AVSS.n4267 AVSS.n4081 0.191827
R10549 AVSS.n6085 AVSS.n231 0.191827
R10550 AVSS.n833 AVSS.n832 0.190551
R10551 AVSS.n1292 AVSS.n1291 0.190551
R10552 AVSS.n3216 AVSS.n3215 0.190551
R10553 AVSS.n1482 AVSS.n1481 0.190551
R10554 AVSS.n4902 AVSS.n4901 0.190551
R10555 AVSS.n3303 AVSS.n1623 0.190551
R10556 AVSS.n553 AVSS.n552 0.190551
R10557 AVSS.n5101 AVSS.n5100 0.190551
R10558 AVSS.n6303 AVSS.n1 0.190551
R10559 AVSS.n5547 AVSS.n5546 0.190551
R10560 AVSS.n5819 AVSS.n5818 0.190551
R10561 AVSS.n4331 AVSS.n3677 0.190551
R10562 AVSS.n4298 AVSS.n3888 0.190551
R10563 AVSS.n4265 AVSS.n4205 0.190551
R10564 AVSS.n262 AVSS.n147 0.190551
R10565 AVSS.n282 AVSS.n281 0.180177
R10566 AVSS.n284 AVSS.n283 0.180177
R10567 AVSS.n6042 AVSS.n5931 0.175972
R10568 AVSS.n6051 AVSS.n6050 0.175972
R10569 AVSS.n6039 AVSS 0.167167
R10570 AVSS.n2539 AVSS.n1823 0.161214
R10571 AVSS.n2590 AVSS.n1738 0.160444
R10572 AVSS.n2510 AVSS.n1749 0.159726
R10573 AVSS.n2561 AVSS.n1748 0.159726
R10574 AVSS.n6064 AVSS.n286 0.156677
R10575 AVSS.n6004 AVSS.n5935 0.152674
R10576 AVSS.n6026 AVSS.n5934 0.152674
R10577 AVSS.n5977 AVSS 0.151362
R10578 AVSS AVSS.t67 0.146625
R10579 AVSS.n6074 AVSS.t64 0.143939
R10580 AVSS.n6047 AVSS 0.138
R10581 AVSS.n2193 AVSS.n2192 0.133312
R10582 AVSS.n4984 AVSS.n1066 0.133312
R10583 AVSS.n4721 AVSS.n1715 0.13201
R10584 AVSS.n4670 AVSS.n2775 0.13201
R10585 AVSS.n2191 AVSS.n2190 0.130708
R10586 AVSS.n4722 AVSS.n4721 0.130708
R10587 AVSS.n4983 AVSS.n4982 0.130708
R10588 AVSS.n4670 AVSS.n4669 0.130708
R10589 AVSS.n2192 AVSS.n2191 0.129406
R10590 AVSS.n4722 AVSS.n1624 0.129406
R10591 AVSS.n4984 AVSS.n4983 0.129406
R10592 AVSS.n4669 AVSS.n4668 0.129406
R10593 AVSS.n5818 AVSS.n5726 0.129327
R10594 AVSS.n554 AVSS.n553 0.129327
R10595 AVSS.n833 AVSS.n42 0.128051
R10596 AVSS.n6211 AVSS.n147 0.128051
R10597 AVSS.n1482 AVSS.n555 0.128051
R10598 AVSS.n4902 AVSS.n1595 0.128051
R10599 AVSS.n4723 AVSS.n1623 0.128051
R10600 AVSS.n4343 AVSS.n4342 0.128051
R10601 AVSS.n4342 AVSS.n3510 0.128051
R10602 AVSS.n5100 AVSS.n420 0.128051
R10603 AVSS.n5547 AVSS.n24 0.128051
R10604 AVSS.n5819 AVSS.n31 0.128051
R10605 AVSS.n3670 AVSS.n3653 0.128051
R10606 AVSS.n4332 AVSS.n4331 0.128051
R10607 AVSS.n4299 AVSS.n4298 0.128051
R10608 AVSS.n4266 AVSS.n4265 0.128051
R10609 AVSS.n6084 AVSS.n262 0.128051
R10610 AVSS.n6215 AVSS.n6214 0.126783
R10611 AVSS.n6219 AVSS.n6218 0.126783
R10612 AVSS.n6223 AVSS.n6222 0.126783
R10613 AVSS.n5726 AVSS.n42 0.126776
R10614 AVSS.n555 AVSS.n554 0.126776
R10615 AVSS.n1595 AVSS.n1594 0.126776
R10616 AVSS.n4808 AVSS.n4723 0.126776
R10617 AVSS.n4344 AVSS.n4343 0.126776
R10618 AVSS.n552 AVSS.n420 0.126776
R10619 AVSS.n5195 AVSS.n0 0.126776
R10620 AVSS.n5394 AVSS.n24 0.126776
R10621 AVSS.n4300 AVSS.n4299 0.126776
R10622 AVSS.n4267 AVSS.n4266 0.126776
R10623 AVSS.n6085 AVSS.n6084 0.126776
R10624 AVSS.n4333 AVSS.n4332 0.1255
R10625 AVSS AVSS.n6303 0.124224
R10626 AVSS.n6023 AVSS.n6006 0.115315
R10627 AVSS.n6007 AVSS.n6005 0.115315
R10628 AVSS.n6224 AVSS.n6223 0.115224
R10629 AVSS.n6220 AVSS.n6219 0.115224
R10630 AVSS.n6216 AVSS.n6215 0.115224
R10631 AVSS.n6068 AVSS.t70 0.106544
R10632 AVSS.n285 AVSS.t72 0.106544
R10633 AVSS.n279 AVSS.t54 0.106544
R10634 AVSS.n286 AVSS.t56 0.106544
R10635 AVSS.n283 AVSS.t58 0.106544
R10636 AVSS.n281 AVSS.t60 0.106544
R10637 AVSS.n6070 AVSS.t74 0.106544
R10638 AVSS.n6072 AVSS.t62 0.106544
R10639 AVSS.n1292 AVSS.n46 0.0974388
R10640 AVSS.n3216 AVSS.n50 0.0974388
R10641 AVSS.n6212 AVSS.n6211 0.0974388
R10642 AVSS.n738 AVSS.n46 0.0961633
R10643 AVSS.n1197 AVSS.n50 0.0961633
R10644 AVSS.n6212 AVSS.n55 0.0961633
R10645 AVSS.n5953 AVSS 0.0956087
R10646 AVSS.n6040 AVSS.n5932 0.0841694
R10647 AVSS.n6048 AVSS.n5932 0.0841694
R10648 AVSS.n6066 AVSS.n6065 0.0765918
R10649 AVSS.n6065 AVSS.n6064 0.0765918
R10650 AVSS.n5936 AVSS.n5935 0.0755
R10651 AVSS.n6026 AVSS.n5937 0.0755
R10652 AVSS.n6073 AVSS 0.0754063
R10653 AVSS.n3663 AVSS.n3659 0.0706531
R10654 AVSS.n6076 AVSS.n54 0.0557303
R10655 AVSS.n6009 AVSS 0.0548478
R10656 AVSS.n6067 AVSS.n6066 0.0530918
R10657 AVSS.n6073 AVSS.n6072 0.0511182
R10658 AVSS.n6071 AVSS.n6070 0.0511182
R10659 AVSS.n6069 AVSS.n6068 0.0511182
R10660 AVSS.n6062 AVSS.n289 0.0497701
R10661 AVSS.n6072 AVSS.n6071 0.0473173
R10662 AVSS.n6070 AVSS.n6069 0.0473173
R10663 AVSS.n6068 AVSS.n6067 0.0472041
R10664 AVSS.n3658 AVSS.n3657 0.0440606
R10665 AVSS.n461 AVSS.n458 0.043017
R10666 AVSS.n457 AVSS.n452 0.043017
R10667 AVSS.n5042 AVSS.n452 0.043017
R10668 AVSS.n6242 AVSS.n32 0.0428729
R10669 AVSS.n40 AVSS.n32 0.0428729
R10670 AVSS.n6228 AVSS.n39 0.0428729
R10671 AVSS.n6240 AVSS.n34 0.0401825
R10672 AVSS.n6233 AVSS.n6232 0.0401825
R10673 AVSS.n5034 AVSS.n459 0.040057
R10674 AVSS.n5036 AVSS.n453 0.040057
R10675 AVSS.n6075 AVSS.n6074 0.0378951
R10676 AVSS.n6232 AVSS.n6226 0.0342302
R10677 AVSS.n3657 AVSS.n3652 0.033737
R10678 AVSS.n6040 AVSS 0.033
R10679 AVSS.n5984 AVSS.n291 0.0311931
R10680 AVSS.n5976 AVSS.n292 0.0311931
R10681 AVSS.n3667 AVSS.n3659 0.030803
R10682 AVSS.n5028 AVSS.n459 0.0285854
R10683 AVSS.n3675 AVSS.n3641 0.0261503
R10684 AVSS.n5987 AVSS.n5986 0.0260494
R10685 AVSS.n5989 AVSS.n5969 0.0260494
R10686 AVSS.n3672 AVSS.n3670 0.0256047
R10687 AVSS.n5035 AVSS.n458 0.0247347
R10688 AVSS.n41 AVSS.n40 0.0246525
R10689 AVSS.n3668 AVSS.n3658 0.0246141
R10690 AVSS.n3662 AVSS.n3661 0.0246141
R10691 AVSS.n3665 AVSS.n3655 0.0246141
R10692 AVSS.n3668 AVSS.n3667 0.0246141
R10693 AVSS.n3661 AVSS.n3656 0.0246141
R10694 AVSS.n3662 AVSS.n3655 0.0246141
R10695 AVSS.n6074 AVSS.n6073 0.024
R10696 AVSS.n41 AVSS.n34 0.023119
R10697 AVSS.n5035 AVSS.n5034 0.0230475
R10698 AVSS.n5048 AVSS.n5044 0.0209918
R10699 AVSS.n5049 AVSS.n5048 0.0209918
R10700 AVSS.n5061 AVSS.n5049 0.0209918
R10701 AVSS.n5061 AVSS.n5060 0.0209918
R10702 AVSS.n5060 AVSS.n5056 0.0209918
R10703 AVSS.n5054 AVSS.n5050 0.0209918
R10704 AVSS.n5050 AVSS.n23 0.0209918
R10705 AVSS.n6262 AVSS.n23 0.0209918
R10706 AVSS.n6262 AVSS.n6261 0.0209918
R10707 AVSS.n6261 AVSS.n6257 0.0209918
R10708 AVSS.n6255 AVSS.n25 0.0209918
R10709 AVSS.n6250 AVSS.n25 0.0209918
R10710 AVSS.n6250 AVSS.n6249 0.0209918
R10711 AVSS.n6249 AVSS.n28 0.0209918
R10712 AVSS.n6244 AVSS.n28 0.0209918
R10713 AVSS.n4112 AVSS.n4098 0.0209583
R10714 AVSS.n4107 AVSS.n4098 0.0209583
R10715 AVSS.n4107 AVSS.n4106 0.0209583
R10716 AVSS.n4106 AVSS.n4100 0.0209583
R10717 AVSS.n4100 AVSS.n263 0.0209583
R10718 AVSS.n4086 AVSS.n4085 0.0209583
R10719 AVSS.n4091 AVSS.n4085 0.0209583
R10720 AVSS.n4092 AVSS.n4091 0.0209583
R10721 AVSS.n4092 AVSS.n4082 0.0209583
R10722 AVSS.n4097 AVSS.n4082 0.0209583
R10723 AVSS.n3875 AVSS.n3874 0.0209583
R10724 AVSS.n3880 AVSS.n3874 0.0209583
R10725 AVSS.n3881 AVSS.n3880 0.0209583
R10726 AVSS.n3881 AVSS.n3871 0.0209583
R10727 AVSS.n3886 AVSS.n3871 0.0209583
R10728 AVSS.n3659 AVSS.n3653 0.0209082
R10729 AVSS.n6082 AVSS.n264 0.019586
R10730 AVSS.n3671 AVSS.n3647 0.0190286
R10731 AVSS.n3651 AVSS.n3647 0.0190286
R10732 AVSS.n3645 AVSS.n3641 0.0190286
R10733 AVSS.n3652 AVSS.n3651 0.0190286
R10734 AVSS.n3646 AVSS.n3645 0.0190286
R10735 AVSS.n3672 AVSS.n3671 0.0190286
R10736 AVSS.n5035 AVSS.n457 0.0187823
R10737 AVSS.n41 AVSS.n39 0.0187203
R10738 AVSS.n6233 AVSS.n41 0.0175635
R10739 AVSS.n5036 AVSS.n5035 0.0175095
R10740 AVSS.n6223 AVSS.n45 0.0161593
R10741 AVSS.n6219 AVSS.n49 0.0161593
R10742 AVSS.n6215 AVSS.n53 0.0161593
R10743 AVSS.n6076 AVSS.n275 0.0155538
R10744 AVSS.n588 AVSS.n585 0.014716
R10745 AVSS.n578 AVSS.n44 0.014716
R10746 AVSS.n579 AVSS.n576 0.014716
R10747 AVSS.n582 AVSS.n574 0.014716
R10748 AVSS.n585 AVSS.n575 0.014716
R10749 AVSS.n578 AVSS.n575 0.014716
R10750 AVSS.n579 AVSS.n45 0.014716
R10751 AVSS.n582 AVSS.n576 0.014716
R10752 AVSS.n1109 AVSS.n1106 0.014716
R10753 AVSS.n1099 AVSS.n48 0.014716
R10754 AVSS.n1100 AVSS.n1097 0.014716
R10755 AVSS.n1103 AVSS.n1095 0.014716
R10756 AVSS.n1106 AVSS.n1096 0.014716
R10757 AVSS.n1099 AVSS.n1096 0.014716
R10758 AVSS.n1100 AVSS.n49 0.014716
R10759 AVSS.n1103 AVSS.n1097 0.014716
R10760 AVSS.n4494 AVSS.n4491 0.014716
R10761 AVSS.n4484 AVSS.n52 0.014716
R10762 AVSS.n4485 AVSS.n4482 0.014716
R10763 AVSS.n4488 AVSS.n4480 0.014716
R10764 AVSS.n4491 AVSS.n4481 0.014716
R10765 AVSS.n4484 AVSS.n4481 0.014716
R10766 AVSS.n4485 AVSS.n53 0.014716
R10767 AVSS.n4488 AVSS.n4482 0.014716
R10768 AVSS.n6078 AVSS.n276 0.0144215
R10769 AVSS.n6077 AVSS.n278 0.0144215
R10770 AVSS.n274 AVSS.n264 0.0144215
R10771 AVSS.n278 AVSS.n276 0.0144215
R10772 AVSS.n275 AVSS.n274 0.0144215
R10773 AVSS.n6079 AVSS.n6078 0.0144215
R10774 AVSS.n287 AVSS 0.014087
R10775 AVSS.n6077 AVSS.n6076 0.012328
R10776 AVSS.n6223 AVSS.n44 0.0123132
R10777 AVSS.n6219 AVSS.n48 0.0123132
R10778 AVSS.n6215 AVSS.n52 0.0123132
R10779 AVSS.n5026 AVSS.n558 0.0112179
R10780 AVSS.n566 AVSS.n565 0.0112179
R10781 AVSS.n568 AVSS.n563 0.0112179
R10782 AVSS.n5024 AVSS.n567 0.0112179
R10783 AVSS.n5023 AVSS.n562 0.0112179
R10784 AVSS.n564 AVSS.n558 0.0112179
R10785 AVSS.n565 AVSS.n564 0.0112179
R10786 AVSS.n568 AVSS.n566 0.0112179
R10787 AVSS.n567 AVSS.n563 0.0112179
R10788 AVSS.n5024 AVSS.n5023 0.0112179
R10789 AVSS.n1619 AVSS.n1618 0.0112179
R10790 AVSS.n1607 AVSS.n1606 0.0112179
R10791 AVSS.n1611 AVSS.n1604 0.0112179
R10792 AVSS.n1609 AVSS.n1608 0.0112179
R10793 AVSS.n1621 AVSS.n1596 0.0112179
R10794 AVSS.n1618 AVSS.n1605 0.0112179
R10795 AVSS.n1606 AVSS.n1605 0.0112179
R10796 AVSS.n1611 AVSS.n1607 0.0112179
R10797 AVSS.n1608 AVSS.n1604 0.0112179
R10798 AVSS.n1609 AVSS.n1596 0.0112179
R10799 AVSS.n3416 AVSS.n3415 0.0112179
R10800 AVSS.n3407 AVSS.n3406 0.0112179
R10801 AVSS.n3410 AVSS.n3404 0.0112179
R10802 AVSS.n3409 AVSS.n3408 0.0112179
R10803 AVSS.n3418 AVSS.n3396 0.0112179
R10804 AVSS.n3415 AVSS.n3405 0.0112179
R10805 AVSS.n3406 AVSS.n3405 0.0112179
R10806 AVSS.n3410 AVSS.n3407 0.0112179
R10807 AVSS.n3408 AVSS.n3404 0.0112179
R10808 AVSS.n3409 AVSS.n3396 0.0112179
R10809 AVSS.n3675 AVSS.n3674 0.0109769
R10810 AVSS.n6082 AVSS.n6081 0.0082957
R10811 AVSS AVSS.n0 0.00432653
R10812 AVSS.n3657 AVSS.n3656 0.00428788
R10813 AVSS.n3657 AVSS.n3646 0.00339017
R10814 AVSS.n6067 AVSS.t69 0.00329016
R10815 AVSS.n280 AVSS.t65 0.00317698
R10816 AVSS.n282 AVSS.t59 0.00317698
R10817 AVSS.n284 AVSS.t57 0.00317698
R10818 AVSS.n6073 AVSS.t63 0.00317698
R10819 AVSS.n6071 AVSS.t61 0.00317698
R10820 AVSS.n6069 AVSS.t73 0.00317698
R10821 AVSS.n6066 AVSS.t53 0.00317698
R10822 AVSS.n6065 AVSS.t71 0.00317698
R10823 AVSS.n6064 AVSS.t55 0.00317698
R10824 AVSS.n2683 AVSS.n2591 0.00180208
R10825 TRIM0.t2 TRIM0 190.643
R10826 TRIM0.t1 TRIM0.n1 190.585
R10827 TRIM0.n1 TRIM0.t0 190.585
R10828 TRIM0 TRIM0.t3 190.553
R10829 TRIM0.t0 TRIM0.n0 119.778
R10830 TRIM0.n0 TRIM0.t2 119.778
R10831 TRIM0.t3 TRIM0.n2 119.778
R10832 TRIM0.n2 TRIM0.t1 119.778
R10833 TRIM0.n2 TRIM0.n0 19.6878
R10834 TRIM0.n1 TRIM0 13.1688
R10835 bjt_0.B.n195 bjt_0.B.n194 83.5719
R10836 bjt_0.B.n37 bjt_0.B.n35 83.5719
R10837 bjt_0.B.n100 bjt_0.B.n98 83.5719
R10838 bjt_0.B.n185 bjt_0.B.n184 83.5719
R10839 bjt_0.B.n183 bjt_0.B.n182 83.5719
R10840 bjt_0.B.n181 bjt_0.B.n180 83.5719
R10841 bjt_0.B.n61 bjt_0.B.n60 83.5719
R10842 bjt_0.B.n59 bjt_0.B.n58 83.5719
R10843 bjt_0.B.n57 bjt_0.B.n56 83.5719
R10844 bjt_0.B.n165 bjt_0.B.n66 83.5719
R10845 bjt_0.B.n158 bjt_0.B.n67 83.5719
R10846 bjt_0.B.n160 bjt_0.B.n159 83.5719
R10847 bjt_0.B.n152 bjt_0.B.n71 83.5719
R10848 bjt_0.B.n145 bjt_0.B.n72 83.5719
R10849 bjt_0.B.n147 bjt_0.B.n146 83.5719
R10850 bjt_0.B.n136 bjt_0.B.n135 83.5719
R10851 bjt_0.B.n134 bjt_0.B.n133 83.5719
R10852 bjt_0.B.n132 bjt_0.B.n131 83.5719
R10853 bjt_0.B.n117 bjt_0.B.n90 83.5719
R10854 bjt_0.B.n124 bjt_0.B.n123 83.5719
R10855 bjt_0.B.n126 bjt_0.B.n125 83.5719
R10856 bjt_0.B.n107 bjt_0.B.n106 83.5719
R10857 bjt_0.B.n96 bjt_0.B.n93 83.5719
R10858 bjt_0.B.n112 bjt_0.B.n92 83.5719
R10859 bjt_0.B.n194 bjt_0.B.n193 73.3165
R10860 bjt_0.B.n186 bjt_0.B.n185 73.3165
R10861 bjt_0.B.n62 bjt_0.B.n61 73.3165
R10862 bjt_0.B.n167 bjt_0.B.n66 73.3165
R10863 bjt_0.B.n154 bjt_0.B.n71 73.3165
R10864 bjt_0.B.n137 bjt_0.B.n136 73.3165
R10865 bjt_0.B.n118 bjt_0.B.n90 73.3165
R10866 bjt_0.B.n106 bjt_0.B.n105 73.3165
R10867 bjt_0.B.n102 bjt_0.B.n98 73.19
R10868 bjt_0.B.n181 bjt_0.B.n43 73.19
R10869 bjt_0.B.n57 bjt_0.B.n49 73.19
R10870 bjt_0.B.n159 bjt_0.B.n157 73.19
R10871 bjt_0.B.n146 bjt_0.B.n144 73.19
R10872 bjt_0.B.n132 bjt_0.B.n80 73.19
R10873 bjt_0.B.n125 bjt_0.B.n87 73.19
R10874 bjt_0.B.n114 bjt_0.B.n92 73.19
R10875 bjt_0.B.n3 bjt_0.B.t16 43.9266
R10876 bjt_0.B.n16 bjt_0.B.t3 43.5116
R10877 bjt_0.B.n10 bjt_0.B.t37 43.5116
R10878 bjt_0.B.n2 bjt_0.B.t12 43.3041
R10879 bjt_0.B.n26 bjt_0.B.t1 43.3041
R10880 bjt_0.B.n3 bjt_0.B.t4 43.2216
R10881 bjt_0.B.n5 bjt_0.B.t18 43.2216
R10882 bjt_0.B.n17 bjt_0.B.t41 43.2216
R10883 bjt_0.B.n19 bjt_0.B.t36 43.2216
R10884 bjt_0.B.n22 bjt_0.B.t39 43.2216
R10885 bjt_0.B.n11 bjt_0.B.t15 43.2216
R10886 bjt_0.B.n13 bjt_0.B.t34 43.2216
R10887 bjt_0.B.n15 bjt_0.B.t0 43.1241
R10888 bjt_0.B.n9 bjt_0.B.t11 43.1241
R10889 bjt_0.B.n24 bjt_0.B.t43 43.0966
R10890 bjt_0.B.n30 bjt_0.B.t33 43.0966
R10891 bjt_0.B.n4 bjt_0.B.t40 43.0416
R10892 bjt_0.B.n6 bjt_0.B.t17 43.0416
R10893 bjt_0.B.n16 bjt_0.B.t8 43.0416
R10894 bjt_0.B.n18 bjt_0.B.t7 43.0416
R10895 bjt_0.B.n19 bjt_0.B.t2 43.0416
R10896 bjt_0.B.n10 bjt_0.B.t19 43.0416
R10897 bjt_0.B.n12 bjt_0.B.t6 43.0416
R10898 bjt_0.B.n14 bjt_0.B.t5 43.0416
R10899 bjt_0.B.n2 bjt_0.B.t10 43.0141
R10900 bjt_0.B.n26 bjt_0.B.t14 43.0141
R10901 bjt_0.B.n20 bjt_0.B.t38 42.9166
R10902 bjt_0.B.n20 bjt_0.B.t35 42.9166
R10903 bjt_0.B.n23 bjt_0.B.t42 42.9166
R10904 bjt_0.B.n29 bjt_0.B.t32 42.9166
R10905 bjt_0.B.n15 bjt_0.B.t13 42.8341
R10906 bjt_0.B.n8 bjt_0.B.t9 42.3691
R10907 bjt_0.B.n194 bjt_0.B.n37 26.074
R10908 bjt_0.B.n185 bjt_0.B.n183 26.074
R10909 bjt_0.B.n61 bjt_0.B.n59 26.074
R10910 bjt_0.B.n158 bjt_0.B.n66 26.074
R10911 bjt_0.B.n145 bjt_0.B.n71 26.074
R10912 bjt_0.B.n136 bjt_0.B.n134 26.074
R10913 bjt_0.B.n124 bjt_0.B.n90 26.074
R10914 bjt_0.B.n106 bjt_0.B.n96 26.074
R10915 bjt_0.B.n98 bjt_0.B.t26 25.7843
R10916 bjt_0.B.t21 bjt_0.B.n181 25.7843
R10917 bjt_0.B.t22 bjt_0.B.n57 25.7843
R10918 bjt_0.B.n159 bjt_0.B.t20 25.7843
R10919 bjt_0.B.n146 bjt_0.B.t24 25.7843
R10920 bjt_0.B.t23 bjt_0.B.n132 25.7843
R10921 bjt_0.B.n125 bjt_0.B.t27 25.7843
R10922 bjt_0.B.t25 bjt_0.B.n92 25.7843
R10923 bjt_0.B.n199 bjt_0.B.n32 22.2712
R10924 bjt_0.B.n1 bjt_0.B.n0 18.0391
R10925 bjt_0.B.n201 bjt_0.B.n200 18.0391
R10926 bjt_0.B.n82 bjt_0.B.n78 9.3005
R10927 bjt_0.B.n82 bjt_0.B.n77 9.3005
R10928 bjt_0.B.n82 bjt_0.B.n79 9.3005
R10929 bjt_0.B.n141 bjt_0.B.n82 9.3005
R10930 bjt_0.B.n84 bjt_0.B.n78 9.3005
R10931 bjt_0.B.n84 bjt_0.B.n77 9.3005
R10932 bjt_0.B.n84 bjt_0.B.n79 9.3005
R10933 bjt_0.B.n141 bjt_0.B.n84 9.3005
R10934 bjt_0.B.n81 bjt_0.B.n78 9.3005
R10935 bjt_0.B.n81 bjt_0.B.n77 9.3005
R10936 bjt_0.B.n81 bjt_0.B.n79 9.3005
R10937 bjt_0.B.n141 bjt_0.B.n81 9.3005
R10938 bjt_0.B.n86 bjt_0.B.n78 9.3005
R10939 bjt_0.B.n86 bjt_0.B.n77 9.3005
R10940 bjt_0.B.n86 bjt_0.B.n79 9.3005
R10941 bjt_0.B.n141 bjt_0.B.n86 9.3005
R10942 bjt_0.B.n142 bjt_0.B.n78 9.3005
R10943 bjt_0.B.n142 bjt_0.B.n77 9.3005
R10944 bjt_0.B.n142 bjt_0.B.n79 9.3005
R10945 bjt_0.B.n142 bjt_0.B.n76 9.3005
R10946 bjt_0.B.n142 bjt_0.B.n141 9.3005
R10947 bjt_0.B.n140 bjt_0.B.n78 9.3005
R10948 bjt_0.B.n140 bjt_0.B.n77 9.3005
R10949 bjt_0.B.n140 bjt_0.B.n79 9.3005
R10950 bjt_0.B.n140 bjt_0.B.n76 9.3005
R10951 bjt_0.B.n141 bjt_0.B.n140 9.3005
R10952 bjt_0.B.n52 bjt_0.B.n47 9.3005
R10953 bjt_0.B.n52 bjt_0.B.n45 9.3005
R10954 bjt_0.B.n52 bjt_0.B.n48 9.3005
R10955 bjt_0.B.n171 bjt_0.B.n52 9.3005
R10956 bjt_0.B.n63 bjt_0.B.n55 9.3005
R10957 bjt_0.B.n55 bjt_0.B.n47 9.3005
R10958 bjt_0.B.n55 bjt_0.B.n48 9.3005
R10959 bjt_0.B.n171 bjt_0.B.n55 9.3005
R10960 bjt_0.B.n51 bjt_0.B.n47 9.3005
R10961 bjt_0.B.n51 bjt_0.B.n48 9.3005
R10962 bjt_0.B.n51 bjt_0.B.n44 9.3005
R10963 bjt_0.B.n171 bjt_0.B.n51 9.3005
R10964 bjt_0.B.n170 bjt_0.B.n47 9.3005
R10965 bjt_0.B.n170 bjt_0.B.n45 9.3005
R10966 bjt_0.B.n170 bjt_0.B.n48 9.3005
R10967 bjt_0.B.n170 bjt_0.B.n44 9.3005
R10968 bjt_0.B.n171 bjt_0.B.n170 9.3005
R10969 bjt_0.B.n63 bjt_0.B.n50 9.3005
R10970 bjt_0.B.n50 bjt_0.B.n47 9.3005
R10971 bjt_0.B.n50 bjt_0.B.n45 9.3005
R10972 bjt_0.B.n50 bjt_0.B.n48 9.3005
R10973 bjt_0.B.n50 bjt_0.B.n44 9.3005
R10974 bjt_0.B.n171 bjt_0.B.n50 9.3005
R10975 bjt_0.B.n172 bjt_0.B.n47 9.3005
R10976 bjt_0.B.n172 bjt_0.B.n45 9.3005
R10977 bjt_0.B.n172 bjt_0.B.n48 9.3005
R10978 bjt_0.B.n172 bjt_0.B.n44 9.3005
R10979 bjt_0.B.n172 bjt_0.B.n171 9.3005
R10980 bjt_0.B.n175 bjt_0.B.n41 9.3005
R10981 bjt_0.B.n175 bjt_0.B.n39 9.3005
R10982 bjt_0.B.n175 bjt_0.B.n42 9.3005
R10983 bjt_0.B.n190 bjt_0.B.n175 9.3005
R10984 bjt_0.B.n177 bjt_0.B.n41 9.3005
R10985 bjt_0.B.n177 bjt_0.B.n39 9.3005
R10986 bjt_0.B.n177 bjt_0.B.n42 9.3005
R10987 bjt_0.B.n190 bjt_0.B.n177 9.3005
R10988 bjt_0.B.n174 bjt_0.B.n41 9.3005
R10989 bjt_0.B.n174 bjt_0.B.n39 9.3005
R10990 bjt_0.B.n174 bjt_0.B.n42 9.3005
R10991 bjt_0.B.n190 bjt_0.B.n174 9.3005
R10992 bjt_0.B.n189 bjt_0.B.n41 9.3005
R10993 bjt_0.B.n189 bjt_0.B.n39 9.3005
R10994 bjt_0.B.n189 bjt_0.B.n42 9.3005
R10995 bjt_0.B.n190 bjt_0.B.n189 9.3005
R10996 bjt_0.B.n173 bjt_0.B.n41 9.3005
R10997 bjt_0.B.n173 bjt_0.B.n39 9.3005
R10998 bjt_0.B.n173 bjt_0.B.n42 9.3005
R10999 bjt_0.B.n173 bjt_0.B.n38 9.3005
R11000 bjt_0.B.n190 bjt_0.B.n173 9.3005
R11001 bjt_0.B.n191 bjt_0.B.n41 9.3005
R11002 bjt_0.B.n191 bjt_0.B.n39 9.3005
R11003 bjt_0.B.n191 bjt_0.B.n42 9.3005
R11004 bjt_0.B.n191 bjt_0.B.n38 9.3005
R11005 bjt_0.B.n191 bjt_0.B.n190 9.3005
R11006 bjt_0.B.n21 bjt_0.B.n20 6.333
R11007 bjt_0.B.n24 bjt_0.B.n23 6.1255
R11008 bjt_0.B.n27 bjt_0.B.n25 6.1255
R11009 bjt_0.B.n30 bjt_0.B.n29 6.1255
R11010 bjt_0.B.n32 bjt_0.B.n7 5.5255
R11011 bjt_0.B.n201 bjt_0.B.n199 5.28993
R11012 bjt_0.B.n199 bjt_0.B.n198 5.08174
R11013 bjt_0.B.n83 bjt_0.B.n76 4.64588
R11014 bjt_0.B.n138 bjt_0.B.n130 4.64588
R11015 bjt_0.B.n85 bjt_0.B.n76 4.64588
R11016 bjt_0.B.n138 bjt_0.B.n75 4.64588
R11017 bjt_0.B.n139 bjt_0.B.n138 4.64588
R11018 bjt_0.B.n53 bjt_0.B.n44 4.64588
R11019 bjt_0.B.n54 bjt_0.B.n45 4.64588
R11020 bjt_0.B.n64 bjt_0.B.n63 4.64588
R11021 bjt_0.B.n63 bjt_0.B.n46 4.64588
R11022 bjt_0.B.n176 bjt_0.B.n38 4.64588
R11023 bjt_0.B.n187 bjt_0.B.n179 4.64588
R11024 bjt_0.B.n178 bjt_0.B.n38 4.64588
R11025 bjt_0.B.n188 bjt_0.B.n187 4.64588
R11026 bjt_0.B.n187 bjt_0.B.n40 4.64588
R11027 bjt_0.B.n0 bjt_0.B.t31 4.3505
R11028 bjt_0.B.n0 bjt_0.B.t30 4.3505
R11029 bjt_0.B.n200 bjt_0.B.t29 4.3505
R11030 bjt_0.B.n200 bjt_0.B.t28 4.3505
R11031 bjt_0.B.n144 bjt_0.B.n143 2.36574
R11032 bjt_0.B.n129 bjt_0.B.n87 2.36574
R11033 bjt_0.B.n103 bjt_0.B.n102 2.36206
R11034 bjt_0.B.n157 bjt_0.B.n156 2.36206
R11035 bjt_0.B.n115 bjt_0.B.n114 2.36206
R11036 bjt_0.B.n193 bjt_0.B.n192 2.19824
R11037 bjt_0.B.n168 bjt_0.B.n167 2.19742
R11038 bjt_0.B.n155 bjt_0.B.n154 2.19742
R11039 bjt_0.B.n118 bjt_0.B.n116 2.19742
R11040 bjt_0.B.n105 bjt_0.B.n104 2.19742
R11041 bjt_0.B.n95 bjt_0.B.n94 1.5505
R11042 bjt_0.B.n109 bjt_0.B.n108 1.5505
R11043 bjt_0.B.n111 bjt_0.B.n110 1.5505
R11044 bjt_0.B.n113 bjt_0.B.n91 1.5505
R11045 bjt_0.B.n120 bjt_0.B.n119 1.5505
R11046 bjt_0.B.n122 bjt_0.B.n121 1.5505
R11047 bjt_0.B.n89 bjt_0.B.n88 1.5505
R11048 bjt_0.B.n128 bjt_0.B.n127 1.5505
R11049 bjt_0.B.n153 bjt_0.B.n70 1.5505
R11050 bjt_0.B.n151 bjt_0.B.n150 1.5505
R11051 bjt_0.B.n149 bjt_0.B.n148 1.5505
R11052 bjt_0.B.n74 bjt_0.B.n73 1.5505
R11053 bjt_0.B.n166 bjt_0.B.n65 1.5505
R11054 bjt_0.B.n164 bjt_0.B.n163 1.5505
R11055 bjt_0.B.n162 bjt_0.B.n161 1.5505
R11056 bjt_0.B.n69 bjt_0.B.n68 1.5505
R11057 bjt_0.B.n36 bjt_0.B.n34 1.5505
R11058 bjt_0.B.n197 bjt_0.B.n196 1.5505
R11059 bjt_0.B.n99 bjt_0.B.n33 1.5505
R11060 bjt_0.B.n101 bjt_0.B.n97 1.5505
R11061 bjt_0.B bjt_0.B.n1 1.39954
R11062 bjt_0.B.n101 bjt_0.B.n100 1.25468
R11063 bjt_0.B.n180 bjt_0.B.n38 1.25468
R11064 bjt_0.B.n56 bjt_0.B.n44 1.25468
R11065 bjt_0.B.n160 bjt_0.B.n69 1.25468
R11066 bjt_0.B.n147 bjt_0.B.n74 1.25468
R11067 bjt_0.B.n131 bjt_0.B.n76 1.25468
R11068 bjt_0.B.n127 bjt_0.B.n126 1.25468
R11069 bjt_0.B.n113 bjt_0.B.n112 1.25468
R11070 bjt_0.B.n193 bjt_0.B.n36 1.19225
R11071 bjt_0.B.n186 bjt_0.B.n41 1.19225
R11072 bjt_0.B.n62 bjt_0.B.n47 1.19225
R11073 bjt_0.B.n167 bjt_0.B.n166 1.19225
R11074 bjt_0.B.n154 bjt_0.B.n153 1.19225
R11075 bjt_0.B.n137 bjt_0.B.n78 1.19225
R11076 bjt_0.B.n119 bjt_0.B.n118 1.19225
R11077 bjt_0.B.n105 bjt_0.B.n95 1.19225
R11078 bjt_0.B.n99 bjt_0.B.n35 1.07024
R11079 bjt_0.B.n182 bjt_0.B.n42 1.07024
R11080 bjt_0.B.n58 bjt_0.B.n48 1.07024
R11081 bjt_0.B.n161 bjt_0.B.n67 1.07024
R11082 bjt_0.B.n148 bjt_0.B.n72 1.07024
R11083 bjt_0.B.n133 bjt_0.B.n79 1.07024
R11084 bjt_0.B.n123 bjt_0.B.n89 1.07024
R11085 bjt_0.B.n111 bjt_0.B.n93 1.07024
R11086 bjt_0.B.n102 bjt_0.B.n101 1.0237
R11087 bjt_0.B.n43 bjt_0.B.n38 1.0237
R11088 bjt_0.B.n49 bjt_0.B.n44 1.0237
R11089 bjt_0.B.n157 bjt_0.B.n69 1.0237
R11090 bjt_0.B.n144 bjt_0.B.n74 1.0237
R11091 bjt_0.B.n80 bjt_0.B.n76 1.0237
R11092 bjt_0.B.n127 bjt_0.B.n87 1.0237
R11093 bjt_0.B.n114 bjt_0.B.n113 1.0237
R11094 bjt_0.B bjt_0.B.n201 0.990885
R11095 bjt_0.B.n195 bjt_0.B.n36 0.959578
R11096 bjt_0.B.n184 bjt_0.B.n41 0.959578
R11097 bjt_0.B.n60 bjt_0.B.n47 0.959578
R11098 bjt_0.B.n166 bjt_0.B.n165 0.959578
R11099 bjt_0.B.n153 bjt_0.B.n152 0.959578
R11100 bjt_0.B.n135 bjt_0.B.n78 0.959578
R11101 bjt_0.B.n119 bjt_0.B.n117 0.959578
R11102 bjt_0.B.n107 bjt_0.B.n95 0.959578
R11103 bjt_0.B.n1 bjt_0.B 0.928385
R11104 bjt_0.B.n190 bjt_0.B.n43 0.812055
R11105 bjt_0.B.n171 bjt_0.B.n49 0.812055
R11106 bjt_0.B.n141 bjt_0.B.n80 0.812055
R11107 bjt_0.B.n196 bjt_0.B.n35 0.77514
R11108 bjt_0.B.n182 bjt_0.B.n39 0.77514
R11109 bjt_0.B.n58 bjt_0.B.n45 0.77514
R11110 bjt_0.B.n164 bjt_0.B.n67 0.77514
R11111 bjt_0.B.n151 bjt_0.B.n72 0.77514
R11112 bjt_0.B.n133 bjt_0.B.n77 0.77514
R11113 bjt_0.B.n123 bjt_0.B.n122 0.77514
R11114 bjt_0.B.n108 bjt_0.B.n93 0.77514
R11115 bjt_0.B.n116 bjt_0.B.n115 0.759783
R11116 bjt_0.B.n156 bjt_0.B.n155 0.759783
R11117 bjt_0.B.n173 bjt_0.B.n172 0.759783
R11118 bjt_0.B.n140 bjt_0.B.n129 0.749947
R11119 bjt_0.B.n169 bjt_0.B.n168 0.749947
R11120 bjt_0.B.n192 bjt_0.B.n191 0.749947
R11121 bjt_0.B.n143 bjt_0.B.n142 0.747079
R11122 bjt_0.B.n7 bjt_0.B.n6 0.7055
R11123 bjt_0.B.n19 bjt_0.B.n18 0.7055
R11124 bjt_0.B.n187 bjt_0.B.n186 0.647417
R11125 bjt_0.B.n63 bjt_0.B.n62 0.647417
R11126 bjt_0.B.n138 bjt_0.B.n137 0.647417
R11127 bjt_0.B.n100 bjt_0.B.n99 0.590702
R11128 bjt_0.B.n180 bjt_0.B.n42 0.590702
R11129 bjt_0.B.n56 bjt_0.B.n48 0.590702
R11130 bjt_0.B.n161 bjt_0.B.n160 0.590702
R11131 bjt_0.B.n148 bjt_0.B.n147 0.590702
R11132 bjt_0.B.n131 bjt_0.B.n79 0.590702
R11133 bjt_0.B.n126 bjt_0.B.n89 0.590702
R11134 bjt_0.B.n112 bjt_0.B.n111 0.590702
R11135 bjt_0.B bjt_0.B.n195 0.572258
R11136 bjt_0.B.n184 bjt_0.B 0.572258
R11137 bjt_0.B.n60 bjt_0.B 0.572258
R11138 bjt_0.B.n165 bjt_0.B 0.572258
R11139 bjt_0.B.n152 bjt_0.B 0.572258
R11140 bjt_0.B.n135 bjt_0.B 0.572258
R11141 bjt_0.B.n117 bjt_0.B 0.572258
R11142 bjt_0.B bjt_0.B.n107 0.572258
R11143 bjt_0.B.n25 bjt_0.B.n24 0.4155
R11144 bjt_0.B.n31 bjt_0.B.n30 0.4155
R11145 bjt_0.B bjt_0.B.n103 0.382495
R11146 bjt_0.B.n104 bjt_0.B 0.377788
R11147 bjt_0.B.n196 bjt_0.B 0.314045
R11148 bjt_0.B bjt_0.B.n39 0.314045
R11149 bjt_0.B bjt_0.B.n45 0.314045
R11150 bjt_0.B bjt_0.B.n164 0.314045
R11151 bjt_0.B bjt_0.B.n151 0.314045
R11152 bjt_0.B bjt_0.B.n77 0.314045
R11153 bjt_0.B.n122 bjt_0.B 0.314045
R11154 bjt_0.B.n108 bjt_0.B 0.314045
R11155 bjt_0.B.n4 bjt_0.B.n3 0.2905
R11156 bjt_0.B.n5 bjt_0.B.n4 0.2905
R11157 bjt_0.B.n6 bjt_0.B.n5 0.2905
R11158 bjt_0.B.n17 bjt_0.B.n16 0.2905
R11159 bjt_0.B.n18 bjt_0.B.n17 0.2905
R11160 bjt_0.B.n23 bjt_0.B.n22 0.2905
R11161 bjt_0.B.n11 bjt_0.B.n10 0.2905
R11162 bjt_0.B.n12 bjt_0.B.n11 0.2905
R11163 bjt_0.B.n13 bjt_0.B.n12 0.2905
R11164 bjt_0.B.n14 bjt_0.B.n13 0.2905
R11165 bjt_0.B.t26 bjt_0.B.n37 0.290206
R11166 bjt_0.B.n183 bjt_0.B.t21 0.290206
R11167 bjt_0.B.n59 bjt_0.B.t22 0.290206
R11168 bjt_0.B.t20 bjt_0.B.n158 0.290206
R11169 bjt_0.B.t24 bjt_0.B.n145 0.290206
R11170 bjt_0.B.n134 bjt_0.B.t23 0.290206
R11171 bjt_0.B.t27 bjt_0.B.n124 0.290206
R11172 bjt_0.B.n96 bjt_0.B.t25 0.290206
R11173 bjt_0.B.n28 bjt_0.B 0.2805
R11174 bjt_0.B.n9 bjt_0.B.n8 0.2655
R11175 bjt_0.B.n32 bjt_0.B.n31 0.2655
R11176 bjt_0.B bjt_0.B.n14 0.218
R11177 bjt_0.B.n28 bjt_0.B.n27 0.208
R11178 bjt_0.B.n29 bjt_0.B.n28 0.208
R11179 bjt_0.B.n7 bjt_0.B.n2 0.083
R11180 bjt_0.B.n21 bjt_0.B.n19 0.083
R11181 bjt_0.B.n22 bjt_0.B.n21 0.083
R11182 bjt_0.B.n25 bjt_0.B.n15 0.083
R11183 bjt_0.B.n31 bjt_0.B.n9 0.083
R11184 bjt_0.B.n27 bjt_0.B.n26 0.083
R11185 bjt_0.B.n32 bjt_0.B.n8 0.0779254
R11186 bjt_0.B.n115 bjt_0.B.n91 0.0209918
R11187 bjt_0.B.n110 bjt_0.B.n91 0.0209918
R11188 bjt_0.B.n110 bjt_0.B.n109 0.0209918
R11189 bjt_0.B.n109 bjt_0.B.n94 0.0209918
R11190 bjt_0.B.n104 bjt_0.B.n94 0.0209918
R11191 bjt_0.B.n128 bjt_0.B.n88 0.0209918
R11192 bjt_0.B.n121 bjt_0.B.n88 0.0209918
R11193 bjt_0.B.n121 bjt_0.B.n120 0.0209918
R11194 bjt_0.B.n120 bjt_0.B.n116 0.0209918
R11195 bjt_0.B.n149 bjt_0.B.n73 0.0209918
R11196 bjt_0.B.n150 bjt_0.B.n149 0.0209918
R11197 bjt_0.B.n150 bjt_0.B.n70 0.0209918
R11198 bjt_0.B.n155 bjt_0.B.n70 0.0209918
R11199 bjt_0.B.n156 bjt_0.B.n68 0.0209918
R11200 bjt_0.B.n162 bjt_0.B.n68 0.0209918
R11201 bjt_0.B.n163 bjt_0.B.n162 0.0209918
R11202 bjt_0.B.n163 bjt_0.B.n65 0.0209918
R11203 bjt_0.B.n168 bjt_0.B.n65 0.0209918
R11204 bjt_0.B.n103 bjt_0.B.n97 0.0209918
R11205 bjt_0.B.n97 bjt_0.B.n33 0.0209918
R11206 bjt_0.B.n197 bjt_0.B.n34 0.0209918
R11207 bjt_0.B.n192 bjt_0.B.n34 0.0201721
R11208 bjt_0.B.n129 bjt_0.B.n128 0.0173033
R11209 bjt_0.B.n143 bjt_0.B.n73 0.0173033
R11210 bjt_0.B.n170 bjt_0.B.n169 0.0173033
R11211 bjt_0.B.n140 bjt_0.B.n139 0.0112346
R11212 bjt_0.B.n84 bjt_0.B.n83 0.0112346
R11213 bjt_0.B.n130 bjt_0.B.n81 0.0112346
R11214 bjt_0.B.n86 bjt_0.B.n85 0.0112346
R11215 bjt_0.B.n142 bjt_0.B.n75 0.0112346
R11216 bjt_0.B.n139 bjt_0.B.n82 0.0112346
R11217 bjt_0.B.n83 bjt_0.B.n82 0.0112346
R11218 bjt_0.B.n130 bjt_0.B.n84 0.0112346
R11219 bjt_0.B.n85 bjt_0.B.n81 0.0112346
R11220 bjt_0.B.n86 bjt_0.B.n75 0.0112346
R11221 bjt_0.B.n172 bjt_0.B.n46 0.0112346
R11222 bjt_0.B.n55 bjt_0.B.n53 0.0112346
R11223 bjt_0.B.n54 bjt_0.B.n51 0.0112346
R11224 bjt_0.B.n170 bjt_0.B.n64 0.0112346
R11225 bjt_0.B.n52 bjt_0.B.n46 0.0112346
R11226 bjt_0.B.n53 bjt_0.B.n52 0.0112346
R11227 bjt_0.B.n55 bjt_0.B.n54 0.0112346
R11228 bjt_0.B.n64 bjt_0.B.n51 0.0112346
R11229 bjt_0.B.n191 bjt_0.B.n40 0.0112346
R11230 bjt_0.B.n177 bjt_0.B.n176 0.0112346
R11231 bjt_0.B.n179 bjt_0.B.n174 0.0112346
R11232 bjt_0.B.n189 bjt_0.B.n178 0.0112346
R11233 bjt_0.B.n188 bjt_0.B.n173 0.0112346
R11234 bjt_0.B.n175 bjt_0.B.n40 0.0112346
R11235 bjt_0.B.n176 bjt_0.B.n175 0.0112346
R11236 bjt_0.B.n179 bjt_0.B.n177 0.0112346
R11237 bjt_0.B.n178 bjt_0.B.n174 0.0112346
R11238 bjt_0.B.n189 bjt_0.B.n188 0.0112346
R11239 bjt_0.B.n198 bjt_0.B.n33 0.0107459
R11240 bjt_0.B.n198 bjt_0.B.n197 0.0107459
R11241 bjt_0.B.n169 bjt_0.B.n50 0.00418852
R11242 digital_0.S1.n41 digital_0.S1.t44 762.783
R11243 digital_0.S1.n41 digital_0.S1.t49 762.783
R11244 digital_0.S1.n37 digital_0.S1.t47 762.783
R11245 digital_0.S1.n37 digital_0.S1.t52 762.783
R11246 digital_0.S1.n42 digital_0.S1.n41 161.3
R11247 digital_0.S1.n38 digital_0.S1.n37 161.3
R11248 digital_0.S1.n4 digital_0.S1.t0 47.7875
R11249 digital_0.S1.n0 digital_0.S1.t55 47.7865
R11250 digital_0.S1.n20 digital_0.S1.t36 47.7865
R11251 digital_0.S1.n0 digital_0.S1.t59 47.6925
R11252 digital_0.S1.n2 digital_0.S1.t26 47.6925
R11253 digital_0.S1.n20 digital_0.S1.t20 47.6925
R11254 digital_0.S1.n4 digital_0.S1.t7 47.6925
R11255 digital_0.S1.n1 digital_0.S1.t9 47.5125
R11256 digital_0.S1.n48 digital_0.S1.t32 43.9066
R11257 digital_0.S1.n13 digital_0.S1.t58 43.7466
R11258 digital_0.S1.n26 digital_0.S1.t10 43.5116
R11259 digital_0.S1.n6 digital_0.S1.t2 43.5116
R11260 digital_0.S1.n32 digital_0.S1.t19 43.3041
R11261 digital_0.S1.n25 digital_0.S1.t13 43.3041
R11262 digital_0.S1.n11 digital_0.S1.t24 43.3041
R11263 digital_0.S1.n27 digital_0.S1.t11 43.2216
R11264 digital_0.S1.n29 digital_0.S1.t37 43.2216
R11265 digital_0.S1.n7 digital_0.S1.t16 43.2216
R11266 digital_0.S1.n9 digital_0.S1.t17 43.2216
R11267 digital_0.S1.n31 digital_0.S1.t18 43.1241
R11268 digital_0.S1.n5 digital_0.S1.t12 43.1241
R11269 digital_0.S1.n12 digital_0.S1.t23 43.1241
R11270 digital_0.S1.n51 digital_0.S1.t5 43.0966
R11271 digital_0.S1.n23 digital_0.S1.t28 43.0966
R11272 digital_0.S1.n15 digital_0.S1.t35 43.0966
R11273 digital_0.S1.n48 digital_0.S1.t57 43.0592
R11274 digital_0.S1.n26 digital_0.S1.t33 43.0416
R11275 digital_0.S1.n28 digital_0.S1.t8 43.0416
R11276 digital_0.S1.n30 digital_0.S1.t29 43.0416
R11277 digital_0.S1.n6 digital_0.S1.t54 43.0416
R11278 digital_0.S1.n8 digital_0.S1.t25 43.0416
R11279 digital_0.S1.n10 digital_0.S1.t56 43.0416
R11280 digital_0.S1.n13 digital_0.S1.t3 43.0416
R11281 digital_0.S1.n32 digital_0.S1.t22 43.0141
R11282 digital_0.S1.n25 digital_0.S1.t15 43.0141
R11283 digital_0.S1.n11 digital_0.S1.t43 43.0141
R11284 digital_0.S1.n52 digital_0.S1.t4 42.9166
R11285 digital_0.S1.n19 digital_0.S1.t27 42.9166
R11286 digital_0.S1.n14 digital_0.S1.t34 42.9166
R11287 digital_0.S1.n31 digital_0.S1.t21 42.8341
R11288 digital_0.S1.n5 digital_0.S1.t14 42.8341
R11289 digital_0.S1.n12 digital_0.S1.t42 42.8341
R11290 digital_0.S1.n48 digital_0.S1 42.8155
R11291 digital_0.S1.n38 digital_0.S1.t48 23.2859
R11292 digital_0.S1.n38 digital_0.S1.t53 23.2859
R11293 digital_0.S1.n42 digital_0.S1.t46 23.2669
R11294 digital_0.S1.n42 digital_0.S1.t51 23.2669
R11295 digital_0.S1.n39 digital_0.S1.n36 18.9359
R11296 digital_0.S1.n39 digital_0.S1.n35 18.9359
R11297 digital_0.S1.n40 digital_0.S1.n34 18.9169
R11298 digital_0.S1 digital_0.S1.n44 18.8194
R11299 digital_0.S1 digital_0.S1.n33 18.7973
R11300 digital_0.S1.n47 digital_0.S1.n46 18.0391
R11301 digital_0.S1.n56 digital_0.S1.n4 11.1039
R11302 digital_0.S1.n21 digital_0.S1.n20 10.3058
R11303 digital_0.S1.n52 digital_0.S1.n51 6.1255
R11304 digital_0.S1.n50 digital_0.S1.n49 6.1255
R11305 digital_0.S1.n15 digital_0.S1.n14 6.1255
R11306 digital_0.S1.n17 digital_0.S1.n16 6.1255
R11307 digital_0.S1.n46 digital_0.S1.t30 4.3505
R11308 digital_0.S1.n46 digital_0.S1.t1 4.3505
R11309 digital_0.S1.n44 digital_0.S1.t31 4.3505
R11310 digital_0.S1.n44 digital_0.S1.t6 4.3505
R11311 digital_0.S1.t53 digital_0.S1.n36 4.3505
R11312 digital_0.S1.n36 digital_0.S1.t41 4.3505
R11313 digital_0.S1.t48 digital_0.S1.n35 4.3505
R11314 digital_0.S1.n35 digital_0.S1.t39 4.3505
R11315 digital_0.S1.n34 digital_0.S1.t40 4.3505
R11316 digital_0.S1.n34 digital_0.S1.t50 4.3505
R11317 digital_0.S1.n33 digital_0.S1.t38 4.3505
R11318 digital_0.S1.n33 digital_0.S1.t45 4.3505
R11319 digital_0.S1.n45 digital_0.S1.n43 3.59185
R11320 digital_0.S1.n21 digital_0.S1.n3 3.14473
R11321 digital_0.S1.n55 digital_0.S1.n54 2.44883
R11322 digital_0.S1.n55 digital_0.S1.n24 2.44883
R11323 digital_0.S1.n23 digital_0.S1.n22 2.44883
R11324 digital_0.S1.n22 digital_0.S1.n19 2.44883
R11325 digital_0.S1 digital_0.S1.n56 2.27213
R11326 digital_0.S1.n49 digital_0.S1.n48 1.9305
R11327 digital_0.S1.n40 digital_0.S1.n39 1.10293
R11328 digital_0.S1.n47 digital_0.S1.n45 0.941788
R11329 digital_0.S1.n3 digital_0.S1.n2 0.873096
R11330 digital_0.S1 digital_0.S1.n3 0.873096
R11331 digital_0.S1 digital_0.S1.n47 0.74103
R11332 digital_0.S1.n14 digital_0.S1.n13 0.7055
R11333 digital_0.S1.n53 digital_0.S1.n30 0.498
R11334 digital_0.S1.n18 digital_0.S1.n10 0.498
R11335 digital_0.S1.n51 digital_0.S1.n50 0.4155
R11336 digital_0.S1.n24 digital_0.S1.n23 0.4155
R11337 digital_0.S1.n16 digital_0.S1.n15 0.4155
R11338 digital_0.S1.n27 digital_0.S1.n26 0.2905
R11339 digital_0.S1.n28 digital_0.S1.n27 0.2905
R11340 digital_0.S1.n29 digital_0.S1.n28 0.2905
R11341 digital_0.S1.n30 digital_0.S1.n29 0.2905
R11342 digital_0.S1.n7 digital_0.S1.n6 0.2905
R11343 digital_0.S1.n8 digital_0.S1.n7 0.2905
R11344 digital_0.S1.n9 digital_0.S1.n8 0.2905
R11345 digital_0.S1.n10 digital_0.S1.n9 0.2905
R11346 digital_0.S1.n1 digital_0.S1.n0 0.274538
R11347 digital_0.S1.n2 digital_0.S1.n1 0.274538
R11348 digital_0.S1.n54 digital_0.S1.n53 0.208
R11349 digital_0.S1.n53 digital_0.S1.n52 0.208
R11350 digital_0.S1.n18 digital_0.S1.n17 0.208
R11351 digital_0.S1.n19 digital_0.S1.n18 0.208
R11352 digital_0.S1.n39 digital_0.S1.n38 0.190155
R11353 digital_0.S1.n22 digital_0.S1.n21 0.1805
R11354 digital_0.S1.n56 digital_0.S1.n55 0.1805
R11355 digital_0.S1.n45 digital_0.S1 0.161485
R11356 digital_0.S1.n40 digital_0.S1 0.120065
R11357 digital_0.S1.n49 digital_0.S1.n32 0.083
R11358 digital_0.S1.n50 digital_0.S1.n31 0.083
R11359 digital_0.S1.n54 digital_0.S1.n25 0.083
R11360 digital_0.S1.n24 digital_0.S1.n5 0.083
R11361 digital_0.S1.n17 digital_0.S1.n11 0.083
R11362 digital_0.S1.n16 digital_0.S1.n12 0.083
R11363 digital_0.S1.n43 digital_0.S1.n40 0.0768889
R11364 digital_0.S1.n43 digital_0.S1.n42 0.0768889
R11365 DVSS.n45 DVSS.n8 8471
R11366 DVSS.n28 DVSS.n4 8471
R11367 DVSS.n61 DVSS.n4 8471
R11368 DVSS.n59 DVSS.n8 8471
R11369 DVSS.n39 DVSS.n24 5886.82
R11370 DVSS.n24 DVSS.n3 5886.82
R11371 DVSS.n53 DVSS.n11 5886.82
R11372 DVSS.n53 DVSS.n12 5886.82
R11373 DVSS.n51 DVSS.n25 5886.82
R11374 DVSS.n51 DVSS.n9 5886.82
R11375 DVSS.n37 DVSS.n29 3870.47
R11376 DVSS.n37 DVSS.n31 3870.47
R11377 DVSS.n33 DVSS.n29 3870.47
R11378 DVSS.n33 DVSS.n31 3870.47
R11379 DVSS.n22 DVSS.n14 3870.47
R11380 DVSS.n22 DVSS.n16 3870.47
R11381 DVSS.n18 DVSS.n14 3870.47
R11382 DVSS.n18 DVSS.n16 3870.47
R11383 DVSS.n45 DVSS.n25 2584.18
R11384 DVSS.n47 DVSS.n25 2584.18
R11385 DVSS.n47 DVSS.n11 2584.18
R11386 DVSS.n44 DVSS.n11 2584.18
R11387 DVSS.n44 DVSS.n39 2584.18
R11388 DVSS.n39 DVSS.n28 2584.18
R11389 DVSS.n59 DVSS.n9 2584.18
R11390 DVSS.n9 DVSS.n6 2584.18
R11391 DVSS.n12 DVSS.n6 2584.18
R11392 DVSS.n12 DVSS.n7 2584.18
R11393 DVSS.n7 DVSS.n3 2584.18
R11394 DVSS.n61 DVSS.n3 2584.18
R11395 DVSS.n27 DVSS.n26 550.4
R11396 DVSS.n41 DVSS.n40 550.4
R11397 DVSS.n58 DVSS 549.271
R11398 DVSS.n54 DVSS.n10 382.495
R11399 DVSS.n50 DVSS.n49 382.495
R11400 DVSS.n42 DVSS.n0 382.495
R11401 DVSS.n55 DVSS 381.365
R11402 DVSS.n57 DVSS 381.365
R11403 DVSS DVSS.n63 381.365
R11404 DVSS.n40 DVSS.n2 338.825
R11405 DVSS.n36 DVSS.n32 251.482
R11406 DVSS.n36 DVSS.n35 251.482
R11407 DVSS.n34 DVSS.n32 251.482
R11408 DVSS.n21 DVSS.n17 251.482
R11409 DVSS.n19 DVSS.n17 251.482
R11410 DVSS.n20 DVSS.n19 251.482
R11411 DVSS.n35 DVSS 214.965
R11412 DVSS DVSS.n20 214.965
R11413 DVSS.n62 DVSS.n2 211.577
R11414 DVSS.t2 DVSS.t5 178.518
R11415 DVSS.t9 DVSS.t7 178.518
R11416 DVSS.t6 DVSS.t8 178.518
R11417 DVSS.t1 DVSS.t4 178.518
R11418 DVSS.n49 DVSS.n27 167.906
R11419 DVSS.n49 DVSS.n48 167.906
R11420 DVSS.n48 DVSS.n10 167.906
R11421 DVSS.n43 DVSS.n10 167.906
R11422 DVSS.n43 DVSS.n42 167.906
R11423 DVSS.n42 DVSS.n41 167.906
R11424 DVSS.n58 DVSS.n57 167.906
R11425 DVSS.n57 DVSS.n56 167.906
R11426 DVSS.n56 DVSS.n55 167.906
R11427 DVSS.n55 DVSS.n1 167.906
R11428 DVSS.n63 DVSS.n1 167.906
R11429 DVSS.n63 DVSS.n62 167.906
R11430 DVSS.n38 DVSS.t5 148.594
R11431 DVSS.t7 DVSS.n13 148.594
R11432 DVSS.n23 DVSS.t8 148.594
R11433 DVSS.n30 DVSS.t2 133.114
R11434 DVSS.n15 DVSS.t1 133.114
R11435 DVSS.n52 DVSS.n13 114.54
R11436 DVSS.n52 DVSS.n23 114.54
R11437 DVSS.n19 DVSS.n18 97.5005
R11438 DVSS.n18 DVSS.n5 97.5005
R11439 DVSS.n22 DVSS.n21 97.5005
R11440 DVSS.n23 DVSS.n22 97.5005
R11441 DVSS.n34 DVSS.n33 97.5005
R11442 DVSS.n33 DVSS.n13 97.5005
R11443 DVSS.n37 DVSS.n36 97.5005
R11444 DVSS.n38 DVSS.n37 97.5005
R11445 DVSS DVSS.n5 93.9029
R11446 DVSS.t0 DVSS.t9 71.2013
R11447 DVSS.t3 DVSS.t6 71.2013
R11448 DVSS.n30 DVSS.t0 61.9142
R11449 DVSS.n15 DVSS.t3 61.9142
R11450 DVSS.t4 DVSS 54.6909
R11451 DVSS.n20 DVSS.n16 48.7505
R11452 DVSS.n16 DVSS.n15 48.7505
R11453 DVSS.n17 DVSS.n14 48.7505
R11454 DVSS.n15 DVSS.n14 48.7505
R11455 DVSS.n35 DVSS.n31 48.7505
R11456 DVSS.n31 DVSS.n30 48.7505
R11457 DVSS.n32 DVSS.n29 48.7505
R11458 DVSS.n30 DVSS.n29 48.7505
R11459 DVSS.n45 DVSS.n27 48.7505
R11460 DVSS.n46 DVSS.n45 48.7505
R11461 DVSS.n48 DVSS.n47 48.7505
R11462 DVSS.n47 DVSS.n46 48.7505
R11463 DVSS.n44 DVSS.n43 48.7505
R11464 DVSS.n46 DVSS.n44 48.7505
R11465 DVSS.n41 DVSS.n28 48.7505
R11466 DVSS.n46 DVSS.n28 48.7505
R11467 DVSS.n62 DVSS.n61 48.7505
R11468 DVSS.n61 DVSS.n60 48.7505
R11469 DVSS.n7 DVSS.n1 48.7505
R11470 DVSS.n60 DVSS.n7 48.7505
R11471 DVSS.n56 DVSS.n6 48.7505
R11472 DVSS.n60 DVSS.n6 48.7505
R11473 DVSS.n59 DVSS.n58 48.7505
R11474 DVSS.n60 DVSS.n59 48.7505
R11475 DVSS DVSS.n34 36.5181
R11476 DVSS.n21 DVSS 36.5181
R11477 DVSS.n46 DVSS.n38 30.9573
R11478 DVSS.n60 DVSS.n5 30.9573
R11479 DVSS.n2 DVSS 24.4519
R11480 DVSS.n54 DVSS.n53 20.1729
R11481 DVSS.n53 DVSS.n52 20.1729
R11482 DVSS.n51 DVSS.n50 20.1729
R11483 DVSS.n52 DVSS.n51 20.1729
R11484 DVSS.n26 DVSS.n8 20.1729
R11485 DVSS.n52 DVSS.n8 20.1729
R11486 DVSS.n24 DVSS.n0 20.1729
R11487 DVSS.n52 DVSS.n24 20.1729
R11488 DVSS.n40 DVSS.n4 20.1729
R11489 DVSS.n52 DVSS.n4 20.1729
R11490 DVSS DVSS.n54 1.12991
R11491 DVSS.n50 DVSS 1.12991
R11492 DVSS.n26 DVSS 1.12991
R11493 DVSS DVSS.n0 1.12991
R11494 TRIM3.t2 TRIM3 190.643
R11495 TRIM3 TRIM3.t3 190.609
R11496 TRIM3.t1 TRIM3.n1 190.585
R11497 TRIM3.n1 TRIM3.t0 190.585
R11498 TRIM3.t0 TRIM3.n0 119.778
R11499 TRIM3.n0 TRIM3.t2 119.778
R11500 TRIM3.t3 TRIM3.n2 119.778
R11501 TRIM3.n2 TRIM3.t1 119.778
R11502 TRIM3.n1 TRIM3 20.1784
R11503 TRIM3.n2 TRIM3.n0 19.6878
R11504 digital_0.S3.n9 digital_0.S3.t17 762.783
R11505 digital_0.S3.n9 digital_0.S3.t12 762.783
R11506 digital_0.S3.n5 digital_0.S3.t15 762.783
R11507 digital_0.S3.n5 digital_0.S3.t20 762.783
R11508 digital_0.S3.n10 digital_0.S3.n9 161.3
R11509 digital_0.S3.n6 digital_0.S3.n5 161.3
R11510 digital_0.S3.n0 digital_0.S3.t8 57.4691
R11511 digital_0.S3.n19 digital_0.S3.t10 54.9333
R11512 digital_0.S3.n17 digital_0.S3.t22 54.8559
R11513 digital_0.S3.n16 digital_0.S3.t7 53.9629
R11514 digital_0.S3.n17 digital_0.S3.t4 51.4723
R11515 digital_0.S3.n19 digital_0.S3.t23 50.9842
R11516 digital_0.S3.n16 digital_0.S3 37.4963
R11517 digital_0.S3.n6 digital_0.S3.t16 23.2859
R11518 digital_0.S3.n6 digital_0.S3.t21 23.2859
R11519 digital_0.S3.n10 digital_0.S3.t19 23.2669
R11520 digital_0.S3.n10 digital_0.S3.t14 23.2669
R11521 digital_0.S3.n7 digital_0.S3.n4 18.9359
R11522 digital_0.S3.n7 digital_0.S3.n3 18.9359
R11523 digital_0.S3.n8 digital_0.S3.n2 18.9169
R11524 digital_0.S3 digital_0.S3.n12 18.8194
R11525 digital_0.S3 digital_0.S3.n1 18.7973
R11526 digital_0.S3.n15 digital_0.S3.n14 18.0391
R11527 digital_0.S3.n14 digital_0.S3.t0 4.3505
R11528 digital_0.S3.n14 digital_0.S3.t1 4.3505
R11529 digital_0.S3.n12 digital_0.S3.t3 4.3505
R11530 digital_0.S3.n12 digital_0.S3.t2 4.3505
R11531 digital_0.S3.t21 digital_0.S3.n4 4.3505
R11532 digital_0.S3.n4 digital_0.S3.t9 4.3505
R11533 digital_0.S3.t16 digital_0.S3.n3 4.3505
R11534 digital_0.S3.n3 digital_0.S3.t6 4.3505
R11535 digital_0.S3.n2 digital_0.S3.t11 4.3505
R11536 digital_0.S3.n2 digital_0.S3.t13 4.3505
R11537 digital_0.S3.n1 digital_0.S3.t5 4.3505
R11538 digital_0.S3.n1 digital_0.S3.t18 4.3505
R11539 digital_0.S3.n13 digital_0.S3.n11 3.58944
R11540 digital_0.S3.n21 digital_0.S3.n16 2.96885
R11541 digital_0.S3.n20 digital_0.S3.n18 1.59711
R11542 digital_0.S3.n8 digital_0.S3.n7 1.10293
R11543 digital_0.S3.n15 digital_0.S3.n13 0.941788
R11544 digital_0.S3 digital_0.S3.n0 0.940018
R11545 digital_0.S3 digital_0.S3.n21 0.89017
R11546 digital_0.S3.n20 digital_0.S3.n19 0.771744
R11547 digital_0.S3.n18 digital_0.S3.n17 0.771744
R11548 digital_0.S3 digital_0.S3.n15 0.722091
R11549 digital_0.S3.n7 digital_0.S3.n6 0.190155
R11550 digital_0.S3.n21 digital_0.S3.n20 0.171
R11551 digital_0.S3.n18 digital_0.S3.n0 0.171
R11552 digital_0.S3.n13 digital_0.S3 0.161485
R11553 digital_0.S3.n8 digital_0.S3 0.120065
R11554 digital_0.S3.n11 digital_0.S3.n8 0.0768889
R11555 digital_0.S3.n11 digital_0.S3.n10 0.0768889
R11556 digital_0.D3.n9 digital_0.D3.t2 762.783
R11557 digital_0.D3.n9 digital_0.D3.t7 762.783
R11558 digital_0.D3.n6 digital_0.D3.t0 762.783
R11559 digital_0.D3.n6 digital_0.D3.t5 762.783
R11560 digital_0.D3.n10 digital_0.D3.n9 161.3
R11561 digital_0.D3.n7 digital_0.D3.n6 161.3
R11562 digital_0.D3 digital_0.D3.t14 60.3223
R11563 digital_0.D3.n1 digital_0.D3.t16 53.6908
R11564 digital_0.D3.n0 digital_0.D3.t15 42.3691
R11565 digital_0.D3.n10 digital_0.D3.t4 23.2859
R11566 digital_0.D3.n10 digital_0.D3.t9 23.2859
R11567 digital_0.D3.n7 digital_0.D3.t1 23.2859
R11568 digital_0.D3.n7 digital_0.D3.t6 23.2859
R11569 digital_0.D3.n13 digital_0.D3.n12 20.3847
R11570 digital_0.D3.n11 digital_0.D3.n3 18.9359
R11571 digital_0.D3.n8 digital_0.D3.n5 18.9359
R11572 digital_0.D3.n8 digital_0.D3.n4 18.9359
R11573 digital_0.D3.n12 digital_0.D3.n2 17.6641
R11574 digital_0.D3.n1 digital_0.D3.n0 17.55
R11575 digital_0.D3 digital_0.D3.n13 4.97324
R11576 digital_0.D3.n2 digital_0.D3.t10 4.3505
R11577 digital_0.D3.n2 digital_0.D3.t3 4.3505
R11578 digital_0.D3.n3 digital_0.D3.t12 4.3505
R11579 digital_0.D3.n3 digital_0.D3.t8 4.3505
R11580 digital_0.D3.t6 digital_0.D3.n5 4.3505
R11581 digital_0.D3.n5 digital_0.D3.t13 4.3505
R11582 digital_0.D3.t1 digital_0.D3.n4 4.3505
R11583 digital_0.D3.n4 digital_0.D3.t11 4.3505
R11584 digital_0.D3.n11 digital_0.D3.n8 1.11257
R11585 digital_0.D3.n12 digital_0.D3 0.752915
R11586 digital_0.D3.n12 digital_0.D3 0.715778
R11587 digital_0.D3.n0 digital_0.D3 0.454827
R11588 digital_0.D3.n13 digital_0.D3.n1 0.27253
R11589 digital_0.D3.n8 digital_0.D3.n7 0.190155
R11590 digital_0.D3.n11 digital_0.D3.n10 0.190155
R11591 digital_0.D3 digital_0.D3.n11 0.139087
R11592 resistor_op_tt_0.C.n10 resistor_op_tt_0.C.t8 402.695
R11593 resistor_op_tt_0.C.n1 resistor_op_tt_0.C.t5 402.695
R11594 resistor_op_tt_0.C.n17 resistor_op_tt_0.C.t10 371.644
R11595 resistor_op_tt_0.C.n14 resistor_op_tt_0.C.t13 371.644
R11596 resistor_op_tt_0.C.t9 resistor_op_tt_0.C.n10 227.323
R11597 resistor_op_tt_0.C.n1 resistor_op_tt_0.C.t7 227.323
R11598 resistor_op_tt_0.C.n12 resistor_op_tt_0.C.n11 199.65
R11599 resistor_op_tt_0.C.n3 resistor_op_tt_0.C.n2 199.65
R11600 resistor_op_tt_0.C.n17 resistor_op_tt_0.C.t12 115.525
R11601 resistor_op_tt_0.C.t14 resistor_op_tt_0.C.n14 115.525
R11602 resistor_op_tt_0.C.n19 resistor_op_tt_0.C.n18 97.1505
R11603 resistor_op_tt_0.C.n16 resistor_op_tt_0.C.n15 97.1505
R11604 resistor_op_tt_0.C.n23 resistor_op_tt_0.C.t0 42.3701
R11605 resistor_op_tt_0.C.n0 resistor_op_tt_0.C.t4 42.3691
R11606 resistor_op_tt_0.C.n11 resistor_op_tt_0.C.t9 28.5655
R11607 resistor_op_tt_0.C.n11 resistor_op_tt_0.C.t15 28.5655
R11608 resistor_op_tt_0.C.n2 resistor_op_tt_0.C.t3 28.5655
R11609 resistor_op_tt_0.C.n2 resistor_op_tt_0.C.t6 28.5655
R11610 resistor_op_tt_0.C.n21 resistor_op_tt_0.C.n13 19.9821
R11611 resistor_op_tt_0.C.n18 resistor_op_tt_0.C.t1 19.3338
R11612 resistor_op_tt_0.C.n18 resistor_op_tt_0.C.t11 19.3338
R11613 resistor_op_tt_0.C.n15 resistor_op_tt_0.C.t14 19.3338
R11614 resistor_op_tt_0.C.n15 resistor_op_tt_0.C.t2 19.3338
R11615 resistor_op_tt_0.C.n6 resistor_op_tt_0.C.n5 16.2244
R11616 resistor_op_tt_0.C.n5 resistor_op_tt_0.C.n4 15.0885
R11617 resistor_op_tt_0.C.n7 resistor_op_tt_0.C.n6 15.0885
R11618 resistor_op_tt_0.C.n8 resistor_op_tt_0.C 13.1344
R11619 resistor_op_tt_0.C.n7 resistor_op_tt_0.C.t19 11.5219
R11620 resistor_op_tt_0.C.n6 resistor_op_tt_0.C.t17 11.5219
R11621 resistor_op_tt_0.C.n5 resistor_op_tt_0.C.t18 11.5219
R11622 resistor_op_tt_0.C.n4 resistor_op_tt_0.C.t16 11.5219
R11623 resistor_op_tt_0.C.n13 resistor_op_tt_0.C 10.4548
R11624 resistor_op_tt_0.C.n21 resistor_op_tt_0.C.n20 9.4191
R11625 resistor_op_tt_0.C.n20 resistor_op_tt_0.C 6.02835
R11626 resistor_op_tt_0.C.n9 resistor_op_tt_0.C.n8 5.97406
R11627 resistor_op_tt_0.C resistor_op_tt_0.C.n16 4.06088
R11628 resistor_op_tt_0.C.n8 resistor_op_tt_0.C.n7 2.87144
R11629 resistor_op_tt_0.C.n22 resistor_op_tt_0.C.n0 2.76169
R11630 resistor_op_tt_0.C.n23 resistor_op_tt_0.C.n22 2.58877
R11631 resistor_op_tt_0.C.n20 resistor_op_tt_0.C.n19 2.2505
R11632 resistor_op_tt_0.C.n9 resistor_op_tt_0.C.n3 2.2505
R11633 resistor_op_tt_0.C.n13 resistor_op_tt_0.C.n12 2.2505
R11634 resistor_op_tt_0.C resistor_op_tt_0.C.n0 1.038
R11635 resistor_op_tt_0.C.n19 resistor_op_tt_0.C.n17 0.64517
R11636 resistor_op_tt_0.C.n16 resistor_op_tt_0.C.n14 0.64517
R11637 resistor_op_tt_0.C.n12 resistor_op_tt_0.C.n10 0.610083
R11638 resistor_op_tt_0.C.n3 resistor_op_tt_0.C.n1 0.610083
R11639 resistor_op_tt_0.C resistor_op_tt_0.C.n23 0.573
R11640 resistor_op_tt_0.C resistor_op_tt_0.C.n9 0.291365
R11641 resistor_op_tt_0.C.n22 resistor_op_tt_0.C.n21 0.268208
R11642 resistor_op_tt_0.C.n4 resistor_op_tt_0.C 0.199458
R11643 pmos_iptat_0.G.t28 pmos_iptat_0.G.t29 516.596
R11644 pmos_iptat_0.G.n19 pmos_iptat_0.G.t2 402.716
R11645 pmos_iptat_0.G.n8 pmos_iptat_0.G.t9 402.695
R11646 pmos_iptat_0.G.n14 pmos_iptat_0.G.t4 402.695
R11647 pmos_iptat_0.G.n31 pmos_iptat_0.G.t15 402.695
R11648 pmos_iptat_0.G.n3 pmos_iptat_0.G.t6 387.759
R11649 pmos_iptat_0.G.n2 pmos_iptat_0.G.t12 387.759
R11650 pmos_iptat_0.G.t24 pmos_iptat_0.G.t26 376.724
R11651 pmos_iptat_0.G.t26 pmos_iptat_0.G.t23 376.724
R11652 pmos_iptat_0.G.t25 pmos_iptat_0.G.t23 376.724
R11653 pmos_iptat_0.G.n8 pmos_iptat_0.G.t11 227.323
R11654 pmos_iptat_0.G.t5 pmos_iptat_0.G.n14 227.323
R11655 pmos_iptat_0.G.n31 pmos_iptat_0.G.t17 227.323
R11656 pmos_iptat_0.G.t3 pmos_iptat_0.G.n19 227.322
R11657 pmos_iptat_0.G.n32 pmos_iptat_0.G.n30 199.65
R11658 pmos_iptat_0.G.n10 pmos_iptat_0.G.n9 199.65
R11659 pmos_iptat_0.G.n21 pmos_iptat_0.G.n20 199.65
R11660 pmos_iptat_0.G.n16 pmos_iptat_0.G.n15 199.65
R11661 pmos_iptat_0.G.n0 pmos_iptat_0.G.t1 83.7522
R11662 pmos_iptat_0.G.n1 pmos_iptat_0.G.t0 83.7522
R11663 pmos_iptat_0.G.n0 pmos_iptat_0.G.t7 83.7172
R11664 pmos_iptat_0.G.n1 pmos_iptat_0.G.t14 83.7172
R11665 pmos_iptat_0.G.n3 pmos_iptat_0.G.t8 82.8128
R11666 pmos_iptat_0.G.n2 pmos_iptat_0.G.t13 82.8128
R11667 pmos_iptat_0.G.t25 pmos_iptat_0.G.t24 31.1858
R11668 pmos_iptat_0.G.n30 pmos_iptat_0.G.t20 28.5655
R11669 pmos_iptat_0.G.n30 pmos_iptat_0.G.t16 28.5655
R11670 pmos_iptat_0.G.n9 pmos_iptat_0.G.t19 28.5655
R11671 pmos_iptat_0.G.n9 pmos_iptat_0.G.t10 28.5655
R11672 pmos_iptat_0.G.n20 pmos_iptat_0.G.t3 28.5655
R11673 pmos_iptat_0.G.n20 pmos_iptat_0.G.t21 28.5655
R11674 pmos_iptat_0.G.n15 pmos_iptat_0.G.t5 28.5655
R11675 pmos_iptat_0.G.n15 pmos_iptat_0.G.t18 28.5655
R11676 pmos_iptat_0.G pmos_iptat_0.G.n1 22.8082
R11677 pmos_iptat_0.G.n36 pmos_iptat_0.G.n5 22.7477
R11678 pmos_iptat_0.G.n22 pmos_iptat_0.G.n11 20.4188
R11679 pmos_iptat_0.G.n5 pmos_iptat_0.G.t27 14.4193
R11680 pmos_iptat_0.G.n34 pmos_iptat_0.G.n33 13.7577
R11681 pmos_iptat_0.G.n35 pmos_iptat_0.G.t28 12.765
R11682 pmos_iptat_0.G.t26 pmos_iptat_0.G.n26 11.5219
R11683 pmos_iptat_0.G.t23 pmos_iptat_0.G.n12 11.5219
R11684 pmos_iptat_0.G.n27 pmos_iptat_0.G.t25 11.5219
R11685 pmos_iptat_0.G.t24 pmos_iptat_0.G.n23 11.5219
R11686 pmos_iptat_0.G.t25 pmos_iptat_0.G.n7 11.5219
R11687 pmos_iptat_0.G.n24 pmos_iptat_0.G.t23 11.5219
R11688 pmos_iptat_0.G.t26 pmos_iptat_0.G.n25 11.5219
R11689 pmos_iptat_0.G.t24 pmos_iptat_0.G.n13 11.5219
R11690 pmos_iptat_0.G.n37 pmos_iptat_0.G.t29 11.5219
R11691 pmos_iptat_0.G.n5 pmos_iptat_0.G.n4 8.86552
R11692 pmos_iptat_0.G.n26 pmos_iptat_0.G.n12 5.59289
R11693 pmos_iptat_0.G.n25 pmos_iptat_0.G.n24 5.59289
R11694 pmos_iptat_0.G.n27 pmos_iptat_0.G.n12 5.43549
R11695 pmos_iptat_0.G.n26 pmos_iptat_0.G.n23 5.43549
R11696 pmos_iptat_0.G.n24 pmos_iptat_0.G.n7 5.43549
R11697 pmos_iptat_0.G.n25 pmos_iptat_0.G.n13 5.43549
R11698 pmos_iptat_0.G.n17 pmos_iptat_0.G.n6 3.70483
R11699 pmos_iptat_0.G.n34 pmos_iptat_0.G.n6 2.58223
R11700 pmos_iptat_0.G.n4 pmos_iptat_0.G.n0 2.2505
R11701 pmos_iptat_0.G.n22 pmos_iptat_0.G.n21 2.2505
R11702 pmos_iptat_0.G.n11 pmos_iptat_0.G.n10 2.2505
R11703 pmos_iptat_0.G.n17 pmos_iptat_0.G.n16 2.2505
R11704 pmos_iptat_0.G.n33 pmos_iptat_0.G.n32 2.2505
R11705 pmos_iptat_0.G.n36 pmos_iptat_0.G.n35 2.238
R11706 pmos_iptat_0.G.n28 pmos_iptat_0.G.n11 1.8484
R11707 pmos_iptat_0.G.n33 pmos_iptat_0.G.n29 1.8484
R11708 pmos_iptat_0.G.n18 pmos_iptat_0.G.n17 1.8484
R11709 pmos_iptat_0.G pmos_iptat_0.G.n22 1.82411
R11710 pmos_iptat_0.G.n28 pmos_iptat_0.G.n27 1.37277
R11711 pmos_iptat_0.G.n23 pmos_iptat_0.G 1.37277
R11712 pmos_iptat_0.G.n29 pmos_iptat_0.G.n7 1.37277
R11713 pmos_iptat_0.G.n18 pmos_iptat_0.G.n13 1.37277
R11714 pmos_iptat_0.G pmos_iptat_0.G.t22 1.37035
R11715 pmos_iptat_0.G.n37 pmos_iptat_0.G.n36 1.24361
R11716 pmos_iptat_0.G pmos_iptat_0.G.n37 1.19762
R11717 pmos_iptat_0.G pmos_iptat_0.G.n18 1.00708
R11718 pmos_iptat_0.G.n29 pmos_iptat_0.G.n28 0.9828
R11719 pmos_iptat_0.G.n1 pmos_iptat_0.G.n2 0.697467
R11720 pmos_iptat_0.G.n0 pmos_iptat_0.G.n3 0.697467
R11721 pmos_iptat_0.G.n21 pmos_iptat_0.G.n19 0.611736
R11722 pmos_iptat_0.G.n10 pmos_iptat_0.G.n8 0.610083
R11723 pmos_iptat_0.G.n16 pmos_iptat_0.G.n14 0.610083
R11724 pmos_iptat_0.G.n32 pmos_iptat_0.G.n31 0.610083
R11725 pmos_iptat_0.G.t27 pmos_iptat_0.G 0.605135
R11726 pmos_iptat_0.G.n4 pmos_iptat_0.G 0.296173
R11727 pmos_iptat_0.G.n36 pmos_iptat_0.G.n6 0.234474
R11728 pmos_iptat_0.G.n35 pmos_iptat_0.G.n34 0.234474
R11729 pmos_startup_0.D4 pmos_startup_0.D4.t0 402.317
R11730 pmos_startup_0.D4.t1 pmos_startup_0.D4 227.351
R11731 pmos_startup_0.D4 pmos_startup_0.D4.n2 199.68
R11732 pmos_startup_0.D4 pmos_startup_0.D4.t6 152.062
R11733 pmos_startup_0.D4.n1 pmos_startup_0.D4 85.4335
R11734 pmos_startup_0.D4.n0 pmos_startup_0.D4.t3 37.3555
R11735 pmos_startup_0.D4.n0 pmos_startup_0.D4.t4 37.3555
R11736 pmos_startup_0.D4.n1 pmos_startup_0.D4.t5 37.3555
R11737 pmos_startup_0.D4.t6 pmos_startup_0.D4.n1 37.3555
R11738 pmos_startup_0.D4.n1 pmos_startup_0.D4.n0 34.9455
R11739 pmos_startup_0.D4.n2 pmos_startup_0.D4.t1 28.5655
R11740 pmos_startup_0.D4.n2 pmos_startup_0.D4.t2 28.5655
R11741 pmos_startup_0.D3.n1 pmos_startup_0.D3.t5 402.317
R11742 pmos_startup_0.D3.n4 pmos_startup_0.D3.t9 387.824
R11743 pmos_startup_0.D3.n12 pmos_startup_0.D3.t7 387.824
R11744 pmos_startup_0.D3.n16 pmos_startup_0.D3.t0 387.824
R11745 pmos_startup_0.D3.n8 pmos_startup_0.D3.t2 387.824
R11746 pmos_startup_0.D3.n1 pmos_startup_0.D3.t6 227.351
R11747 pmos_startup_0.D3.n3 pmos_startup_0.D3.n0 199.65
R11748 pmos_startup_0.D3.t8 pmos_startup_0.D3.n12 82.8079
R11749 pmos_startup_0.D3.n16 pmos_startup_0.D3.t1 82.8079
R11750 pmos_startup_0.D3.n8 pmos_startup_0.D3.t4 82.8079
R11751 pmos_startup_0.D3.n4 pmos_startup_0.D3.t11 82.8079
R11752 pmos_startup_0.D3.n6 pmos_startup_0.D3.n5 66.3172
R11753 pmos_startup_0.D3.n14 pmos_startup_0.D3.n13 66.3172
R11754 pmos_startup_0.D3.n17 pmos_startup_0.D3.n15 66.3172
R11755 pmos_startup_0.D3.n9 pmos_startup_0.D3.n7 66.3172
R11756 pmos_startup_0.D3.t6 pmos_startup_0.D3.n3 28.5655
R11757 pmos_startup_0.D3.n3 pmos_startup_0.D3.t13 28.5655
R11758 pmos_startup_0.D3.n5 pmos_startup_0.D3.t15 17.4005
R11759 pmos_startup_0.D3.n5 pmos_startup_0.D3.t10 17.4005
R11760 pmos_startup_0.D3.n13 pmos_startup_0.D3.t8 17.4005
R11761 pmos_startup_0.D3.n13 pmos_startup_0.D3.t17 17.4005
R11762 pmos_startup_0.D3.t1 pmos_startup_0.D3.n15 17.4005
R11763 pmos_startup_0.D3.n15 pmos_startup_0.D3.t16 17.4005
R11764 pmos_startup_0.D3.n7 pmos_startup_0.D3.t14 17.4005
R11765 pmos_startup_0.D3.n7 pmos_startup_0.D3.t3 17.4005
R11766 pmos_startup_0.D3.n2 pmos_startup_0.D3.t18 17.1143
R11767 pmos_startup_0.D3.n11 pmos_startup_0.D3.n0 16.1238
R11768 pmos_startup_0.D3.n2 pmos_startup_0.D3.t12 11.5219
R11769 pmos_startup_0.D3.n1 pmos_startup_0.D3.n0 0.581685
R11770 pmos_startup_0.D3 pmos_startup_0.D3.n18 4.5005
R11771 pmos_startup_0.D3.n11 pmos_startup_0.D3.n10 4.5005
R11772 pmos_startup_0.D3 pmos_startup_0.D3.n2 2.72479
R11773 pmos_startup_0.D3 pmos_startup_0.D3.n11 0.896333
R11774 pmos_startup_0.D3.n6 pmos_startup_0.D3.n4 0.612666
R11775 pmos_startup_0.D3.n14 pmos_startup_0.D3.n12 0.612666
R11776 pmos_startup_0.D3.n17 pmos_startup_0.D3.n16 0.612666
R11777 pmos_startup_0.D3.n9 pmos_startup_0.D3.n8 0.612666
R11778 pmos_startup_0.D3.n0 pmos_startup_0.D3 0.275849
R11779 pmos_startup_0.D3.n18 pmos_startup_0.D3.n14 0.217727
R11780 pmos_startup_0.D3.n18 pmos_startup_0.D3.n17 0.217727
R11781 pmos_startup_0.D3.n10 pmos_startup_0.D3.n9 0.217727
R11782 pmos_startup_0.D3.n10 pmos_startup_0.D3.n6 0.217727
R11783 pmos_current_bgr_2_0.D4.n16 pmos_current_bgr_2_0.D4.t14 402.51
R11784 pmos_current_bgr_2_0.D4.n7 pmos_current_bgr_2_0.D4.t9 402.51
R11785 pmos_current_bgr_2_0.D4.n5 pmos_current_bgr_2_0.D4.t6 387.759
R11786 pmos_current_bgr_2_0.D4.n4 pmos_current_bgr_2_0.D4.t11 387.759
R11787 pmos_current_bgr_2_0.D4.t10 pmos_current_bgr_2_0.D4.n7 227.337
R11788 pmos_current_bgr_2_0.D4.n16 pmos_current_bgr_2_0.D4.t16 227.337
R11789 pmos_current_bgr_2_0.D4.n10 pmos_current_bgr_2_0.D4.n8 200.034
R11790 pmos_current_bgr_2_0.D4.n15 pmos_current_bgr_2_0.D4.n3 200.034
R11791 pmos_current_bgr_2_0.D4.n0 pmos_current_bgr_2_0.D4.t1 83.7522
R11792 pmos_current_bgr_2_0.D4.n1 pmos_current_bgr_2_0.D4.t0 83.7522
R11793 pmos_current_bgr_2_0.D4.n0 pmos_current_bgr_2_0.D4.t7 83.7172
R11794 pmos_current_bgr_2_0.D4.n1 pmos_current_bgr_2_0.D4.t13 83.7172
R11795 pmos_current_bgr_2_0.D4.n5 pmos_current_bgr_2_0.D4.t8 82.8128
R11796 pmos_current_bgr_2_0.D4.n4 pmos_current_bgr_2_0.D4.t12 82.8128
R11797 pmos_current_bgr_2_0.D4.n8 pmos_current_bgr_2_0.D4.t10 28.5655
R11798 pmos_current_bgr_2_0.D4.n8 pmos_current_bgr_2_0.D4.t3 28.5655
R11799 pmos_current_bgr_2_0.D4.n3 pmos_current_bgr_2_0.D4.t5 28.5655
R11800 pmos_current_bgr_2_0.D4.n3 pmos_current_bgr_2_0.D4.t15 28.5655
R11801 pmos_current_bgr_2_0.D4.n6 pmos_current_bgr_2_0.D4.n1 13.1825
R11802 pmos_current_bgr_2_0.D4 pmos_current_bgr_2_0.D4.n17 12.5576
R11803 pmos_current_bgr_2_0.D4.n14 pmos_current_bgr_2_0.D4.t4 11.5219
R11804 pmos_current_bgr_2_0.D4.n13 pmos_current_bgr_2_0.D4.t18 11.5219
R11805 pmos_current_bgr_2_0.D4.n2 pmos_current_bgr_2_0.D4.t17 11.5219
R11806 pmos_current_bgr_2_0.D4.n9 pmos_current_bgr_2_0.D4.t2 11.5219
R11807 pmos_current_bgr_2_0.D4.n13 pmos_current_bgr_2_0.D4.n12 8.96517
R11808 pmos_current_bgr_2_0.D4.n12 pmos_current_bgr_2_0.D4.n6 8.79224
R11809 pmos_current_bgr_2_0.D4.n12 pmos_current_bgr_2_0.D4.n11 5.92985
R11810 pmos_current_bgr_2_0.D4.n9 pmos_current_bgr_2_0.D4.n2 5.59289
R11811 pmos_current_bgr_2_0.D4.n14 pmos_current_bgr_2_0.D4.n13 5.59289
R11812 pmos_current_bgr_2_0.D4.n10 pmos_current_bgr_2_0.D4.n9 2.7967
R11813 pmos_current_bgr_2_0.D4.n15 pmos_current_bgr_2_0.D4.n14 2.7967
R11814 pmos_current_bgr_2_0.D4 pmos_current_bgr_2_0.D4.n0 2.61108
R11815 pmos_current_bgr_2_0.D4 pmos_current_bgr_2_0.D4.n2 2.46246
R11816 pmos_current_bgr_2_0.D4.n11 pmos_current_bgr_2_0.D4.n7 0.979361
R11817 pmos_current_bgr_2_0.D4.n17 pmos_current_bgr_2_0.D4.n16 0.979361
R11818 pmos_current_bgr_2_0.D4.n6 pmos_current_bgr_2_0.D4 0.951721
R11819 pmos_current_bgr_2_0.D4.n1 pmos_current_bgr_2_0.D4.n4 0.697467
R11820 pmos_current_bgr_2_0.D4.n0 pmos_current_bgr_2_0.D4.n5 0.697467
R11821 pmos_current_bgr_2_0.D4.n11 pmos_current_bgr_2_0.D4.n10 0.23963
R11822 pmos_current_bgr_2_0.D4.n17 pmos_current_bgr_2_0.D4.n15 0.23963
R11823 a_n4883_22159.t0 a_n4883_22159.t1 95.4796
R11824 a_n547_22325.t0 a_n547_22325.t1 95.4796
R11825 a_n17355_21661.t0 a_n17355_21661.t1 86.3178
R11826 a_n13555_21661.t0 a_n13555_21661.t1 95.4786
R11827 a_n13555_21329.t0 a_n13555_21329.t1 95.4796
R11828 a_n9219_21163.t0 a_n9219_21163.t1 95.4786
R11829 a_n13555_20997.t0 a_n13555_20997.t1 86.2637
R11830 a_n9219_20997.t0 a_n9219_20997.t1 86.2627
R11831 a_n9219_19433.t0 a_n9219_19433.t1 86.2637
R11832 a_n4883_19433.t0 a_n4883_19433.t1 86.2627
R11833 resistor_op_tt_0.A.n2 resistor_op_tt_0.A.t1 90.1607
R11834 resistor_op_tt_0.A.n1 resistor_op_tt_0.A.t2 87.6722
R11835 resistor_op_tt_0.A.n0 resistor_op_tt_0.A.t0 47.8785
R11836 resistor_op_tt_0.A resistor_op_tt_0.A.t3 47.6906
R11837 resistor_op_tt_0.A.n1 resistor_op_tt_0.A.n0 17.1313
R11838 resistor_op_tt_0.A.n2 resistor_op_tt_0.A.n1 1.7055
R11839 resistor_op_tt_0.A.n0 resistor_op_tt_0.A 0.279346
R11840 resistor_op_tt_0.A resistor_op_tt_0.A.n2 0.0189918
R11841 a_n4883_22325.t0 a_n4883_22325.t1 86.5527
R11842 a_n547_22159.t0 a_n547_22159.t1 86.5537
R11843 a_n17355_21495.t0 a_n17355_21495.t1 87.5628
R11844 a_n13555_21495.t0 a_n13555_21495.t1 86.5537
R11845 a_n9219_20595.t0 a_n9219_20595.t1 86.2627
R11846 a_n4883_20595.t0 a_n4883_20595.t1 86.2627
R11847 a_n4883_19931.t0 a_n4883_19931.t1 86.2637
R11848 a_n547_19931.t0 a_n547_19931.t1 86.2627
R11849 digital_0.S2.n10 digital_0.S2.t20 762.783
R11850 digital_0.S2.n10 digital_0.S2.t15 762.783
R11851 digital_0.S2.n6 digital_0.S2.t18 762.783
R11852 digital_0.S2.n6 digital_0.S2.t13 762.783
R11853 digital_0.S2.n11 digital_0.S2.n10 161.3
R11854 digital_0.S2.n7 digital_0.S2.n6 161.3
R11855 digital_0.S2.n20 digital_0.S2.t8 62.1591
R11856 digital_0.S2.n17 digital_0.S2.t30 50.9537
R11857 digital_0.S2.n0 digital_0.S2.t29 50.9537
R11858 digital_0.S2.n17 digital_0.S2.t26 50.711
R11859 digital_0.S2.n0 digital_0.S2.t3 50.711
R11860 digital_0.S2.n24 digital_0.S2.t0 48.6901
R11861 digital_0.S2.n22 digital_0.S2.t7 47.9666
R11862 digital_0.S2.n18 digital_0.S2.t9 47.7865
R11863 digital_0.S2.n18 digital_0.S2.t23 47.6925
R11864 digital_0.S2.n23 digital_0.S2.t28 47.6925
R11865 digital_0.S2.n24 digital_0.S2.t25 47.6059
R11866 digital_0.S2.n19 digital_0.S2.t31 47.5125
R11867 digital_0.S2.n22 digital_0.S2.t4 47.5125
R11868 digital_0.S2.n25 digital_0.S2.t24 47.4258
R11869 digital_0.S2.n7 digital_0.S2.t19 23.2859
R11870 digital_0.S2.n7 digital_0.S2.t14 23.2859
R11871 digital_0.S2.n11 digital_0.S2.t22 23.2669
R11872 digital_0.S2.n11 digital_0.S2.t17 23.2669
R11873 digital_0.S2.n8 digital_0.S2.n5 18.9359
R11874 digital_0.S2.n8 digital_0.S2.n4 18.9359
R11875 digital_0.S2.n9 digital_0.S2.n3 18.9169
R11876 digital_0.S2 digital_0.S2.n13 18.8194
R11877 digital_0.S2 digital_0.S2.n2 18.7973
R11878 digital_0.S2.n16 digital_0.S2.n15 18.0391
R11879 digital_0.S2.n29 digital_0.S2 11.46
R11880 digital_0.S2.n26 digital_0.S2.n25 6.43319
R11881 digital_0.S2.n25 digital_0.S2.n24 5.65435
R11882 digital_0.S2.n27 digital_0.S2.n21 5.45883
R11883 digital_0.S2.n15 digital_0.S2.t6 4.3505
R11884 digital_0.S2.n15 digital_0.S2.t5 4.3505
R11885 digital_0.S2.n13 digital_0.S2.t11 4.3505
R11886 digital_0.S2.n13 digital_0.S2.t27 4.3505
R11887 digital_0.S2.t14 digital_0.S2.n5 4.3505
R11888 digital_0.S2.n5 digital_0.S2.t12 4.3505
R11889 digital_0.S2.t19 digital_0.S2.n4 4.3505
R11890 digital_0.S2.n4 digital_0.S2.t10 4.3505
R11891 digital_0.S2.n3 digital_0.S2.t2 4.3505
R11892 digital_0.S2.n3 digital_0.S2.t16 4.3505
R11893 digital_0.S2.n2 digital_0.S2.t1 4.3505
R11894 digital_0.S2.n2 digital_0.S2.t21 4.3505
R11895 digital_0.S2.n14 digital_0.S2.n12 3.58944
R11896 digital_0.S2.n28 digital_0.S2.n17 3.19711
R11897 digital_0.S2.n1 digital_0.S2.n0 2.96069
R11898 digital_0.S2.n21 digital_0.S2.n20 2.72967
R11899 digital_0.S2.n27 digital_0.S2.n26 2.72967
R11900 digital_0.S2.n20 digital_0.S2.n19 1.27213
R11901 digital_0.S2.n9 digital_0.S2.n8 1.10293
R11902 digital_0.S2.n16 digital_0.S2.n14 0.941788
R11903 digital_0.S2 digital_0.S2.n1 0.911204
R11904 digital_0.S2.n26 digital_0.S2.n23 0.873096
R11905 digital_0.S2 digital_0.S2.n16 0.725879
R11906 digital_0.S2 digital_0.S2.n29 0.64704
R11907 digital_0.S2.n19 digital_0.S2.n18 0.274538
R11908 digital_0.S2.n23 digital_0.S2.n22 0.274538
R11909 digital_0.S2.n8 digital_0.S2.n7 0.190155
R11910 digital_0.S2.n21 digital_0.S2.n1 0.171
R11911 digital_0.S2.n28 digital_0.S2.n27 0.171
R11912 digital_0.S2.n14 digital_0.S2 0.161485
R11913 digital_0.S2.n9 digital_0.S2 0.120065
R11914 digital_0.S2.n12 digital_0.S2.n9 0.0768889
R11915 digital_0.S2.n12 digital_0.S2.n11 0.0768889
R11916 digital_0.S2.n29 digital_0.S2.n28 0.0382093
R11917 resistor_op_tt_0.D resistor_op_tt_0.D.t0 47.7647
R11918 resistor_op_tt_0.D.n2 resistor_op_tt_0.D.t3 47.5642
R11919 resistor_op_tt_0.D.n2 resistor_op_tt_0.D.n1 17.4377
R11920 resistor_op_tt_0.D resistor_op_tt_0.D.n2 0.853153
R11921 resistor_op_tt_0.D.n0 resistor_op_tt_0.D.t5 0.311679
R11922 resistor_op_tt_0.D.n1 resistor_op_tt_0.D.n0 0.180177
R11923 resistor_op_tt_0.D.t4 resistor_op_tt_0.D.t6 0.168944
R11924 resistor_op_tt_0.D.t7 resistor_op_tt_0.D.t4 0.118567
R11925 resistor_op_tt_0.D.t5 resistor_op_tt_0.D.t6 0.118
R11926 resistor_op_tt_0.D.n1 resistor_op_tt_0.D.t2 0.106544
R11927 resistor_op_tt_0.D.t5 resistor_op_tt_0.D 0.0974375
R11928 resistor_op_tt_0.D resistor_op_tt_0.D.t7 0.0720062
R11929 resistor_op_tt_0.D.n0 resistor_op_tt_0.D.t1 0.00317698
R11930 IPTAT.n0 IPTAT.t5 280.783
R11931 IPTAT.n0 IPTAT.t0 280.783
R11932 IPTAT.n6 IPTAT.t7 280.783
R11933 IPTAT.n6 IPTAT.t2 280.783
R11934 IPTAT.n7 IPTAT.t9 228.726
R11935 IPTAT.n7 IPTAT.t4 228.726
R11936 IPTAT.t6 IPTAT.n1 228.689
R11937 IPTAT.t1 IPTAT.n1 228.689
R11938 IPTAT.n9 IPTAT.n3 200.124
R11939 IPTAT.n9 IPTAT.n2 200.124
R11940 IPTAT.n8 IPTAT.n5 200.124
R11941 IPTAT.n8 IPTAT.n4 200.124
R11942 IPTAT.n1 IPTAT.n0 161.3
R11943 IPTAT.n7 IPTAT.n6 161.3
R11944 IPTAT.n3 IPTAT.t1 28.5655
R11945 IPTAT.n3 IPTAT.t12 28.5655
R11946 IPTAT.n2 IPTAT.t6 28.5655
R11947 IPTAT.n2 IPTAT.t10 28.5655
R11948 IPTAT.n5 IPTAT.t11 28.5655
R11949 IPTAT.n5 IPTAT.t3 28.5655
R11950 IPTAT.n4 IPTAT.t13 28.5655
R11951 IPTAT.n4 IPTAT.t8 28.5655
R11952 IPTAT.n7 IPTAT 17.5245
R11953 IPTAT.n9 IPTAT.n8 11.1853
R11954 IPTAT IPTAT.n1 0.234196
R11955 IPTAT.n8 IPTAT.n7 0.141804
R11956 IPTAT IPTAT.n9 0.00593478
R11957 DVDD.n9 DVDD.n5 13419.6
R11958 DVDD.n9 DVDD.n4 13419.6
R11959 DVDD.n16 DVDD.n4 11204
R11960 DVDD.n16 DVDD.n5 10991.4
R11961 DVDD.n15 DVDD.n6 6947.03
R11962 DVDD.n10 DVDD.n6 6947.03
R11963 DVDD.n10 DVDD.n7 6947.03
R11964 DVDD.n15 DVDD.n7 6947.03
R11965 DVDD.n19 DVDD.n2 4454.12
R11966 DVDD.n19 DVDD.n3 4454.12
R11967 DVDD.n21 DVDD.n2 4454.12
R11968 DVDD.n21 DVDD.n3 4454.12
R11969 DVDD.n14 DVDD.n8 1620.33
R11970 DVDD.n14 DVDD.n13 1620.33
R11971 DVDD.n11 DVDD.n8 1620.33
R11972 DVDD.n13 DVDD.n12 943.812
R11973 DVDD.n12 DVDD.n11 676.519
R11974 DVDD.n18 DVDD.n0 475.106
R11975 DVDD.n18 DVDD.n1 475.106
R11976 DVDD.n22 DVDD.n1 475.106
R11977 DVDD DVDD.n0 278.589
R11978 DVDD.t1 DVDD.n3 238.605
R11979 DVDD.t0 DVDD.n17 228.327
R11980 DVDD.n20 DVDD.t0 201.825
R11981 DVDD.n20 DVDD.t1 201.825
R11982 DVDD DVDD.n22 196.518
R11983 DVDD.n17 DVDD.n16 133.19
R11984 DVDD.n16 DVDD.n15 51.8889
R11985 DVDD.n12 DVDD 22.8033
R11986 DVDD.n22 DVDD.n21 10.8829
R11987 DVDD.n21 DVDD.n20 10.8829
R11988 DVDD.n19 DVDD.n18 10.8829
R11989 DVDD.n20 DVDD.n19 10.8829
R11990 DVDD.n3 DVDD.n1 10.2783
R11991 DVDD.n2 DVDD.n0 10.2783
R11992 DVDD.n17 DVDD.n2 10.2783
R11993 DVDD.n15 DVDD.n14 5.0005
R11994 DVDD.n11 DVDD.n10 5.0005
R11995 DVDD.n10 DVDD.n9 5.0005
R11996 DVDD.n8 DVDD.n6 2.10277
R11997 DVDD.n6 DVDD.n4 2.10277
R11998 DVDD.n13 DVDD.n7 2.10277
R11999 DVDD.n7 DVDD.n5 2.10277
R12000 a_3789_22325.t0 a_3789_22325.t1 86.5537
R12001 pmos_current_bgr_0.D1 pmos_current_bgr_0.D1.n1 202.694
R12002 pmos_current_bgr_0.D1.n2 pmos_current_bgr_0.D1.n0 201.903
R12003 pmos_current_bgr_0.D1.n3 pmos_current_bgr_0.D1.t0 42.5516
R12004 pmos_current_bgr_0.D1.n0 pmos_current_bgr_0.D1.t3 28.5655
R12005 pmos_current_bgr_0.D1.n0 pmos_current_bgr_0.D1.t1 28.5655
R12006 pmos_current_bgr_0.D1.n1 pmos_current_bgr_0.D1.t2 28.5655
R12007 pmos_current_bgr_0.D1.n1 pmos_current_bgr_0.D1.t4 28.5655
R12008 pmos_current_bgr_0.D1.n3 pmos_current_bgr_0.D1.n2 9.83481
R12009 pmos_current_bgr_0.D1 pmos_current_bgr_0.D1.n3 0.336214
R12010 pmos_current_bgr_0.D1.n2 pmos_current_bgr_0.D1 0.317979
R12011 a_n9219_21827.t0 a_n9219_21827.t1 86.5537
R12012 digital_0.SVBGSC.n1 digital_0.SVBGSC.n0 66.3172
R12013 digital_0.SVBGSC digital_0.SVBGSC.t1 54.9705
R12014 digital_0.SVBGSC.n2 digital_0.SVBGSC.n1 46.003
R12015 digital_0.SVBGSC.n2 digital_0.SVBGSC.t2 42.5516
R12016 digital_0.SVBGSC.n0 digital_0.SVBGSC.t3 17.4005
R12017 digital_0.SVBGSC.n0 digital_0.SVBGSC.t0 17.4005
R12018 digital_0.SVBGSC digital_0.SVBGSC.n2 3.13129
R12019 digital_0.SVBGSC.n1 digital_0.SVBGSC 0.224058
R12020 digital_0.SVBGSC.n1 digital_0.SVBGSC 0.221654
R12021 a_n4883_19765.t0 a_n4883_19765.t1 86.2637
R12022 a_n547_19765.t0 a_n547_19765.t1 86.2627
R12023 differential_pair_0.S.n2 differential_pair_0.S.t9 387.759
R12024 differential_pair_0.S.n7 differential_pair_0.S.t6 387.759
R12025 differential_pair_0.S.n5 differential_pair_0.S.n4 97.7157
R12026 differential_pair_0.S differential_pair_0.S.n3 97.4875
R12027 differential_pair_0.S.n1 differential_pair_0.S.t4 83.7522
R12028 differential_pair_0.S.n0 differential_pair_0.S.t5 83.7522
R12029 differential_pair_0.S.n1 differential_pair_0.S.t10 83.7172
R12030 differential_pair_0.S.n0 differential_pair_0.S.t8 83.7172
R12031 differential_pair_0.S.n7 differential_pair_0.S.t7 82.8128
R12032 differential_pair_0.S.n2 differential_pair_0.S.t11 82.8128
R12033 differential_pair_0.S.n3 differential_pair_0.S.t3 19.3338
R12034 differential_pair_0.S.n3 differential_pair_0.S.t0 19.3338
R12035 differential_pair_0.S.n4 differential_pair_0.S.t1 19.3338
R12036 differential_pair_0.S.n4 differential_pair_0.S.t2 19.3338
R12037 differential_pair_0.S.n5 differential_pair_0.S 17.4
R12038 differential_pair_0.S.n6 differential_pair_0.S 10.2251
R12039 differential_pair_0.S.n8 differential_pair_0.S.n6 8.59468
R12040 differential_pair_0.S.n6 differential_pair_0.S.n5 7.13003
R12041 differential_pair_0.S differential_pair_0.S.n8 6.6764
R12042 differential_pair_0.S differential_pair_0.S.n1 4.04356
R12043 differential_pair_0.S.n8 differential_pair_0.S.n0 3.9555
R12044 differential_pair_0.S.n1 differential_pair_0.S.n2 0.697467
R12045 differential_pair_0.S.n0 differential_pair_0.S.n7 0.697467
R12046 a_n4883_20429.t0 a_n4883_20429.t1 86.2637
R12047 a_n547_20429.t0 a_n547_20429.t1 86.2627
R12048 a_3789_22159.t0 a_3789_22159.t1 95.4786
R12049 a_8125_21993.t0 a_8125_21993.t1 95.6986
R12050 a_n4883_21329.t0 a_n4883_21329.t1 95.4786
R12051 a_3789_19931.t0 a_3789_19931.t1 86.2627
R12052 differential_pair_0.D4.n0 differential_pair_0.D4.t10 402.385
R12053 differential_pair_0.D4.n3 differential_pair_0.D4.t8 387.854
R12054 differential_pair_0.D4.n9 differential_pair_0.D4.t13 371.644
R12055 differential_pair_0.D4.n5 differential_pair_0.D4.t6 371.644
R12056 differential_pair_0.D4.n0 differential_pair_0.D4.t12 227.345
R12057 differential_pair_0.D4.t9 differential_pair_0.D4.n3 227.323
R12058 differential_pair_0.D4.n12 differential_pair_0.D4.n4 199.65
R12059 differential_pair_0.D4.n2 differential_pair_0.D4.n1 199.65
R12060 differential_pair_0.D4.t7 differential_pair_0.D4.n5 115.525
R12061 differential_pair_0.D4.n9 differential_pair_0.D4.t15 115.525
R12062 differential_pair_0.D4.n10 differential_pair_0.D4.n8 97.1505
R12063 differential_pair_0.D4.n7 differential_pair_0.D4.n6 97.1505
R12064 differential_pair_0.D4.n4 differential_pair_0.D4.t9 28.5655
R12065 differential_pair_0.D4.n4 differential_pair_0.D4.t3 28.5655
R12066 differential_pair_0.D4.n1 differential_pair_0.D4.t5 28.5655
R12067 differential_pair_0.D4.n1 differential_pair_0.D4.t11 28.5655
R12068 differential_pair_0.D4.n12 differential_pair_0.D4.n11 22.2572
R12069 differential_pair_0.D4.n8 differential_pair_0.D4.t0 19.3338
R12070 differential_pair_0.D4.n8 differential_pair_0.D4.t14 19.3338
R12071 differential_pair_0.D4.n6 differential_pair_0.D4.t7 19.3338
R12072 differential_pair_0.D4.n6 differential_pair_0.D4.t1 19.3338
R12073 differential_pair_0.D4.n13 differential_pair_0.D4.t16 11.5219
R12074 differential_pair_0.D4.n13 differential_pair_0.D4.t2 11.5219
R12075 differential_pair_0.D4.n14 differential_pair_0.D4.t4 11.5219
R12076 differential_pair_0.D4.n14 differential_pair_0.D4.t17 11.5219
R12077 differential_pair_0.D4.n11 differential_pair_0.D4 6.02466
R12078 differential_pair_0.D4 differential_pair_0.D4.n7 5.78569
R12079 differential_pair_0.D4.n11 differential_pair_0.D4.n10 3.9555
R12080 differential_pair_0.D4.n14 differential_pair_0.D4.n13 3.52397
R12081 differential_pair_0.D4.n13 differential_pair_0.D4.n12 2.60463
R12082 differential_pair_0.D4 differential_pair_0.D4.n14 1.81387
R12083 differential_pair_0.D4.n7 differential_pair_0.D4.n5 0.64517
R12084 differential_pair_0.D4.n10 differential_pair_0.D4.n9 0.64517
R12085 differential_pair_0.D4.n12 differential_pair_0.D4.n3 0.610341
R12086 differential_pair_0.D4.n2 differential_pair_0.D4.n0 0.586682
R12087 differential_pair_0.D4 differential_pair_0.D4.n2 0.346501
R12088 a_n4883_19599.t0 a_n4883_19599.t1 86.2637
R12089 a_n547_19599.t0 a_n547_19599.t1 86.2637
R12090 a_n4883_21661.t0 a_n4883_21661.t1 86.4732
R12091 a_n4883_22491.t0 a_n4883_22491.t1 86.2627
R12092 a_n547_22491.t0 a_n547_22491.t1 86.2637
R12093 a_8125_21827.t0 a_8125_21827.t1 86.7887
R12094 a_8125_19931.t0 a_8125_19931.t1 85.9587
R12095 VENA VENA.t1 118.347
R12096 VENA VENA.t0 118.347
R12097 VENA.n0 VENA.t2 118.005
R12098 VENA.n1 VENA.t3 118.005
R12099 VENA.n2 VENA 17.0005
R12100 VENA.n2 VENA.n1 1.13803
R12101 VENA VENA.n0 1.11546
R12102 VENA.n0 VENA 0.359196
R12103 VENA.n1 VENA 0.359196
R12104 VENA VENA.n2 0.0230694
R12105 VBGSC.n0 VBGSC.t3 387.61
R12106 VBGSC.n6 VBGSC.t0 380.147
R12107 VBGSC.n0 VBGSC.t4 83.1367
R12108 VBGSC.n5 VBGSC.t2 79.0672
R12109 VBGSC.n2 VBGSC.n1 66.7492
R12110 VBGSC.n8 VBGSC.n3 66.7492
R12111 VBGSC.n6 VBGSC.n5 58.3534
R12112 VBGSC.n1 VBGSC.t5 17.4005
R12113 VBGSC.n1 VBGSC.t6 17.4005
R12114 VBGSC.n3 VBGSC.t7 17.4005
R12115 VBGSC.n3 VBGSC.t1 17.4005
R12116 VBGSC.n4 VBGSC 13.2374
R12117 VBGSC.n7 VBGSC.n6 9.3005
R12118 VBGSC.n5 VBGSC.n4 4.6505
R12119 VBGSC VBGSC.n0 0.77179
R12120 VBGSC VBGSC.n2 0.652674
R12121 VBGSC VBGSC.n8 0.6255
R12122 VBGSC.n7 VBGSC.n4 0.390968
R12123 VBGSC.n8 VBGSC.n7 0.1255
R12124 VBGSC.n2 VBGSC 0.00321739
R12125 VBGTC.n0 VBGTC.t3 387.61
R12126 VBGTC.n6 VBGTC.t0 380.147
R12127 VBGTC.n0 VBGTC.t4 83.1367
R12128 VBGTC.n5 VBGTC.t2 79.0672
R12129 VBGTC.n2 VBGTC.n1 66.7492
R12130 VBGTC.n8 VBGTC.n3 66.7492
R12131 VBGTC.n6 VBGTC.n5 58.3534
R12132 VBGTC.n1 VBGTC.t5 17.4005
R12133 VBGTC.n1 VBGTC.t7 17.4005
R12134 VBGTC.n3 VBGTC.t6 17.4005
R12135 VBGTC.n3 VBGTC.t1 17.4005
R12136 VBGTC.n4 VBGTC 15.3456
R12137 VBGTC.n7 VBGTC.n6 9.3005
R12138 VBGTC.n5 VBGTC.n4 4.6505
R12139 VBGTC.n2 VBGTC.n0 0.774507
R12140 VBGTC VBGTC.n2 0.6255
R12141 VBGTC.n7 VBGTC.n4 0.390968
R12142 VBGTC.n8 VBGTC.n7 0.1255
R12143 VBGTC VBGTC.n8 0.0521304
R12144 a_3789_19765.t0 a_3789_19765.t1 86.2637
R12145 TRIM2.t1 TRIM2 190.643
R12146 TRIM2.t2 TRIM2.n1 190.585
R12147 TRIM2.n1 TRIM2.t3 190.585
R12148 TRIM2 TRIM2.t0 190.553
R12149 TRIM2.t3 TRIM2.n0 119.778
R12150 TRIM2.n0 TRIM2.t1 119.778
R12151 TRIM2.t0 TRIM2.n2 119.778
R12152 TRIM2.n2 TRIM2.t2 119.778
R12153 TRIM2.n2 TRIM2.n0 19.6878
R12154 TRIM2.n1 TRIM2 17.8418
R12155 differential_pair_0.PLUS.n1 differential_pair_0.PLUS.t3 67.3793
R12156 differential_pair_0.PLUS.n2 differential_pair_0.PLUS.t0 42.9618
R12157 differential_pair_0.PLUS.n0 differential_pair_0.PLUS.t1 42.894
R12158 differential_pair_0.PLUS.n1 differential_pair_0.PLUS.n0 14.0048
R12159 differential_pair_0.PLUS differential_pair_0.PLUS.t2 11.4392
R12160 differential_pair_0.PLUS.t3 differential_pair_0.PLUS 10.5356
R12161 differential_pair_0.PLUS.n2 differential_pair_0.PLUS.n1 8.02474
R12162 differential_pair_0.PLUS.n0 differential_pair_0.PLUS 0.0768889
R12163 differential_pair_0.PLUS differential_pair_0.PLUS.n2 0.0334861
R12164 a_n13555_21163.t0 a_n13555_21163.t1 86.5527
R12165 a_3789_20429.t0 a_3789_20429.t1 86.2637
R12166 a_n9219_20263.t0 a_n9219_20263.t1 86.2627
R12167 a_n4883_20263.t0 a_n4883_20263.t1 86.2627
R12168 a_8125_19599.t0 a_8125_19599.t1 85.9587
R12169 ENA.n1 ENA.n0 119.07
R12170 ENA.n2 ENA.t3 79.1268
R12171 ENA ENA.t1 78.5248
R12172 ENA.t0 ENA 78.4541
R12173 ENA.n2 ENA.t2 77.8672
R12174 ENA.n0 ENA.t0 24.1005
R12175 ENA.n1 ENA.t1 24.1005
R12176 ENA.t2 ENA.n1 24.1005
R12177 ENA.n0 ENA.t3 24.1005
R12178 ENA ENA.n2 0.157443
R12179 AVDD.n3 AVDD.n2 100.111
R12180 AVDD.n1 AVDD.n0 100.111
R12181 AVDD.n2 AVDD.t3 14.283
R12182 AVDD.n2 AVDD.t2 14.283
R12183 AVDD.n0 AVDD.t0 14.283
R12184 AVDD.n0 AVDD.t1 14.283
R12185 AVDD.n1 AVDD 4.42603
R12186 AVDD AVDD.n3 0.517787
R12187 AVDD AVDD.n1 0.273106
R12188 AVDD.n3 AVDD 0.254489
R12189 a_8125_20263.t0 a_8125_20263.t1 85.9587
R12190 TRIM1.t2 TRIM1 190.643
R12191 TRIM1.t1 TRIM1.n1 190.585
R12192 TRIM1.n1 TRIM1.t0 190.585
R12193 TRIM1 TRIM1.t3 190.544
R12194 TRIM1.t0 TRIM1.n0 119.778
R12195 TRIM1.n0 TRIM1.t2 119.778
R12196 TRIM1.t3 TRIM1.n2 119.778
R12197 TRIM1.n2 TRIM1.t1 119.778
R12198 TRIM1.n2 TRIM1.n0 19.6878
R12199 TRIM1.n1 TRIM1 15.5053
R12200 bjt_0.A.n3 bjt_0.A.n2 83.5719
R12201 bjt_0.A.t1 bjt_0.A.n0 65.0307
R12202 bjt_0.A.n2 bjt_0.A.n1 64.9507
R12203 bjt_0.A.n8 bjt_0.A.t0 42.5516
R12204 bjt_0.A.n7 bjt_0.A.t3 26.4846
R12205 bjt_0.A.n8 bjt_0.A.n7 20.3952
R12206 bjt_0.A.t3 bjt_0.A 12.9139
R12207 bjt_0.A bjt_0.A.t2 11.4791
R12208 bjt_0.A.n7 bjt_0.A 10.7496
R12209 bjt_0.A bjt_0.A.n6 4.79788
R12210 bjt_0.A.n3 bjt_0.A.n0 1.56328
R12211 bjt_0.A.n5 bjt_0.A.n4 1.5505
R12212 bjt_0.A.n5 bjt_0.A.n1 1.3347
R12213 bjt_0.A bjt_0.A.n1 1.27399
R12214 bjt_0.A.n4 bjt_0.A.n3 0.77514
R12215 bjt_0.A.n6 bjt_0.A.n0 0.533875
R12216 bjt_0.A bjt_0.A.n8 0.473
R12217 bjt_0.A.n4 bjt_0.A 0.314045
R12218 bjt_0.A.n2 bjt_0.A.t1 0.290206
R12219 bjt_0.A.n6 bjt_0.A.n5 0.00767213
R12220 a_3789_19599.t0 a_3789_19599.t1 86.2627
R12221 a_n547_21993.t0 a_n547_21993.t1 95.4796
R12222 a_3789_21827.t0 a_3789_21827.t1 95.4796
R12223 a_n13555_22159.t0 a_n13555_22159.t1 95.4796
R12224 a_n9219_22325.t0 a_n9219_22325.t1 95.4786
R12225 a_3789_22491.t0 a_3789_22491.t1 86.2637
R12226 a_n9219_20097.t0 a_n9219_20097.t1 86.2637
R12227 a_n4883_20097.t0 a_n4883_20097.t1 86.2637
R12228 a_n547_19433.t0 a_n547_19433.t1 86.2637
R12229 digital_0.SVBGTC.n1 digital_0.SVBGTC.n0 66.3172
R12230 digital_0.SVBGTC digital_0.SVBGTC.t2 43.4301
R12231 digital_0.SVBGTC.n2 digital_0.SVBGTC.t3 42.5516
R12232 digital_0.SVBGTC.n2 digital_0.SVBGTC.n1 40.9088
R12233 digital_0.SVBGTC.n0 digital_0.SVBGTC.t1 17.4005
R12234 digital_0.SVBGTC.n0 digital_0.SVBGTC.t0 17.4005
R12235 digital_0.SVBGTC digital_0.SVBGTC.n2 0.573
R12236 digital_0.SVBGTC.n1 digital_0.SVBGTC 0.221654
R12237 digital_0.SVBGTC.n1 digital_0.SVBGTC 0.221654
R12238 a_n547_20595.t0 a_n547_20595.t1 86.2637
R12239 a_n13555_22325.t0 a_n13555_22325.t1 86.5537
R12240 a_n9219_22159.t0 a_n9219_22159.t1 86.5527
R12241 a_n9219_21661.t0 a_n9219_21661.t1 86.5527
R12242 a_n4883_21495.n0 a_n4883_21495.t1 43.3791
R12243 a_n4883_21495.n1 a_n4883_21495.t3 43.3541
R12244 a_n4883_21495.t0 a_n4883_21495.n1 43.2001
R12245 a_n4883_21495.n0 a_n4883_21495.t2 43.1741
R12246 a_n4883_21495.n1 a_n4883_21495.n0 10.9342
R12247 a_n13019_19765.t0 a_n13019_19765.t1 86.3178
R12248 a_n9219_19931.t0 a_n9219_19931.t1 86.2627
R12249 a_n9219_21993.n1 a_n9219_21993.t3 47.7671
R12250 a_n9219_21993.n0 a_n9219_21993.t1 47.7671
R12251 a_n9219_21993.t0 a_n9219_21993.n1 47.588
R12252 a_n9219_21993.n0 a_n9219_21993.t2 47.587
R12253 a_n9219_21993.n1 a_n9219_21993.n0 10.4236
R12254 a_3789_19433.t0 a_3789_19433.t1 86.2637
R12255 a_n9219_19765.t0 a_n9219_19765.t1 86.2627
R12256 a_n9219_20429.t0 a_n9219_20429.t1 86.2627
R12257 a_n4883_21163.t0 a_n4883_21163.t1 86.5527
R12258 a_n547_21329.t0 a_n547_21329.t1 86.5537
R12259 a_3789_20595.t0 a_3789_20595.t1 86.2627
R12260 pmos_startup_0.D2.n1 pmos_startup_0.D2.t2 396.214
R12261 pmos_startup_0.D2.n0 pmos_startup_0.D2.t4 223.565
R12262 pmos_startup_0.D2.n4 pmos_startup_0.D2.n3 199.65
R12263 pmos_startup_0.D2.n1 pmos_startup_0.D2.n0 62.1181
R12264 pmos_startup_0.D2.n5 pmos_startup_0.D2.t1 42.5516
R12265 pmos_startup_0.D2.n3 pmos_startup_0.D2.t0 28.5655
R12266 pmos_startup_0.D2.n3 pmos_startup_0.D2.t3 28.5655
R12267 pmos_startup_0.D2.n5 pmos_startup_0.D2.n4 25.2687
R12268 pmos_startup_0.D2 pmos_startup_0.D2.t5 20.1605
R12269 pmos_startup_0.D2.n2 pmos_startup_0.D2.n1 9.89749
R12270 pmos_startup_0.D2.n4 pmos_startup_0.D2.n0 4.6505
R12271 pmos_startup_0.D2.n2 pmos_startup_0.D2 0.559447
R12272 pmos_startup_0.D2 pmos_startup_0.D2.n5 0.490885
R12273 pmos_startup_0.D2.n4 pmos_startup_0.D2.n2 0.0802101
R12274 a_n9219_19599.t0 a_n9219_19599.t1 86.2627
R12275 a_n13555_21993.t0 a_n13555_21993.t1 86.5527
R12276 a_n13555_22491.t0 a_n13555_22491.t1 86.2637
R12277 a_n9219_22491.t0 a_n9219_22491.t1 86.2627
R12278 a_n547_20263.t0 a_n547_20263.t1 86.2637
R12279 a_n547_21163.t0 a_n547_21163.t1 95.4796
R12280 a_3789_21329.t0 a_3789_21329.t1 95.4796
R12281 a_n9219_21329.t0 a_n9219_21329.t1 86.5537
R12282 a_n4883_20997.t0 a_n4883_20997.t1 86.2637
R12283 a_220_15663.t0 a_220_15663.t1 86.2627
R12284 a_3789_21163.t0 a_3789_21163.t1 86.5527
R12285 a_8125_21329.t0 a_8125_21329.t1 86.7887
R12286 a_n547_20097.t0 a_n547_20097.t1 86.2627
R12287 a_220_14999.n0 a_220_14999.t3 43.3316
R12288 a_220_14999.n1 a_220_14999.t1 43.3316
R12289 a_220_14999.n0 a_220_14999.t2 43.2216
R12290 a_220_14999.t0 a_220_14999.n1 43.2216
R12291 a_220_14999.n1 a_220_14999.n0 0.2905
R12292 a_3789_20263.t0 a_3789_20263.t1 86.2627
R12293 a_n9219_21495.t0 a_n9219_21495.t1 105.778
R12294 a_n547_21495.t0 a_n547_21495.t1 95.4796
R12295 a_3789_21661.t0 a_3789_21661.t1 95.4796
R12296 a_3789_20097.t0 a_3789_20097.t1 86.2637
R12297 a_n13555_21827.t0 a_n13555_21827.t1 95.4786
R12298 a_3789_21495.t0 a_3789_21495.t1 86.5527
R12299 a_220_15165.n0 a_220_15165.t3 47.9666
R12300 a_220_15165.t0 a_220_15165.n1 47.8948
R12301 a_220_15165.n0 a_220_15165.t2 47.5125
R12302 a_220_15165.n1 a_220_15165.t1 47.5125
R12303 a_220_15165.n1 a_220_15165.n0 0.274538
R12304 a_8125_21163.t0 a_8125_21163.t1 95.6986
R12305 a_n547_20997.t0 a_n547_20997.t1 86.2627
R12306 a_n13019_20097.t0 a_n13019_20097.t1 86.3178
R12307 a_3789_20997.t0 a_3789_20997.t1 86.2627
R12308 a_220_14833.t0 a_220_14833.t1 86.2637
C0 TRIM0 VBGSC 0.290536f
C1 bjt_0.A pmos_iptat_0.G 1.34154f
C2 digital_0.D3 resistor_op_tt_0.C 0.642112f
C3 bjt_0.A pmos_current_bgr_2_0.D4 0.439226f
C4 digital_0.S1 digital_0.D3 1.09705f
C5 AVSS digital_0.S2 5.6467f
C6 bjt_0.B digital_0.SVBGTC 0.013521f
C7 pmos_startup_0.D4 digital_0.S3 0.407034f
C8 DVSS AVDD 0.026303f
C9 differential_pair_0.D4 digital_0.S2 0.103746f
C10 digital_0.S1 TRIM0 0.821992f
C11 DVDD ENA 2.01375f
C12 digital_0.S3 pmos_iptat_0.G 0.38912f
C13 TRIM3 digital_0.S3 0.837131f
C14 digital_0.S3 pmos_current_bgr_2_0.D4 0.242603f
C15 AVSS digital_0.D3 5.07156f
C16 VENA digital_0.SVBGSC 0.225908f
C17 TRIM0 VBGTC 0.02382f
C18 bjt_0.A resistor_op_tt_0.A 0.224331f
C19 resistor_op_tt_0.D digital_0.S2 0.035226f
C20 differential_pair_0.D4 digital_0.D3 0.235409f
C21 IPTAT pmos_iptat_0.G 2.63111f
C22 digital_0.S1 digital_0.SVBGTC 0.015728f
C23 AVSS TRIM0 0.074767f
C24 VBGTC digital_0.SVBGTC 0.217701f
C25 DVDD VENA 0.176292f
C26 digital_0.S2 differential_pair_0.PLUS 3.35649f
C27 pmos_startup_0.D3 digital_0.S2 0.131403f
C28 AVSS digital_0.SVBGTC 1.15405f
C29 bjt_0.B resistor_op_tt_0.C 0.124784f
C30 digital_0.S1 bjt_0.B 10.653299f
C31 bjt_0.A differential_pair_0.S 2.16604f
C32 digital_0.S2 pmos_current_bgr_2_0.D3 1.17414f
C33 DVSS TRIM2 1.20602f
C34 digital_0.D3 differential_pair_0.PLUS 0.355881f
C35 pmos_startup_0.D3 digital_0.D3 0.029044f
C36 differential_pair_0.D4 digital_0.SVBGTC 0.014097f
C37 digital_0.S1 VBGSC 0.120116f
C38 DVDD TRIM3 5.47702f
C39 bjt_0.A VREF 0.200895f
C40 TRIM0 ENA 0.187761f
C41 VBGTC VBGSC 0.039872f
C42 digital_0.D3 pmos_current_bgr_2_0.D3 0.840252f
C43 bjt_0.B AVSS 24.3328f
C44 pmos_current_bgr_0.D1 resistor_op_tt_0.C 0.030922f
C45 pmos_startup_0.D4 digital_0.S2 0.195841f
C46 AVSS VBGSC 0.054158f
C47 bjt_0.B differential_pair_0.D4 0.073365f
C48 digital_0.S1 resistor_op_tt_0.C 0.091103f
C49 digital_0.S2 pmos_iptat_0.G 0.154947f
C50 TRIM3 digital_0.S2 0.027722f
C51 digital_0.S1 VBGTC 0.120525f
C52 DVDD AVDD 0.172656f
C53 digital_0.S2 pmos_current_bgr_2_0.D4 0.860291f
C54 TRIM2 digital_0.S3 0.810324f
C55 bjt_0.B resistor_op_tt_0.D 0.346223f
C56 digital_0.SVBGTC differential_pair_0.PLUS 0.010625f
C57 pmos_startup_0.D4 digital_0.D3 0.025699f
C58 pmos_current_bgr_0.D1 AVSS 2.13024f
C59 TRIM0 VENA 0.0528f
C60 AVSS resistor_op_tt_0.C 3.06824f
C61 digital_0.S1 AVSS 15.9884f
C62 digital_0.D3 pmos_iptat_0.G 0.02808f
C63 TRIM3 digital_0.D3 0.853722f
C64 pmos_startup_0.D2 pmos_current_bgr_0.D1 0.120526f
C65 digital_0.D3 pmos_current_bgr_2_0.D4 0.163561f
C66 pmos_startup_0.D2 resistor_op_tt_0.C 0.065453f
C67 pmos_startup_0.D2 digital_0.S1 1.58128f
C68 DVSS digital_0.S3 1.791f
C69 differential_pair_0.D4 resistor_op_tt_0.C 3.37647f
C70 AVSS VBGTC 0.050682f
C71 digital_0.S1 differential_pair_0.D4 0.051294f
C72 bjt_0.B differential_pair_0.PLUS 0.261906f
C73 resistor_op_tt_0.A digital_0.S2 0.026511f
C74 bjt_0.B pmos_startup_0.D3 0.176319f
C75 VBGSC ENA 0.010892f
C76 VENA digital_0.SVBGTC 0.165958f
C77 TRIM2 TRIM1 3.6069f
C78 resistor_op_tt_0.D resistor_op_tt_0.C 0.154415f
C79 digital_0.S1 resistor_op_tt_0.D 0.065113f
C80 bjt_0.A digital_0.S3 0.995483f
C81 bjt_0.B pmos_current_bgr_2_0.D3 0.121734f
C82 resistor_op_tt_0.A digital_0.D3 0.041388f
C83 pmos_startup_0.D2 AVSS 2.75508f
C84 AVSS differential_pair_0.D4 2.68929f
C85 DVSS digital_0.SVBGSC 0.219171f
C86 DVSS TRIM1 1.22775f
C87 pmos_current_bgr_0.D1 differential_pair_0.PLUS 0.486932f
C88 bjt_0.B VENA 0.013339f
C89 digital_0.SVBGTC pmos_current_bgr_2_0.D4 0.024673f
C90 DVDD TRIM2 0.705102f
C91 resistor_op_tt_0.C differential_pair_0.PLUS 1.54711f
C92 AVSS resistor_op_tt_0.D 36.806396f
C93 digital_0.S1 differential_pair_0.PLUS 0.149112f
C94 pmos_startup_0.D3 resistor_op_tt_0.C 0.271361f
C95 digital_0.S1 pmos_startup_0.D3 0.141437f
C96 VENA VBGSC 2.53218f
C97 VBGTC ENA 0.277091f
C98 differential_pair_0.S digital_0.S2 0.424583f
C99 bjt_0.B pmos_startup_0.D4 0.531297f
C100 resistor_op_tt_0.C pmos_current_bgr_2_0.D3 0.936647f
C101 digital_0.S1 pmos_current_bgr_2_0.D3 0.333707f
C102 DVDD DVSS 37.036f
C103 AVSS ENA 0.140855f
C104 bjt_0.B pmos_iptat_0.G 0.604849f
C105 bjt_0.B TRIM3 0.07834f
C106 bjt_0.B pmos_current_bgr_2_0.D4 0.085388f
C107 AVSS differential_pair_0.PLUS 10.5874f
C108 differential_pair_0.S digital_0.D3 0.284266f
C109 AVSS pmos_startup_0.D3 2.70865f
C110 TRIM2 digital_0.S2 0.843265f
C111 TRIM3 VBGSC 0.024016f
C112 digital_0.S1 VENA 0.036749f
C113 digital_0.SVBGSC digital_0.S3 0.168167f
C114 pmos_startup_0.D2 differential_pair_0.PLUS 0.143558f
C115 differential_pair_0.D4 differential_pair_0.PLUS 1.85403f
C116 pmos_startup_0.D2 pmos_startup_0.D3 2.20668f
C117 differential_pair_0.D4 pmos_startup_0.D3 0.085711f
C118 VBGTC VENA 2.9551f
C119 AVSS pmos_current_bgr_2_0.D3 28.122301f
C120 pmos_startup_0.D4 resistor_op_tt_0.C 0.053416f
C121 digital_0.S1 pmos_startup_0.D4 0.143357f
C122 pmos_current_bgr_0.D1 pmos_iptat_0.G 0.732931f
C123 pmos_startup_0.D2 pmos_current_bgr_2_0.D3 0.015501f
C124 differential_pair_0.D4 pmos_current_bgr_2_0.D3 2.57724f
C125 DVSS digital_0.S2 1.81813f
C126 pmos_iptat_0.G resistor_op_tt_0.C 15.1435f
C127 AVSS VENA 0.01642f
C128 digital_0.S1 pmos_iptat_0.G 0.410505f
C129 resistor_op_tt_0.C pmos_current_bgr_2_0.D4 1.34052f
C130 digital_0.S1 pmos_current_bgr_2_0.D4 0.10491f
C131 DVDD digital_0.S3 0.131466f
C132 DVSS digital_0.D3 1.73276f
C133 differential_pair_0.S digital_0.SVBGTC 0.022169f
C134 bjt_0.A digital_0.S2 0.292711f
C135 AVSS pmos_startup_0.D4 2.11275f
C136 pmos_startup_0.D3 differential_pair_0.PLUS 0.12938f
C137 pmos_startup_0.D2 pmos_startup_0.D4 0.110797f
C138 differential_pair_0.D4 pmos_startup_0.D4 0.050767f
C139 AVSS pmos_iptat_0.G 13.536f
C140 AVSS TRIM3 0.022971f
C141 AVSS pmos_current_bgr_2_0.D4 2.90704f
C142 resistor_op_tt_0.A resistor_op_tt_0.C 1.10585f
C143 DVSS TRIM0 1.45712f
C144 bjt_0.A digital_0.D3 0.232573f
C145 pmos_startup_0.D2 pmos_iptat_0.G 1.03404f
C146 differential_pair_0.D4 pmos_iptat_0.G 0.78978f
C147 pmos_current_bgr_2_0.D3 differential_pair_0.PLUS 1.55462f
C148 digital_0.S3 digital_0.S2 4.72495f
C149 DVDD digital_0.SVBGSC 0.081846f
C150 DVDD TRIM1 0.358436f
C151 differential_pair_0.D4 pmos_current_bgr_2_0.D4 3.30024f
C152 pmos_startup_0.D3 pmos_current_bgr_2_0.D3 0.31894f
C153 VENA ENA 0.163316f
C154 VBGTC AVDD 0.331838f
C155 resistor_op_tt_0.D pmos_iptat_0.G 0.111254p
C156 digital_0.D3 digital_0.S3 6.44683f
C157 DVSS digital_0.SVBGTC 0.128562f
C158 AVSS resistor_op_tt_0.A 3.77888f
C159 AVSS AVDD 0.115133f
C160 bjt_0.B TRIM2 0.05547f
C161 pmos_startup_0.D4 differential_pair_0.PLUS 0.034396f
C162 pmos_startup_0.D3 pmos_startup_0.D4 0.77828f
C163 differential_pair_0.D4 resistor_op_tt_0.A 0.192913f
C164 TRIM1 digital_0.S2 0.814485f
C165 digital_0.SVBGSC digital_0.S2 0.023826f
C166 TRIM2 VBGSC 0.036964f
C167 differential_pair_0.S resistor_op_tt_0.C 0.994325f
C168 pmos_iptat_0.G differential_pair_0.PLUS 0.361875f
C169 pmos_startup_0.D3 pmos_iptat_0.G 0.621429f
C170 pmos_current_bgr_2_0.D4 differential_pair_0.PLUS 1.19339f
C171 pmos_current_bgr_0.D1 VREF 1.45117f
C172 pmos_startup_0.D3 pmos_current_bgr_2_0.D4 0.368843f
C173 pmos_startup_0.D4 pmos_current_bgr_2_0.D3 0.543903f
C174 bjt_0.B DVSS 0.19911f
C175 VREF resistor_op_tt_0.C 1.18857f
C176 digital_0.SVBGSC digital_0.D3 1.29194f
C177 pmos_iptat_0.G pmos_current_bgr_2_0.D3 2.39226f
C178 DVSS VBGSC 0.785843f
C179 pmos_current_bgr_2_0.D3 pmos_current_bgr_2_0.D4 5.13521f
C180 digital_0.S1 TRIM2 0.02805f
C181 DVDD digital_0.S2 0.120279f
C182 digital_0.SVBGTC digital_0.S3 0.106412f
C183 AVSS differential_pair_0.S 9.56994f
C184 bjt_0.A bjt_0.B 5.69045f
C185 ENA AVDD 0.756313f
C186 TRIM1 TRIM0 3.1119f
C187 TRIM0 digital_0.SVBGSC 0.044673f
C188 resistor_op_tt_0.A differential_pair_0.PLUS 0.178161f
C189 differential_pair_0.D4 differential_pair_0.S 0.578071f
C190 AVSS VREF 3.73112f
C191 DVDD digital_0.D3 0.242278f
C192 digital_0.S1 DVSS 1.89744f
C193 pmos_startup_0.D4 pmos_iptat_0.G 0.274708f
C194 AVSS TRIM2 0.021887f
C195 resistor_op_tt_0.A pmos_current_bgr_2_0.D3 0.700007f
C196 pmos_startup_0.D4 pmos_current_bgr_2_0.D4 0.488571f
C197 bjt_0.B digital_0.S3 1.15682f
C198 DVSS VBGTC 0.727026f
C199 pmos_current_bgr_0.D1 bjt_0.A 3.26218f
C200 digital_0.SVBGSC digital_0.SVBGTC 6.82108f
C201 DVDD TRIM0 0.297131f
C202 pmos_iptat_0.G pmos_current_bgr_2_0.D4 2.8934f
C203 bjt_0.A resistor_op_tt_0.C 3.03083f
C204 bjt_0.A digital_0.S1 0.647837f
C205 AVSS DVSS 0.119249f
C206 digital_0.D3 digital_0.S2 2.04794f
C207 differential_pair_0.S differential_pair_0.PLUS 2.00341f
C208 bjt_0.B digital_0.SVBGSC 0.125306f
C209 bjt_0.B TRIM1 0.057977f
C210 DVDD digital_0.SVBGTC 0.097878f
C211 digital_0.S3 resistor_op_tt_0.C 0.107236f
C212 digital_0.S1 digital_0.S3 5.41062f
C213 VREF differential_pair_0.PLUS 0.156823f
C214 bjt_0.A AVSS 14.061999f
C215 TRIM1 VBGSC 0.06357f
C216 differential_pair_0.S pmos_current_bgr_2_0.D3 3.0408f
C217 resistor_op_tt_0.A pmos_current_bgr_2_0.D4 0.124876f
C218 VBGSC digital_0.SVBGSC 0.316962f
C219 pmos_startup_0.D2 bjt_0.A 0.767931f
C220 bjt_0.A differential_pair_0.D4 1.99159f
C221 digital_0.S1 IPTAT 0.022613f
C222 bjt_0.B DVDD 0.201231f
C223 AVSS digital_0.S3 6.79901f
C224 bjt_0.A resistor_op_tt_0.D 1.98499f
C225 DVSS ENA 0.136427f
C226 digital_0.SVBGTC digital_0.S2 0.027737f
C227 digital_0.S1 digital_0.SVBGSC 0.128462f
C228 digital_0.S1 TRIM1 0.847144f
C229 pmos_startup_0.D2 digital_0.S3 0.037495f
C230 DVDD VBGSC 0.081251f
C231 differential_pair_0.D4 digital_0.S3 0.190837f
C232 VBGTC digital_0.SVBGSC 0.280586f
C233 differential_pair_0.S pmos_iptat_0.G 1.29567f
C234 AVSS IPTAT 0.920267f
C235 digital_0.SVBGTC digital_0.D3 7.03954f
C236 differential_pair_0.S pmos_current_bgr_2_0.D4 0.861683f
C237 resistor_op_tt_0.D digital_0.S3 0.586743f
C238 bjt_0.A differential_pair_0.PLUS 7.484169f
C239 bjt_0.A pmos_startup_0.D3 0.332112f
C240 VREF pmos_iptat_0.G 4.73595f
C241 bjt_0.B digital_0.S2 6.41383f
C242 AVSS TRIM1 0.021887f
C243 AVSS digital_0.SVBGSC 3.07141f
C244 digital_0.S1 DVDD 0.121251f
C245 DVSS VENA 1.46332f
C246 TRIM3 TRIM2 4.10673f
C247 differential_pair_0.D4 digital_0.SVBGSC 0.010335f
C248 bjt_0.A pmos_current_bgr_2_0.D3 0.251504f
C249 DVDD VBGTC 0.229944f
C250 bjt_0.B digital_0.D3 0.536248f
C251 digital_0.S3 differential_pair_0.PLUS 0.229111f
C252 pmos_startup_0.D3 digital_0.S3 0.892384f
C253 resistor_op_tt_0.A differential_pair_0.S 0.112712f
C254 AVSS DVDD 0.119514f
C255 DVSS TRIM3 1.22291f
C256 digital_0.S2 resistor_op_tt_0.C 0.094543f
C257 digital_0.S3 pmos_current_bgr_2_0.D3 0.076657f
C258 digital_0.S1 digital_0.S2 10.2985f
C259 bjt_0.B TRIM0 0.606702f
C260 bjt_0.A pmos_startup_0.D4 0.117727f
C261 AVDD VSUBS 0.942396f
C262 ENA VSUBS 2.350606f
C263 VBGSC VSUBS 1.661369f
C264 VENA VSUBS 2.859062f
C265 VBGTC VSUBS 1.583076f
C266 TRIM0 VSUBS 1.718918f
C267 TRIM1 VSUBS 2.258568f
C268 TRIM2 VSUBS 2.564478f
C269 TRIM3 VSUBS 3.139189f
C270 IPTAT VSUBS 1.855772f
C271 VREF VSUBS 5.035279f
C272 DVSS VSUBS 6.536457f
C273 AVSS VSUBS 0.214153p
C274 DVDD VSUBS 58.821274f
C275 resistor_op_tt_0.D VSUBS 4.501713f
C276 differential_pair_0.S VSUBS 6.828552f
C277 resistor_op_tt_0.A VSUBS 1.337532f
C278 pmos_startup_0.D4 VSUBS 1.751466f
C279 pmos_startup_0.D3 VSUBS 2.997227f
C280 differential_pair_0.D4 VSUBS 7.794115f
C281 pmos_current_bgr_2_0.D4 VSUBS 7.847576f
C282 pmos_current_bgr_2_0.D3 VSUBS 20.231037f
C283 resistor_op_tt_0.C VSUBS 10.004482f
C284 pmos_iptat_0.G VSUBS 21.0945f
C285 digital_0.S2 VSUBS 8.264129f
C286 digital_0.S3 VSUBS 10.147709f
C287 bjt_0.B VSUBS 4.604816f
C288 digital_0.S1 VSUBS 14.705749f
C289 pmos_startup_0.D2 VSUBS 3.059782f
C290 bjt_0.A VSUBS 12.409239f
C291 differential_pair_0.PLUS VSUBS 8.8754f
C292 digital_0.D3 VSUBS 8.76654f
C293 digital_0.SVBGTC VSUBS 1.966834f
C294 digital_0.SVBGSC VSUBS 4.814141f
C295 pmos_current_bgr_0.D1 VSUBS 1.781014f
C296 pmos_startup_0.D2.t4 VSUBS 0.067616f
C297 pmos_startup_0.D2.n0 VSUBS 0.048045f
C298 pmos_startup_0.D2.t5 VSUBS 3.65855f
C299 pmos_startup_0.D2.t2 VSUBS 0.049302f
C300 pmos_startup_0.D2.n1 VSUBS 0.056657f
C301 pmos_startup_0.D2.n2 VSUBS 0.075243f
C302 pmos_startup_0.D2.t0 VSUBS 0.018695f
C303 pmos_startup_0.D2.t3 VSUBS 0.018695f
C304 pmos_startup_0.D2.n3 VSUBS 0.038453f
C305 pmos_startup_0.D2.n4 VSUBS 1.85272f
C306 pmos_startup_0.D2.t1 VSUBS 0.066332f
C307 pmos_startup_0.D2.n5 VSUBS 2.63737f
C308 digital_0.SVBGTC.t1 VSUBS 0.030862f
C309 digital_0.SVBGTC.t0 VSUBS 0.030862f
C310 digital_0.SVBGTC.n0 VSUBS 0.067002f
C311 digital_0.SVBGTC.n1 VSUBS 6.155879f
C312 digital_0.SVBGTC.t3 VSUBS 0.109501f
C313 digital_0.SVBGTC.n2 VSUBS 6.28177f
C314 digital_0.SVBGTC.t2 VSUBS 0.127956f
C315 bjt_0.A.n0 VSUBS 0.955382f
C316 bjt_0.A.n1 VSUBS 0.780733f
C317 bjt_0.A.t1 VSUBS 0.529178f
C318 bjt_0.A.n2 VSUBS 0.524137f
C319 bjt_0.A.n3 VSUBS 0.241693f
C320 bjt_0.A.n4 VSUBS 0.093529f
C321 bjt_0.A.n5 VSUBS 1.28489f
C322 bjt_0.A.n6 VSUBS 2.2661f
C323 bjt_0.A.t2 VSUBS 2.80784f
C324 bjt_0.A.t3 VSUBS 5.16071f
C325 bjt_0.A.n7 VSUBS 12.019099f
C326 bjt_0.A.t0 VSUBS 0.047006f
C327 bjt_0.A.n8 VSUBS 5.4969f
C328 TRIM1.t2 VSUBS 0.655731f
C329 TRIM1.n0 VSUBS 0.577587f
C330 TRIM1.t0 VSUBS 0.655654f
C331 TRIM1.n1 VSUBS 1.46016f
C332 TRIM1.t1 VSUBS 0.655654f
C333 TRIM1.n2 VSUBS 0.577587f
C334 TRIM1.t3 VSUBS 0.6556f
C335 ENA.t3 VSUBS 0.223539f
C336 ENA.t1 VSUBS 0.222894f
C337 ENA.t0 VSUBS 0.222826f
C338 ENA.n0 VSUBS 0.275486f
C339 ENA.n1 VSUBS 0.275486f
C340 ENA.t2 VSUBS 0.222325f
C341 ENA.n2 VSUBS 0.145498f
C342 differential_pair_0.PLUS.t0 VSUBS 0.059649f
C343 differential_pair_0.PLUS.t1 VSUBS 0.059071f
C344 differential_pair_0.PLUS.n0 VSUBS 1.22709f
C345 differential_pair_0.PLUS.t2 VSUBS 3.51175f
C346 differential_pair_0.PLUS.t3 VSUBS 8.2646f
C347 differential_pair_0.PLUS.n1 VSUBS 7.63385f
C348 differential_pair_0.PLUS.n2 VSUBS 0.408578f
C349 TRIM2.t1 VSUBS 0.723162f
C350 TRIM2.n0 VSUBS 0.636982f
C351 TRIM2.t3 VSUBS 0.723077f
C352 TRIM2.n1 VSUBS 1.76576f
C353 TRIM2.t2 VSUBS 0.723077f
C354 TRIM2.n2 VSUBS 0.636982f
C355 TRIM2.t0 VSUBS 0.723029f
C356 VBGTC.t3 VSUBS 0.048432f
C357 VBGTC.t4 VSUBS 0.063393f
C358 VBGTC.n0 VSUBS 0.115649f
C359 VBGTC.t5 VSUBS 0.018176f
C360 VBGTC.t7 VSUBS 0.018176f
C361 VBGTC.n1 VSUBS 0.040061f
C362 VBGTC.n2 VSUBS 0.231711f
C363 VBGTC.t6 VSUBS 0.018176f
C364 VBGTC.t1 VSUBS 0.018176f
C365 VBGTC.n3 VSUBS 0.040061f
C366 VBGTC.n4 VSUBS 0.876991f
C367 VBGTC.t2 VSUBS 0.060703f
C368 VBGTC.n5 VSUBS 0.050677f
C369 VBGTC.t0 VSUBS 0.04745f
C370 VBGTC.n6 VSUBS 0.051007f
C371 VBGTC.n7 VSUBS 0.036021f
C372 VBGTC.n8 VSUBS 0.131913f
C373 VBGSC.t3 VSUBS 0.0449f
C374 VBGSC.t4 VSUBS 0.058769f
C375 VBGSC.n0 VSUBS 0.106906f
C376 VBGSC.t5 VSUBS 0.01685f
C377 VBGSC.t6 VSUBS 0.01685f
C378 VBGSC.n1 VSUBS 0.03714f
C379 VBGSC.n2 VSUBS 0.145233f
C380 VBGSC.t7 VSUBS 0.01685f
C381 VBGSC.t1 VSUBS 0.01685f
C382 VBGSC.n3 VSUBS 0.03714f
C383 VBGSC.n4 VSUBS 0.670698f
C384 VBGSC.t2 VSUBS 0.056277f
C385 VBGSC.n5 VSUBS 0.046981f
C386 VBGSC.t0 VSUBS 0.043989f
C387 VBGSC.n6 VSUBS 0.047287f
C388 VBGSC.n7 VSUBS 0.033394f
C389 VBGSC.n8 VSUBS 0.150492f
C390 VENA.t1 VSUBS 0.430752f
C391 VENA.t2 VSUBS 0.430184f
C392 VENA.n0 VSUBS 0.244955f
C393 VENA.t0 VSUBS 0.430752f
C394 VENA.t3 VSUBS 0.430184f
C395 VENA.n1 VSUBS 0.246908f
C396 VENA.n2 VSUBS 1.06089f
C397 differential_pair_0.D4.t12 VSUBS 0.052514f
C398 differential_pair_0.D4.t10 VSUBS 0.038632f
C399 differential_pair_0.D4.n0 VSUBS 0.078162f
C400 differential_pair_0.D4.t5 VSUBS 0.014351f
C401 differential_pair_0.D4.t11 VSUBS 0.014351f
C402 differential_pair_0.D4.n1 VSUBS 0.029516f
C403 differential_pair_0.D4.n2 VSUBS 0.185981f
C404 differential_pair_0.D4.t8 VSUBS 0.038012f
C405 differential_pair_0.D4.n3 VSUBS 0.079026f
C406 differential_pair_0.D4.t9 VSUBS 0.066861f
C407 differential_pair_0.D4.t3 VSUBS 0.014351f
C408 differential_pair_0.D4.n4 VSUBS 0.029516f
C409 differential_pair_0.D4.t6 VSUBS 0.036422f
C410 differential_pair_0.D4.n5 VSUBS 0.071725f
C411 differential_pair_0.D4.t7 VSUBS 0.058989f
C412 differential_pair_0.D4.t1 VSUBS 0.012916f
C413 differential_pair_0.D4.n6 VSUBS 0.027345f
C414 differential_pair_0.D4.n7 VSUBS 0.229832f
C415 differential_pair_0.D4.t0 VSUBS 0.012916f
C416 differential_pair_0.D4.t14 VSUBS 0.012916f
C417 differential_pair_0.D4.n8 VSUBS 0.027345f
C418 differential_pair_0.D4.t13 VSUBS 0.036422f
C419 differential_pair_0.D4.t15 VSUBS 0.046073f
C420 differential_pair_0.D4.n9 VSUBS 0.071725f
C421 differential_pair_0.D4.n10 VSUBS 0.200583f
C422 differential_pair_0.D4.n11 VSUBS 1.66219f
C423 differential_pair_0.D4.n12 VSUBS 1.25694f
C424 differential_pair_0.D4.t2 VSUBS 2.53126f
C425 differential_pair_0.D4.t16 VSUBS 2.53126f
C426 differential_pair_0.D4.n13 VSUBS 1.43075f
C427 differential_pair_0.D4.t17 VSUBS 2.53126f
C428 differential_pair_0.D4.t4 VSUBS 2.53126f
C429 differential_pair_0.D4.n14 VSUBS 1.38674f
C430 differential_pair_0.S.n0 VSUBS 0.811557f
C431 differential_pair_0.S.n1 VSUBS 0.816014f
C432 differential_pair_0.S.t4 VSUBS 0.112861f
C433 differential_pair_0.S.t9 VSUBS 0.085609f
C434 differential_pair_0.S.t11 VSUBS 0.111297f
C435 differential_pair_0.S.n2 VSUBS 0.190122f
C436 differential_pair_0.S.t10 VSUBS 0.112775f
C437 differential_pair_0.S.t3 VSUBS 0.028901f
C438 differential_pair_0.S.t0 VSUBS 0.028901f
C439 differential_pair_0.S.n3 VSUBS 0.06169f
C440 differential_pair_0.S.t1 VSUBS 0.028901f
C441 differential_pair_0.S.t2 VSUBS 0.028901f
C442 differential_pair_0.S.n4 VSUBS 0.062151f
C443 differential_pair_0.S.n5 VSUBS 2.52893f
C444 differential_pair_0.S.n6 VSUBS 1.7146f
C445 differential_pair_0.S.t7 VSUBS 0.111297f
C446 differential_pair_0.S.t6 VSUBS 0.085609f
C447 differential_pair_0.S.n7 VSUBS 0.190122f
C448 differential_pair_0.S.t8 VSUBS 0.112775f
C449 differential_pair_0.S.t5 VSUBS 0.112861f
C450 differential_pair_0.S.n8 VSUBS 3.58518f
C451 digital_0.SVBGSC.t3 VSUBS 0.0155f
C452 digital_0.SVBGSC.t0 VSUBS 0.0155f
C453 digital_0.SVBGSC.n0 VSUBS 0.033649f
C454 digital_0.SVBGSC.n1 VSUBS 4.09448f
C455 digital_0.SVBGSC.t2 VSUBS 0.054993f
C456 digital_0.SVBGSC.n2 VSUBS 4.3479f
C457 digital_0.SVBGSC.t1 VSUBS 0.229152f
C458 pmos_current_bgr_0.D1.t3 VSUBS 0.014351f
C459 pmos_current_bgr_0.D1.t1 VSUBS 0.014351f
C460 pmos_current_bgr_0.D1.n0 VSUBS 0.030537f
C461 pmos_current_bgr_0.D1.t2 VSUBS 0.014351f
C462 pmos_current_bgr_0.D1.t4 VSUBS 0.014351f
C463 pmos_current_bgr_0.D1.n1 VSUBS 0.031154f
C464 pmos_current_bgr_0.D1.n2 VSUBS 2.20783f
C465 pmos_current_bgr_0.D1.t0 VSUBS 0.050917f
C466 pmos_current_bgr_0.D1.n3 VSUBS 2.75825f
C467 DVDD.n0 VSUBS 0.163652f
C468 DVDD.n1 VSUBS 0.206823f
C469 DVDD.n2 VSUBS 0.206823f
C470 DVDD.n3 VSUBS 1.61289f
C471 DVDD.n4 VSUBS 5.11721f
C472 DVDD.n5 VSUBS 5.07038f
C473 DVDD.n6 VSUBS 1.51531f
C474 DVDD.n7 VSUBS 1.51531f
C475 DVDD.n8 VSUBS 0.697583f
C476 DVDD.n9 VSUBS 5.78024f
C477 DVDD.n10 VSUBS 1.52611f
C478 DVDD.n11 VSUBS 0.496f
C479 DVDD.n12 VSUBS 1.24171f
C480 DVDD.n13 VSUBS 0.551482f
C481 DVDD.n14 VSUBS 0.699826f
C482 DVDD.n15 VSUBS 2.17798f
C483 DVDD.n16 VSUBS 5.83962f
C484 DVDD.n17 VSUBS 1.76856f
C485 DVDD.t0 VSUBS 2.10432f
C486 DVDD.t1 VSUBS 2.16761f
C487 DVDD.n18 VSUBS 0.206805f
C488 DVDD.n19 VSUBS 0.206805f
C489 DVDD.n20 VSUBS 1.97467f
C490 DVDD.n21 VSUBS 0.206805f
C491 DVDD.n22 VSUBS 0.145606f
C492 IPTAT.t5 VSUBS 0.034151f
C493 IPTAT.t0 VSUBS 0.034151f
C494 IPTAT.n0 VSUBS 0.073722f
C495 IPTAT.n1 VSUBS 0.321222f
C496 IPTAT.t6 VSUBS 0.094234f
C497 IPTAT.t10 VSUBS 0.02011f
C498 IPTAT.n2 VSUBS 0.041615f
C499 IPTAT.t1 VSUBS 0.094234f
C500 IPTAT.t12 VSUBS 0.02011f
C501 IPTAT.n3 VSUBS 0.041615f
C502 IPTAT.t13 VSUBS 0.02011f
C503 IPTAT.t8 VSUBS 0.02011f
C504 IPTAT.n4 VSUBS 0.041615f
C505 IPTAT.t11 VSUBS 0.02011f
C506 IPTAT.t3 VSUBS 0.02011f
C507 IPTAT.n5 VSUBS 0.041615f
C508 IPTAT.t9 VSUBS 0.074148f
C509 IPTAT.t7 VSUBS 0.034151f
C510 IPTAT.t2 VSUBS 0.034151f
C511 IPTAT.n6 VSUBS 0.073722f
C512 IPTAT.t4 VSUBS 0.074148f
C513 IPTAT.n7 VSUBS 1.06005f
C514 IPTAT.n8 VSUBS 0.934835f
C515 IPTAT.n9 VSUBS 0.926861f
C516 resistor_op_tt_0.D.t0 VSUBS 0.030522f
C517 resistor_op_tt_0.D.t3 VSUBS 0.029973f
C518 resistor_op_tt_0.D.t6 VSUBS 21.8311f
C519 resistor_op_tt_0.D.t4 VSUBS 21.488901f
C520 resistor_op_tt_0.D.t7 VSUBS 19.5616f
C521 resistor_op_tt_0.D.t5 VSUBS 20.4635f
C522 resistor_op_tt_0.D.t1 VSUBS 19.5345f
C523 resistor_op_tt_0.D.n0 VSUBS 18.0907f
C524 resistor_op_tt_0.D.t2 VSUBS 20.6365f
C525 resistor_op_tt_0.D.n1 VSUBS 2.03835f
C526 resistor_op_tt_0.D.n2 VSUBS 0.898923f
C527 digital_0.S2.t3 VSUBS 0.139354f
C528 digital_0.S2.t29 VSUBS 0.139844f
C529 digital_0.S2.n0 VSUBS 1.93562f
C530 digital_0.S2.n1 VSUBS 1.428f
C531 digital_0.S2.t1 VSUBS 0.072743f
C532 digital_0.S2.t21 VSUBS 0.072743f
C533 digital_0.S2.n2 VSUBS 0.174202f
C534 digital_0.S2.t2 VSUBS 0.072743f
C535 digital_0.S2.t16 VSUBS 0.072743f
C536 digital_0.S2.n3 VSUBS 0.176639f
C537 digital_0.S2.t10 VSUBS 0.072743f
C538 digital_0.S2.n4 VSUBS 0.177031f
C539 digital_0.S2.t12 VSUBS 0.072743f
C540 digital_0.S2.n5 VSUBS 0.177031f
C541 digital_0.S2.t14 VSUBS 0.348599f
C542 digital_0.S2.t19 VSUBS 0.348599f
C543 digital_0.S2.t18 VSUBS 0.115211f
C544 digital_0.S2.t13 VSUBS 0.115211f
C545 digital_0.S2.n6 VSUBS 0.12377f
C546 digital_0.S2.n7 VSUBS 0.913184f
C547 digital_0.S2.n8 VSUBS 0.891327f
C548 digital_0.S2.n9 VSUBS 0.502374f
C549 digital_0.S2.t17 VSUBS 0.275499f
C550 digital_0.S2.t22 VSUBS 0.275499f
C551 digital_0.S2.t20 VSUBS 0.115211f
C552 digital_0.S2.t15 VSUBS 0.115211f
C553 digital_0.S2.n10 VSUBS 0.12377f
C554 digital_0.S2.n11 VSUBS 0.905809f
C555 digital_0.S2.n12 VSUBS 0.062385f
C556 digital_0.S2.t11 VSUBS 0.072743f
C557 digital_0.S2.t27 VSUBS 0.072743f
C558 digital_0.S2.n13 VSUBS 0.19519f
C559 digital_0.S2.n14 VSUBS 0.282705f
C560 digital_0.S2.t6 VSUBS 0.072743f
C561 digital_0.S2.t5 VSUBS 0.072743f
C562 digital_0.S2.n15 VSUBS 0.164282f
C563 digital_0.S2.n16 VSUBS 0.679035f
C564 digital_0.S2.t26 VSUBS 0.139354f
C565 digital_0.S2.t30 VSUBS 0.139844f
C566 digital_0.S2.n17 VSUBS 2.00243f
C567 digital_0.S2.t9 VSUBS 0.115209f
C568 digital_0.S2.t23 VSUBS 0.112436f
C569 digital_0.S2.n18 VSUBS 0.952998f
C570 digital_0.S2.t31 VSUBS 0.112523f
C571 digital_0.S2.n19 VSUBS 0.554756f
C572 digital_0.S2.t8 VSUBS 0.454339f
C573 digital_0.S2.n20 VSUBS 2.41089f
C574 digital_0.S2.n21 VSUBS 0.774779f
C575 digital_0.S2.t7 VSUBS 0.115113f
C576 digital_0.S2.t4 VSUBS 0.112523f
C577 digital_0.S2.n22 VSUBS 0.953008f
C578 digital_0.S2.t28 VSUBS 0.112436f
C579 digital_0.S2.n23 VSUBS 0.527777f
C580 digital_0.S2.t24 VSUBS 0.111754f
C581 digital_0.S2.t25 VSUBS 0.11167f
C582 digital_0.S2.t0 VSUBS 0.123067f
C583 digital_0.S2.n24 VSUBS 1.42686f
C584 digital_0.S2.n25 VSUBS 1.27991f
C585 digital_0.S2.n26 VSUBS 0.71669f
C586 digital_0.S2.n27 VSUBS 0.774779f
C587 digital_0.S2.n28 VSUBS 1.11676f
C588 digital_0.S2.n29 VSUBS 2.51325f
C589 resistor_op_tt_0.A.t1 VSUBS 0.082092f
C590 resistor_op_tt_0.A.t3 VSUBS 0.112911f
C591 resistor_op_tt_0.A.t0 VSUBS 0.114861f
C592 resistor_op_tt_0.A.n0 VSUBS 1.16243f
C593 resistor_op_tt_0.A.t2 VSUBS 0.070753f
C594 resistor_op_tt_0.A.n1 VSUBS 0.79981f
C595 resistor_op_tt_0.A.n2 VSUBS 0.922604f
C596 pmos_current_bgr_2_0.D4.n0 VSUBS 0.406151f
C597 pmos_current_bgr_2_0.D4.n1 VSUBS 2.68175f
C598 pmos_current_bgr_2_0.D4.t17 VSUBS 2.97636f
C599 pmos_current_bgr_2_0.D4.n2 VSUBS 0.586081f
C600 pmos_current_bgr_2_0.D4.t5 VSUBS 0.016874f
C601 pmos_current_bgr_2_0.D4.t15 VSUBS 0.016874f
C602 pmos_current_bgr_2_0.D4.n3 VSUBS 0.034871f
C603 pmos_current_bgr_2_0.D4.t12 VSUBS 0.058484f
C604 pmos_current_bgr_2_0.D4.t11 VSUBS 0.044985f
C605 pmos_current_bgr_2_0.D4.n4 VSUBS 0.099905f
C606 pmos_current_bgr_2_0.D4.t13 VSUBS 0.059261f
C607 pmos_current_bgr_2_0.D4.t0 VSUBS 0.059306f
C608 pmos_current_bgr_2_0.D4.t1 VSUBS 0.059306f
C609 pmos_current_bgr_2_0.D4.t8 VSUBS 0.058484f
C610 pmos_current_bgr_2_0.D4.t6 VSUBS 0.044985f
C611 pmos_current_bgr_2_0.D4.n5 VSUBS 0.099905f
C612 pmos_current_bgr_2_0.D4.t7 VSUBS 0.059261f
C613 pmos_current_bgr_2_0.D4.n6 VSUBS 2.32398f
C614 pmos_current_bgr_2_0.D4.t9 VSUBS 0.04545f
C615 pmos_current_bgr_2_0.D4.n7 VSUBS 0.119398f
C616 pmos_current_bgr_2_0.D4.t10 VSUBS 0.07862f
C617 pmos_current_bgr_2_0.D4.t3 VSUBS 0.016874f
C618 pmos_current_bgr_2_0.D4.n8 VSUBS 0.034871f
C619 pmos_current_bgr_2_0.D4.t2 VSUBS 2.97636f
C620 pmos_current_bgr_2_0.D4.n9 VSUBS 0.602542f
C621 pmos_current_bgr_2_0.D4.n10 VSUBS 0.25402f
C622 pmos_current_bgr_2_0.D4.n11 VSUBS 0.205232f
C623 pmos_current_bgr_2_0.D4.n12 VSUBS 0.766987f
C624 pmos_current_bgr_2_0.D4.t18 VSUBS 2.97636f
C625 pmos_current_bgr_2_0.D4.n13 VSUBS 0.800822f
C626 pmos_current_bgr_2_0.D4.t4 VSUBS 2.97636f
C627 pmos_current_bgr_2_0.D4.n14 VSUBS 0.602542f
C628 pmos_current_bgr_2_0.D4.n15 VSUBS 0.25402f
C629 pmos_current_bgr_2_0.D4.t14 VSUBS 0.04545f
C630 pmos_current_bgr_2_0.D4.t16 VSUBS 0.061746f
C631 pmos_current_bgr_2_0.D4.n16 VSUBS 0.119398f
C632 pmos_current_bgr_2_0.D4.n17 VSUBS 0.271091f
C633 pmos_startup_0.D3.n0 VSUBS 0.657088f
C634 pmos_startup_0.D3.n1 VSUBS 0.080309f
C635 pmos_startup_0.D3.t18 VSUBS 2.79024f
C636 pmos_startup_0.D3.t12 VSUBS 2.61787f
C637 pmos_startup_0.D3.n2 VSUBS 0.882869f
C638 pmos_startup_0.D3.t13 VSUBS 0.014842f
C639 pmos_startup_0.D3.n3 VSUBS 0.030526f
C640 pmos_startup_0.D3.t6 VSUBS 0.069153f
C641 pmos_startup_0.D3.t5 VSUBS 0.039937f
C642 pmos_startup_0.D3.t9 VSUBS 0.039584f
C643 pmos_startup_0.D3.t11 VSUBS 0.051438f
C644 pmos_startup_0.D3.n4 VSUBS 0.08106f
C645 pmos_startup_0.D3.t15 VSUBS 0.014842f
C646 pmos_startup_0.D3.t10 VSUBS 0.014842f
C647 pmos_startup_0.D3.n5 VSUBS 0.032221f
C648 pmos_startup_0.D3.n6 VSUBS 0.178779f
C649 pmos_startup_0.D3.t14 VSUBS 0.014842f
C650 pmos_startup_0.D3.t3 VSUBS 0.014842f
C651 pmos_startup_0.D3.n7 VSUBS 0.032221f
C652 pmos_startup_0.D3.t4 VSUBS 0.051438f
C653 pmos_startup_0.D3.t2 VSUBS 0.039584f
C654 pmos_startup_0.D3.n8 VSUBS 0.08106f
C655 pmos_startup_0.D3.n9 VSUBS 0.178779f
C656 pmos_startup_0.D3.n10 VSUBS 0.054961f
C657 pmos_startup_0.D3.n11 VSUBS 1.12008f
C658 pmos_startup_0.D3.t7 VSUBS 0.039584f
C659 pmos_startup_0.D3.n12 VSUBS 0.08106f
C660 pmos_startup_0.D3.t8 VSUBS 0.066279f
C661 pmos_startup_0.D3.t17 VSUBS 0.014842f
C662 pmos_startup_0.D3.n13 VSUBS 0.032221f
C663 pmos_startup_0.D3.n14 VSUBS 0.178779f
C664 pmos_startup_0.D3.t16 VSUBS 0.014842f
C665 pmos_startup_0.D3.n15 VSUBS 0.032221f
C666 pmos_startup_0.D3.t1 VSUBS 0.066279f
C667 pmos_startup_0.D3.t0 VSUBS 0.039584f
C668 pmos_startup_0.D3.n16 VSUBS 0.08106f
C669 pmos_startup_0.D3.n17 VSUBS 0.178779f
C670 pmos_startup_0.D3.n18 VSUBS 0.054961f
C671 pmos_startup_0.D4.t3 VSUBS 0.173651f
C672 pmos_startup_0.D4.t4 VSUBS 0.173651f
C673 pmos_startup_0.D4.n0 VSUBS 0.111122f
C674 pmos_startup_0.D4.t5 VSUBS 0.173651f
C675 pmos_startup_0.D4.n1 VSUBS 0.107723f
C676 pmos_startup_0.D4.t6 VSUBS 0.231747f
C677 pmos_startup_0.D4.t0 VSUBS 0.024668f
C678 pmos_startup_0.D4.t1 VSUBS 0.042715f
C679 pmos_startup_0.D4.n2 VSUBS 0.018863f
C680 pmos_iptat_0.G.t22 VSUBS 79.8206f
C681 pmos_iptat_0.G.n0 VSUBS 0.120646f
C682 pmos_iptat_0.G.n1 VSUBS 0.483523f
C683 pmos_iptat_0.G.t29 VSUBS 2.64901f
C684 pmos_iptat_0.G.t13 VSUBS 0.017687f
C685 pmos_iptat_0.G.t12 VSUBS 0.013605f
C686 pmos_iptat_0.G.n2 VSUBS 0.030214f
C687 pmos_iptat_0.G.t14 VSUBS 0.017922f
C688 pmos_iptat_0.G.t0 VSUBS 0.017936f
C689 pmos_iptat_0.G.t1 VSUBS 0.017936f
C690 pmos_iptat_0.G.t8 VSUBS 0.017687f
C691 pmos_iptat_0.G.t6 VSUBS 0.013605f
C692 pmos_iptat_0.G.n3 VSUBS 0.030214f
C693 pmos_iptat_0.G.t7 VSUBS 0.017922f
C694 pmos_iptat_0.G.n4 VSUBS 0.165509f
C695 pmos_iptat_0.G.t27 VSUBS 81.5995f
C696 pmos_iptat_0.G.n5 VSUBS 1.37275f
C697 pmos_iptat_0.G.n6 VSUBS 0.133475f
C698 pmos_iptat_0.G.n7 VSUBS 0.366162f
C699 pmos_iptat_0.G.t11 VSUBS 0.018673f
C700 pmos_iptat_0.G.t9 VSUBS 0.013757f
C701 pmos_iptat_0.G.n8 VSUBS 0.028136f
C702 pmos_iptat_0.G.n9 VSUBS 0.010496f
C703 pmos_iptat_0.G.n10 VSUBS 0.064575f
C704 pmos_iptat_0.G.n11 VSUBS 0.403991f
C705 pmos_iptat_0.G.n12 VSUBS 0.222639f
C706 pmos_iptat_0.G.t23 VSUBS 2.90644f
C707 pmos_iptat_0.G.n13 VSUBS 0.366162f
C708 pmos_iptat_0.G.t4 VSUBS 0.013757f
C709 pmos_iptat_0.G.n14 VSUBS 0.028136f
C710 pmos_iptat_0.G.t5 VSUBS 0.023777f
C711 pmos_iptat_0.G.n15 VSUBS 0.010496f
C712 pmos_iptat_0.G.n16 VSUBS 0.064575f
C713 pmos_iptat_0.G.n17 VSUBS 0.085627f
C714 pmos_iptat_0.G.n18 VSUBS 0.242783f
C715 pmos_iptat_0.G.t2 VSUBS 0.013758f
C716 pmos_iptat_0.G.n19 VSUBS 0.028162f
C717 pmos_iptat_0.G.t3 VSUBS 0.023776f
C718 pmos_iptat_0.G.n20 VSUBS 0.010496f
C719 pmos_iptat_0.G.n21 VSUBS 0.064548f
C720 pmos_iptat_0.G.n22 VSUBS 0.403555f
C721 pmos_iptat_0.G.n23 VSUBS 0.366162f
C722 pmos_iptat_0.G.n24 VSUBS 0.222639f
C723 pmos_iptat_0.G.n25 VSUBS 0.222639f
C724 pmos_iptat_0.G.n26 VSUBS 0.222639f
C725 pmos_iptat_0.G.t26 VSUBS 2.90644f
C726 pmos_iptat_0.G.t24 VSUBS 3.55039f
C727 pmos_iptat_0.G.t25 VSUBS 3.55042f
C728 pmos_iptat_0.G.n27 VSUBS 0.366162f
C729 pmos_iptat_0.G.n28 VSUBS 0.242783f
C730 pmos_iptat_0.G.n29 VSUBS 0.242783f
C731 pmos_iptat_0.G.n30 VSUBS 0.010496f
C732 pmos_iptat_0.G.t15 VSUBS 0.013757f
C733 pmos_iptat_0.G.t17 VSUBS 0.018673f
C734 pmos_iptat_0.G.n31 VSUBS 0.028136f
C735 pmos_iptat_0.G.n32 VSUBS 0.064575f
C736 pmos_iptat_0.G.n33 VSUBS 0.277144f
C737 pmos_iptat_0.G.n34 VSUBS 0.324639f
C738 pmos_iptat_0.G.t28 VSUBS 2.67077f
C739 pmos_iptat_0.G.n35 VSUBS 0.332746f
C740 pmos_iptat_0.G.n36 VSUBS 0.634339f
C741 pmos_iptat_0.G.n37 VSUBS 0.200394f
C742 resistor_op_tt_0.C.t4 VSUBS 0.081337f
C743 resistor_op_tt_0.C.n0 VSUBS 0.568296f
C744 resistor_op_tt_0.C.t7 VSUBS 0.08405f
C745 resistor_op_tt_0.C.t5 VSUBS 0.061921f
C746 resistor_op_tt_0.C.n1 VSUBS 0.126645f
C747 resistor_op_tt_0.C.t3 VSUBS 0.02297f
C748 resistor_op_tt_0.C.t6 VSUBS 0.02297f
C749 resistor_op_tt_0.C.n2 VSUBS 0.047245f
C750 resistor_op_tt_0.C.n3 VSUBS 0.290657f
C751 resistor_op_tt_0.C.t16 VSUBS 4.05164f
C752 resistor_op_tt_0.C.n4 VSUBS 1.76879f
C753 resistor_op_tt_0.C.t18 VSUBS 4.05164f
C754 resistor_op_tt_0.C.n5 VSUBS 2.62749f
C755 resistor_op_tt_0.C.t17 VSUBS 4.05164f
C756 resistor_op_tt_0.C.n6 VSUBS 2.62749f
C757 resistor_op_tt_0.C.t19 VSUBS 4.05164f
C758 resistor_op_tt_0.C.n7 VSUBS 2.24311f
C759 resistor_op_tt_0.C.n8 VSUBS 0.493046f
C760 resistor_op_tt_0.C.n9 VSUBS 0.239302f
C761 resistor_op_tt_0.C.t8 VSUBS 0.061921f
C762 resistor_op_tt_0.C.n10 VSUBS 0.126645f
C763 resistor_op_tt_0.C.t9 VSUBS 0.10702f
C764 resistor_op_tt_0.C.t15 VSUBS 0.02297f
C765 resistor_op_tt_0.C.n11 VSUBS 0.047245f
C766 resistor_op_tt_0.C.n12 VSUBS 0.290657f
C767 resistor_op_tt_0.C.n13 VSUBS 2.38587f
C768 resistor_op_tt_0.C.t13 VSUBS 0.058299f
C769 resistor_op_tt_0.C.n14 VSUBS 0.114806f
C770 resistor_op_tt_0.C.t14 VSUBS 0.09442f
C771 resistor_op_tt_0.C.t2 VSUBS 0.020673f
C772 resistor_op_tt_0.C.n15 VSUBS 0.04377f
C773 resistor_op_tt_0.C.n16 VSUBS 0.32471f
C774 resistor_op_tt_0.C.t12 VSUBS 0.073747f
C775 resistor_op_tt_0.C.t10 VSUBS 0.058299f
C776 resistor_op_tt_0.C.n17 VSUBS 0.114806f
C777 resistor_op_tt_0.C.t1 VSUBS 0.020673f
C778 resistor_op_tt_0.C.t11 VSUBS 0.020673f
C779 resistor_op_tt_0.C.n18 VSUBS 0.04377f
C780 resistor_op_tt_0.C.n19 VSUBS 0.287406f
C781 resistor_op_tt_0.C.n20 VSUBS 1.35946f
C782 resistor_op_tt_0.C.n21 VSUBS 2.03246f
C783 resistor_op_tt_0.C.n22 VSUBS 0.321353f
C784 resistor_op_tt_0.C.t0 VSUBS 0.081339f
C785 resistor_op_tt_0.C.n23 VSUBS 0.519479f
C786 digital_0.D3.t15 VSUBS 0.050267f
C787 digital_0.D3.n0 VSUBS 2.14775f
C788 digital_0.D3.t16 VSUBS 0.093021f
C789 digital_0.D3.n1 VSUBS 2.58248f
C790 digital_0.D3.t10 VSUBS 0.056784f
C791 digital_0.D3.t3 VSUBS 0.056784f
C792 digital_0.D3.n2 VSUBS 0.120004f
C793 digital_0.D3.t12 VSUBS 0.056784f
C794 digital_0.D3.t8 VSUBS 0.056784f
C795 digital_0.D3.n3 VSUBS 0.138191f
C796 digital_0.D3.t11 VSUBS 0.056784f
C797 digital_0.D3.n4 VSUBS 0.138191f
C798 digital_0.D3.t13 VSUBS 0.056784f
C799 digital_0.D3.n5 VSUBS 0.138191f
C800 digital_0.D3.t6 VSUBS 0.272118f
C801 digital_0.D3.t1 VSUBS 0.272118f
C802 digital_0.D3.t0 VSUBS 0.089934f
C803 digital_0.D3.t5 VSUBS 0.089934f
C804 digital_0.D3.n6 VSUBS 0.096615f
C805 digital_0.D3.n7 VSUBS 0.712835f
C806 digital_0.D3.n8 VSUBS 0.696357f
C807 digital_0.D3.t9 VSUBS 0.215335f
C808 digital_0.D3.t4 VSUBS 0.215335f
C809 digital_0.D3.t2 VSUBS 0.089934f
C810 digital_0.D3.t7 VSUBS 0.089934f
C811 digital_0.D3.n9 VSUBS 0.096615f
C812 digital_0.D3.n10 VSUBS 0.712835f
C813 digital_0.D3.n11 VSUBS 0.396792f
C814 digital_0.D3.n12 VSUBS 2.30238f
C815 digital_0.D3.n13 VSUBS 3.85849f
C816 digital_0.D3.t14 VSUBS 0.273644f
C817 digital_0.S3.t8 VSUBS 0.143066f
C818 digital_0.S3.n0 VSUBS 1.83866f
C819 digital_0.S3.t7 VSUBS 0.085393f
C820 digital_0.S3.t5 VSUBS 0.051338f
C821 digital_0.S3.t18 VSUBS 0.051338f
C822 digital_0.S3.n1 VSUBS 0.122943f
C823 digital_0.S3.t11 VSUBS 0.051338f
C824 digital_0.S3.t13 VSUBS 0.051338f
C825 digital_0.S3.n2 VSUBS 0.124663f
C826 digital_0.S3.t6 VSUBS 0.051338f
C827 digital_0.S3.n3 VSUBS 0.12494f
C828 digital_0.S3.t9 VSUBS 0.051338f
C829 digital_0.S3.n4 VSUBS 0.12494f
C830 digital_0.S3.t21 VSUBS 0.246023f
C831 digital_0.S3.t16 VSUBS 0.246023f
C832 digital_0.S3.t15 VSUBS 0.08131f
C833 digital_0.S3.t20 VSUBS 0.08131f
C834 digital_0.S3.n5 VSUBS 0.087351f
C835 digital_0.S3.n6 VSUBS 0.644478f
C836 digital_0.S3.n7 VSUBS 0.629053f
C837 digital_0.S3.n8 VSUBS 0.354549f
C838 digital_0.S3.t14 VSUBS 0.194433f
C839 digital_0.S3.t19 VSUBS 0.194433f
C840 digital_0.S3.t17 VSUBS 0.08131f
C841 digital_0.S3.t12 VSUBS 0.08131f
C842 digital_0.S3.n9 VSUBS 0.087351f
C843 digital_0.S3.n10 VSUBS 0.639273f
C844 digital_0.S3.n11 VSUBS 0.044028f
C845 digital_0.S3.t3 VSUBS 0.051338f
C846 digital_0.S3.t2 VSUBS 0.051338f
C847 digital_0.S3.n12 VSUBS 0.137798f
C848 digital_0.S3.n13 VSUBS 0.199519f
C849 digital_0.S3.t0 VSUBS 0.051338f
C850 digital_0.S3.t1 VSUBS 0.051338f
C851 digital_0.S3.n14 VSUBS 0.115941f
C852 digital_0.S3.n15 VSUBS 0.478936f
C853 digital_0.S3.n16 VSUBS 4.23617f
C854 digital_0.S3.t22 VSUBS 0.191674f
C855 digital_0.S3.t4 VSUBS 0.103553f
C856 digital_0.S3.n17 VSUBS 2.82847f
C857 digital_0.S3.n18 VSUBS 0.701352f
C858 digital_0.S3.t10 VSUBS 0.186677f
C859 digital_0.S3.t23 VSUBS 0.100418f
C860 digital_0.S3.n19 VSUBS 2.61326f
C861 digital_0.S3.n20 VSUBS 0.701352f
C862 digital_0.S3.n21 VSUBS 0.813614f
C863 TRIM3.t2 VSUBS 0.866601f
C864 TRIM3.n0 VSUBS 0.763327f
C865 TRIM3.t0 VSUBS 0.866499f
C866 TRIM3.n1 VSUBS 2.3023f
C867 TRIM3.t1 VSUBS 0.866499f
C868 TRIM3.n2 VSUBS 0.763327f
C869 TRIM3.t3 VSUBS 0.866543f
C870 DVSS.n0 VSUBS 0.062842f
C871 DVSS.n1 VSUBS 0.05501f
C872 DVSS.n2 VSUBS 0.872992f
C873 DVSS.n3 VSUBS 0.117666f
C874 DVSS.n4 VSUBS 0.181602f
C875 DVSS.n5 VSUBS 0.935831f
C876 DVSS.n6 VSUBS 0.05501f
C877 DVSS.n7 VSUBS 0.05501f
C878 DVSS.n8 VSUBS 0.181602f
C879 DVSS.n9 VSUBS 0.117666f
C880 DVSS.n10 VSUBS 0.117666f
C881 DVSS.n11 VSUBS 0.117666f
C882 DVSS.n12 VSUBS 0.117666f
C883 DVSS.n13 VSUBS 1.97221f
C884 DVSS.t8 VSUBS 2.45172f
C885 DVSS.n14 VSUBS 0.083891f
C886 DVSS.t6 VSUBS 1.87166f
C887 DVSS.t3 VSUBS 0.997704f
C888 DVSS.t4 VSUBS 1.51916f
C889 DVSS.t1 VSUBS 2.33571f
C890 DVSS.n15 VSUBS 1.46175f
C891 DVSS.n16 VSUBS 0.083891f
C892 DVSS.n17 VSUBS 0.083891f
C893 DVSS.n18 VSUBS 0.085084f
C894 DVSS.n19 VSUBS 0.085084f
C895 DVSS.n20 VSUBS 0.077681f
C896 DVSS.n21 VSUBS 0.048524f
C897 DVSS.n22 VSUBS 0.085084f
C898 DVSS.n23 VSUBS 1.97221f
C899 DVSS.n24 VSUBS 0.125313f
C900 DVSS.n25 VSUBS 0.117666f
C901 DVSS.n26 VSUBS 0.090986f
C902 DVSS.n27 VSUBS 0.119123f
C903 DVSS.n28 VSUBS 0.119123f
C904 DVSS.t5 VSUBS 0.600507f
C905 DVSS.n29 VSUBS 0.083891f
C906 DVSS.t2 VSUBS 2.33571f
C907 DVSS.t7 VSUBS 2.45172f
C908 DVSS.t9 VSUBS 1.87166f
C909 DVSS.t0 VSUBS 0.997704f
C910 DVSS.n30 VSUBS 1.46175f
C911 DVSS.n31 VSUBS 0.083891f
C912 DVSS.n32 VSUBS 0.083891f
C913 DVSS.n33 VSUBS 0.085084f
C914 DVSS.n34 VSUBS 0.048524f
C915 DVSS.n35 VSUBS 0.077681f
C916 DVSS.n36 VSUBS 0.085084f
C917 DVSS.n37 VSUBS 0.085084f
C918 DVSS.n38 VSUBS 1.14638f
C919 DVSS.n39 VSUBS 0.117666f
C920 DVSS.n40 VSUBS 0.146304f
C921 DVSS.n41 VSUBS 0.119123f
C922 DVSS.n42 VSUBS 0.117666f
C923 DVSS.n43 VSUBS 0.05501f
C924 DVSS.n44 VSUBS 0.05501f
C925 DVSS.n45 VSUBS 0.119123f
C926 DVSS.n46 VSUBS 0.943565f
C927 DVSS.n47 VSUBS 0.05501f
C928 DVSS.n48 VSUBS 0.05501f
C929 DVSS.n49 VSUBS 0.117666f
C930 DVSS.n50 VSUBS 0.062842f
C931 DVSS.n51 VSUBS 0.125313f
C932 DVSS.n52 VSUBS 1.71698f
C933 DVSS.n53 VSUBS 0.125313f
C934 DVSS.n54 VSUBS 0.062842f
C935 DVSS.n55 VSUBS 0.117481f
C936 DVSS.n56 VSUBS 0.05501f
C937 DVSS.n57 VSUBS 0.117481f
C938 DVSS.n58 VSUBS 0.118937f
C939 DVSS.n59 VSUBS 0.119123f
C940 DVSS.n60 VSUBS 0.943565f
C941 DVSS.n61 VSUBS 0.119123f
C942 DVSS.n62 VSUBS 0.062596f
C943 DVSS.n63 VSUBS 0.117481f
C944 digital_0.S1.t55 VSUBS 0.106315f
C945 digital_0.S1.t59 VSUBS 0.103755f
C946 digital_0.S1.n0 VSUBS 0.879423f
C947 digital_0.S1.t9 VSUBS 0.103835f
C948 digital_0.S1.n1 VSUBS 0.449487f
C949 digital_0.S1.t26 VSUBS 0.103755f
C950 digital_0.S1.n2 VSUBS 0.487031f
C951 digital_0.S1.n3 VSUBS 0.306029f
C952 digital_0.S1.t7 VSUBS 0.103755f
C953 digital_0.S1.t0 VSUBS 0.106315f
C954 digital_0.S1.n4 VSUBS 1.56388f
C955 digital_0.S1.t12 VSUBS 0.066388f
C956 digital_0.S1.t14 VSUBS 0.06353f
C957 digital_0.S1.n5 VSUBS 0.852016f
C958 digital_0.S1.t28 VSUBS 0.0644f
C959 digital_0.S1.t27 VSUBS 0.064324f
C960 digital_0.S1.t2 VSUBS 0.068571f
C961 digital_0.S1.t54 VSUBS 0.065521f
C962 digital_0.S1.n6 VSUBS 0.90788f
C963 digital_0.S1.t16 VSUBS 0.065592f
C964 digital_0.S1.n7 VSUBS 0.463785f
C965 digital_0.S1.t25 VSUBS 0.065521f
C966 digital_0.S1.n8 VSUBS 0.463856f
C967 digital_0.S1.t17 VSUBS 0.065592f
C968 digital_0.S1.n9 VSUBS 0.463785f
C969 digital_0.S1.t56 VSUBS 0.065521f
C970 digital_0.S1.n10 VSUBS 0.475864f
C971 digital_0.S1.t24 VSUBS 0.066456f
C972 digital_0.S1.t43 VSUBS 0.06361f
C973 digital_0.S1.n11 VSUBS 0.851869f
C974 digital_0.S1.t23 VSUBS 0.066388f
C975 digital_0.S1.t42 VSUBS 0.06353f
C976 digital_0.S1.n12 VSUBS 0.852016f
C977 digital_0.S1.t35 VSUBS 0.0644f
C978 digital_0.S1.t34 VSUBS 0.064324f
C979 digital_0.S1.t58 VSUBS 0.073113f
C980 digital_0.S1.t3 VSUBS 0.065521f
C981 digital_0.S1.n13 VSUBS 0.977513f
C982 digital_0.S1.n14 VSUBS 0.817366f
C983 digital_0.S1.n15 VSUBS 0.795403f
C984 digital_0.S1.n16 VSUBS 0.383231f
C985 digital_0.S1.n17 VSUBS 0.371223f
C986 digital_0.S1.n18 VSUBS 0.052805f
C987 digital_0.S1.n19 VSUBS 0.620151f
C988 digital_0.S1.t36 VSUBS 0.106315f
C989 digital_0.S1.t20 VSUBS 0.103755f
C990 digital_0.S1.n20 VSUBS 1.51444f
C991 digital_0.S1.n21 VSUBS 0.842469f
C992 digital_0.S1.n22 VSUBS 0.531357f
C993 digital_0.S1.n23 VSUBS 0.632082f
C994 digital_0.S1.n24 VSUBS 0.21991f
C995 digital_0.S1.t13 VSUBS 0.066456f
C996 digital_0.S1.t15 VSUBS 0.06361f
C997 digital_0.S1.n25 VSUBS 0.851869f
C998 digital_0.S1.t10 VSUBS 0.068571f
C999 digital_0.S1.t33 VSUBS 0.065521f
C1000 digital_0.S1.n26 VSUBS 0.90788f
C1001 digital_0.S1.t11 VSUBS 0.065592f
C1002 digital_0.S1.n27 VSUBS 0.463785f
C1003 digital_0.S1.t8 VSUBS 0.065521f
C1004 digital_0.S1.n28 VSUBS 0.463856f
C1005 digital_0.S1.t37 VSUBS 0.065592f
C1006 digital_0.S1.n29 VSUBS 0.463785f
C1007 digital_0.S1.t29 VSUBS 0.065521f
C1008 digital_0.S1.n30 VSUBS 0.475864f
C1009 digital_0.S1.t4 VSUBS 0.064324f
C1010 digital_0.S1.t5 VSUBS 0.0644f
C1011 digital_0.S1.t18 VSUBS 0.066388f
C1012 digital_0.S1.t21 VSUBS 0.06353f
C1013 digital_0.S1.n31 VSUBS 0.852016f
C1014 digital_0.S1.t19 VSUBS 0.066456f
C1015 digital_0.S1.t22 VSUBS 0.06361f
C1016 digital_0.S1.n32 VSUBS 0.851869f
C1017 digital_0.S1.t32 VSUBS 0.072923f
C1018 digital_0.S1.t57 VSUBS 0.064537f
C1019 digital_0.S1.t38 VSUBS 0.067127f
C1020 digital_0.S1.t45 VSUBS 0.067127f
C1021 digital_0.S1.n33 VSUBS 0.160753f
C1022 digital_0.S1.t40 VSUBS 0.067127f
C1023 digital_0.S1.t50 VSUBS 0.067127f
C1024 digital_0.S1.n34 VSUBS 0.163002f
C1025 digital_0.S1.t39 VSUBS 0.067127f
C1026 digital_0.S1.n35 VSUBS 0.163364f
C1027 digital_0.S1.t41 VSUBS 0.067127f
C1028 digital_0.S1.n36 VSUBS 0.163364f
C1029 digital_0.S1.t53 VSUBS 0.321686f
C1030 digital_0.S1.t48 VSUBS 0.321686f
C1031 digital_0.S1.t47 VSUBS 0.106316f
C1032 digital_0.S1.t52 VSUBS 0.106316f
C1033 digital_0.S1.n37 VSUBS 0.114214f
C1034 digital_0.S1.n38 VSUBS 0.842683f
C1035 digital_0.S1.n39 VSUBS 0.822513f
C1036 digital_0.S1.n40 VSUBS 0.463588f
C1037 digital_0.S1.t51 VSUBS 0.25423f
C1038 digital_0.S1.t46 VSUBS 0.25423f
C1039 digital_0.S1.t44 VSUBS 0.106316f
C1040 digital_0.S1.t49 VSUBS 0.106316f
C1041 digital_0.S1.n41 VSUBS 0.114214f
C1042 digital_0.S1.n42 VSUBS 0.835877f
C1043 digital_0.S1.n43 VSUBS 0.057669f
C1044 digital_0.S1.t31 VSUBS 0.067127f
C1045 digital_0.S1.t6 VSUBS 0.067127f
C1046 digital_0.S1.n44 VSUBS 0.180177f
C1047 digital_0.S1.n45 VSUBS 0.26108f
C1048 digital_0.S1.t30 VSUBS 0.067127f
C1049 digital_0.S1.t1 VSUBS 0.067127f
C1050 digital_0.S1.n46 VSUBS 0.151598f
C1051 digital_0.S1.n47 VSUBS 0.628139f
C1052 digital_0.S1.n48 VSUBS 4.19285f
C1053 digital_0.S1.n49 VSUBS 0.477357f
C1054 digital_0.S1.n50 VSUBS 0.383231f
C1055 digital_0.S1.n51 VSUBS 0.795403f
C1056 digital_0.S1.n52 VSUBS 0.783472f
C1057 digital_0.S1.n53 VSUBS 0.052805f
C1058 digital_0.S1.n54 VSUBS 0.207902f
C1059 digital_0.S1.n55 VSUBS 0.531357f
C1060 digital_0.S1.n56 VSUBS 0.838319f
C1061 bjt_0.B.t31 VSUBS 0.03072f
C1062 bjt_0.B.t30 VSUBS 0.03072f
C1063 bjt_0.B.n0 VSUBS 0.069378f
C1064 bjt_0.B.n1 VSUBS 0.276512f
C1065 bjt_0.B.t12 VSUBS 0.030413f
C1066 bjt_0.B.t10 VSUBS 0.029111f
C1067 bjt_0.B.n2 VSUBS 0.389854f
C1068 bjt_0.B.t16 VSUBS 0.033478f
C1069 bjt_0.B.t4 VSUBS 0.030018f
C1070 bjt_0.B.n3 VSUBS 0.435339f
C1071 bjt_0.B.t40 VSUBS 0.029985f
C1072 bjt_0.B.n4 VSUBS 0.212282f
C1073 bjt_0.B.t18 VSUBS 0.030018f
C1074 bjt_0.B.n5 VSUBS 0.212249f
C1075 bjt_0.B.t17 VSUBS 0.029985f
C1076 bjt_0.B.n6 VSUBS 0.224247f
C1077 bjt_0.B.n7 VSUBS 0.16951f
C1078 bjt_0.B.t9 VSUBS 0.027195f
C1079 bjt_0.B.n8 VSUBS 0.142935f
C1080 bjt_0.B.t11 VSUBS 0.030382f
C1081 bjt_0.B.n9 VSUBS 0.213408f
C1082 bjt_0.B.t33 VSUBS 0.029472f
C1083 bjt_0.B.t32 VSUBS 0.029437f
C1084 bjt_0.B.t37 VSUBS 0.031381f
C1085 bjt_0.B.t19 VSUBS 0.029985f
C1086 bjt_0.B.n10 VSUBS 0.415487f
C1087 bjt_0.B.t15 VSUBS 0.030018f
C1088 bjt_0.B.n11 VSUBS 0.212249f
C1089 bjt_0.B.t6 VSUBS 0.029985f
C1090 bjt_0.B.n12 VSUBS 0.212282f
C1091 bjt_0.B.t34 VSUBS 0.030018f
C1092 bjt_0.B.n13 VSUBS 0.212249f
C1093 bjt_0.B.t5 VSUBS 0.029985f
C1094 bjt_0.B.n14 VSUBS 0.210362f
C1095 bjt_0.B.t0 VSUBS 0.030382f
C1096 bjt_0.B.t13 VSUBS 0.029074f
C1097 bjt_0.B.n15 VSUBS 0.389922f
C1098 bjt_0.B.t43 VSUBS 0.029472f
C1099 bjt_0.B.t42 VSUBS 0.029437f
C1100 bjt_0.B.t3 VSUBS 0.031381f
C1101 bjt_0.B.t8 VSUBS 0.029985f
C1102 bjt_0.B.n16 VSUBS 0.415487f
C1103 bjt_0.B.t41 VSUBS 0.030018f
C1104 bjt_0.B.n17 VSUBS 0.212249f
C1105 bjt_0.B.t7 VSUBS 0.029985f
C1106 bjt_0.B.n18 VSUBS 0.223272f
C1107 bjt_0.B.t36 VSUBS 0.030018f
C1108 bjt_0.B.t2 VSUBS 0.029985f
C1109 bjt_0.B.n19 VSUBS 0.408045f
C1110 bjt_0.B.t35 VSUBS 0.029437f
C1111 bjt_0.B.t38 VSUBS 0.029437f
C1112 bjt_0.B.n20 VSUBS 0.552712f
C1113 bjt_0.B.n21 VSUBS 0.175384f
C1114 bjt_0.B.t39 VSUBS 0.030018f
C1115 bjt_0.B.n22 VSUBS 0.209122f
C1116 bjt_0.B.n23 VSUBS 0.361679f
C1117 bjt_0.B.n24 VSUBS 0.364013f
C1118 bjt_0.B.n25 VSUBS 0.175384f
C1119 bjt_0.B.t14 VSUBS 0.029111f
C1120 bjt_0.B.t1 VSUBS 0.030413f
C1121 bjt_0.B.n26 VSUBS 0.389854f
C1122 bjt_0.B.n27 VSUBS 0.169889f
C1123 bjt_0.B.n28 VSUBS 0.018406f
C1124 bjt_0.B.n29 VSUBS 0.358553f
C1125 bjt_0.B.n30 VSUBS 0.364013f
C1126 bjt_0.B.n31 VSUBS 0.020193f
C1127 bjt_0.B.n32 VSUBS 2.19018f
C1128 bjt_0.B.n33 VSUBS 0.12116f
C1129 bjt_0.B.n34 VSUBS 0.158316f
C1130 bjt_0.B.n35 VSUBS 0.091896f
C1131 bjt_0.B.n36 VSUBS 0.120559f
C1132 bjt_0.B.n37 VSUBS 0.081939f
C1133 bjt_0.B.n38 VSUBS 0.13816f
C1134 bjt_0.B.n39 VSUBS 0.054219f
C1135 bjt_0.B.n41 VSUBS 0.120559f
C1136 bjt_0.B.n42 VSUBS 0.082707f
C1137 bjt_0.B.n43 VSUBS 0.151051f
C1138 bjt_0.B.n44 VSUBS 0.13816f
C1139 bjt_0.B.n45 VSUBS 0.054219f
C1140 bjt_0.B.n47 VSUBS 0.120559f
C1141 bjt_0.B.n48 VSUBS 0.082707f
C1142 bjt_0.B.n49 VSUBS 0.151051f
C1143 bjt_0.B.n50 VSUBS 0.092082f
C1144 bjt_0.B.n51 VSUBS 0.161547f
C1145 bjt_0.B.n52 VSUBS 0.161547f
C1146 bjt_0.B.n55 VSUBS 0.161547f
C1147 bjt_0.B.n56 VSUBS 0.091896f
C1148 bjt_0.B.n57 VSUBS 0.368278f
C1149 bjt_0.B.t22 VSUBS 0.081038f
C1150 bjt_0.B.n58 VSUBS 0.091896f
C1151 bjt_0.B.n59 VSUBS 0.081939f
C1152 bjt_0.B.n60 VSUBS 0.076274f
C1153 bjt_0.B.n61 VSUBS 0.367989f
C1154 bjt_0.B.n62 VSUBS 0.167689f
C1155 bjt_0.B.n63 VSUBS 0.295935f
C1156 bjt_0.B.n65 VSUBS 0.161547f
C1157 bjt_0.B.n66 VSUBS 0.367989f
C1158 bjt_0.B.n67 VSUBS 0.091896f
C1159 bjt_0.B.n68 VSUBS 0.161547f
C1160 bjt_0.B.n69 VSUBS 0.13816f
C1161 bjt_0.B.n70 VSUBS 0.161547f
C1162 bjt_0.B.n71 VSUBS 0.367989f
C1163 bjt_0.B.n72 VSUBS 0.091896f
C1164 bjt_0.B.n73 VSUBS 0.147007f
C1165 bjt_0.B.n74 VSUBS 0.13816f
C1166 bjt_0.B.n76 VSUBS 0.13816f
C1167 bjt_0.B.n77 VSUBS 0.054219f
C1168 bjt_0.B.n78 VSUBS 0.120559f
C1169 bjt_0.B.n79 VSUBS 0.082707f
C1170 bjt_0.B.n80 VSUBS 0.151051f
C1171 bjt_0.B.n81 VSUBS 0.161547f
C1172 bjt_0.B.n82 VSUBS 0.161547f
C1173 bjt_0.B.n84 VSUBS 0.161547f
C1174 bjt_0.B.n86 VSUBS 0.161547f
C1175 bjt_0.B.n87 VSUBS 0.339297f
C1176 bjt_0.B.n88 VSUBS 0.161547f
C1177 bjt_0.B.n89 VSUBS 0.082707f
C1178 bjt_0.B.n90 VSUBS 0.367989f
C1179 bjt_0.B.n91 VSUBS 0.161547f
C1180 bjt_0.B.n92 VSUBS 0.368278f
C1181 bjt_0.B.n93 VSUBS 0.091896f
C1182 bjt_0.B.n94 VSUBS 0.161547f
C1183 bjt_0.B.n95 VSUBS 0.120559f
C1184 bjt_0.B.t25 VSUBS 0.081038f
C1185 bjt_0.B.n96 VSUBS 0.081939f
C1186 bjt_0.B.n97 VSUBS 0.161547f
C1187 bjt_0.B.t26 VSUBS 0.081038f
C1188 bjt_0.B.n98 VSUBS 0.368278f
C1189 bjt_0.B.n99 VSUBS 0.082707f
C1190 bjt_0.B.n100 VSUBS 0.091896f
C1191 bjt_0.B.n101 VSUBS 0.13816f
C1192 bjt_0.B.n102 VSUBS 0.339f
C1193 bjt_0.B.n103 VSUBS 0.322648f
C1194 bjt_0.B.n104 VSUBS 0.331416f
C1195 bjt_0.B.n105 VSUBS 0.376481f
C1196 bjt_0.B.n106 VSUBS 0.367989f
C1197 bjt_0.B.n107 VSUBS 0.076274f
C1198 bjt_0.B.n108 VSUBS 0.054219f
C1199 bjt_0.B.n109 VSUBS 0.161547f
C1200 bjt_0.B.n110 VSUBS 0.161547f
C1201 bjt_0.B.n111 VSUBS 0.082707f
C1202 bjt_0.B.n112 VSUBS 0.091896f
C1203 bjt_0.B.n113 VSUBS 0.13816f
C1204 bjt_0.B.n114 VSUBS 0.339f
C1205 bjt_0.B.n115 VSUBS 0.393558f
C1206 bjt_0.B.n116 VSUBS 0.403211f
C1207 bjt_0.B.n117 VSUBS 0.076274f
C1208 bjt_0.B.n118 VSUBS 0.376481f
C1209 bjt_0.B.n119 VSUBS 0.120559f
C1210 bjt_0.B.n120 VSUBS 0.161547f
C1211 bjt_0.B.n121 VSUBS 0.161547f
C1212 bjt_0.B.n122 VSUBS 0.054219f
C1213 bjt_0.B.n123 VSUBS 0.091896f
C1214 bjt_0.B.n124 VSUBS 0.081939f
C1215 bjt_0.B.t27 VSUBS 0.081038f
C1216 bjt_0.B.n125 VSUBS 0.368278f
C1217 bjt_0.B.n126 VSUBS 0.091896f
C1218 bjt_0.B.n127 VSUBS 0.13816f
C1219 bjt_0.B.n128 VSUBS 0.147007f
C1220 bjt_0.B.n129 VSUBS 0.410105f
C1221 bjt_0.B.n131 VSUBS 0.091896f
C1222 bjt_0.B.n132 VSUBS 0.368278f
C1223 bjt_0.B.t23 VSUBS 0.081038f
C1224 bjt_0.B.n133 VSUBS 0.091896f
C1225 bjt_0.B.n134 VSUBS 0.081939f
C1226 bjt_0.B.n135 VSUBS 0.076274f
C1227 bjt_0.B.n136 VSUBS 0.367989f
C1228 bjt_0.B.n137 VSUBS 0.167689f
C1229 bjt_0.B.n138 VSUBS 0.295935f
C1230 bjt_0.B.n140 VSUBS 0.313763f
C1231 bjt_0.B.n141 VSUBS 0.286357f
C1232 bjt_0.B.n142 VSUBS 0.291999f
C1233 bjt_0.B.n143 VSUBS 0.409253f
C1234 bjt_0.B.n144 VSUBS 0.339297f
C1235 bjt_0.B.n145 VSUBS 0.081939f
C1236 bjt_0.B.t24 VSUBS 0.081038f
C1237 bjt_0.B.n146 VSUBS 0.368278f
C1238 bjt_0.B.n147 VSUBS 0.091896f
C1239 bjt_0.B.n148 VSUBS 0.082707f
C1240 bjt_0.B.n149 VSUBS 0.161547f
C1241 bjt_0.B.n150 VSUBS 0.161547f
C1242 bjt_0.B.n151 VSUBS 0.054219f
C1243 bjt_0.B.n152 VSUBS 0.076274f
C1244 bjt_0.B.n153 VSUBS 0.120559f
C1245 bjt_0.B.n154 VSUBS 0.376481f
C1246 bjt_0.B.n155 VSUBS 0.403211f
C1247 bjt_0.B.n156 VSUBS 0.393558f
C1248 bjt_0.B.n157 VSUBS 0.339f
C1249 bjt_0.B.n158 VSUBS 0.081939f
C1250 bjt_0.B.t20 VSUBS 0.081038f
C1251 bjt_0.B.n159 VSUBS 0.368278f
C1252 bjt_0.B.n160 VSUBS 0.091896f
C1253 bjt_0.B.n161 VSUBS 0.082707f
C1254 bjt_0.B.n162 VSUBS 0.161547f
C1255 bjt_0.B.n163 VSUBS 0.161547f
C1256 bjt_0.B.n164 VSUBS 0.054219f
C1257 bjt_0.B.n165 VSUBS 0.076274f
C1258 bjt_0.B.n166 VSUBS 0.120559f
C1259 bjt_0.B.n167 VSUBS 0.376481f
C1260 bjt_0.B.n168 VSUBS 0.400906f
C1261 bjt_0.B.n169 VSUBS 0.219913f
C1262 bjt_0.B.n170 VSUBS 0.147007f
C1263 bjt_0.B.n171 VSUBS 0.286357f
C1264 bjt_0.B.n172 VSUBS 0.316068f
C1265 bjt_0.B.n173 VSUBS 0.29515f
C1266 bjt_0.B.n174 VSUBS 0.161547f
C1267 bjt_0.B.n175 VSUBS 0.161547f
C1268 bjt_0.B.n177 VSUBS 0.161547f
C1269 bjt_0.B.n180 VSUBS 0.091896f
C1270 bjt_0.B.n181 VSUBS 0.368278f
C1271 bjt_0.B.t21 VSUBS 0.081038f
C1272 bjt_0.B.n182 VSUBS 0.091896f
C1273 bjt_0.B.n183 VSUBS 0.081939f
C1274 bjt_0.B.n184 VSUBS 0.076274f
C1275 bjt_0.B.n185 VSUBS 0.367989f
C1276 bjt_0.B.n186 VSUBS 0.167689f
C1277 bjt_0.B.n187 VSUBS 0.295935f
C1278 bjt_0.B.n189 VSUBS 0.161547f
C1279 bjt_0.B.n190 VSUBS 0.286357f
C1280 bjt_0.B.n191 VSUBS 0.313763f
C1281 bjt_0.B.n192 VSUBS 0.410374f
C1282 bjt_0.B.n193 VSUBS 0.376552f
C1283 bjt_0.B.n194 VSUBS 0.367989f
C1284 bjt_0.B.n195 VSUBS 0.076274f
C1285 bjt_0.B.n196 VSUBS 0.054219f
C1286 bjt_0.B.n197 VSUBS 0.12116f
C1287 bjt_0.B.n198 VSUBS 1.09766f
C1288 bjt_0.B.n199 VSUBS 3.71191f
C1289 bjt_0.B.t29 VSUBS 0.03072f
C1290 bjt_0.B.t28 VSUBS 0.03072f
C1291 bjt_0.B.n200 VSUBS 0.069378f
C1292 bjt_0.B.n201 VSUBS 0.443356f
C1293 TRIM0.t2 VSUBS 0.31673f
C1294 TRIM0.n0 VSUBS 0.278984f
C1295 TRIM0.t0 VSUBS 0.316692f
C1296 TRIM0.n1 VSUBS 0.637208f
C1297 TRIM0.t1 VSUBS 0.316692f
C1298 TRIM0.n2 VSUBS 0.278984f
C1299 TRIM0.t3 VSUBS 0.316671f
C1300 AVSS.n0 VSUBS 0.026777f
C1301 AVSS.n1 VSUBS 0.075408f
C1302 AVSS.n3 VSUBS 0.018889f
C1303 AVSS.n4 VSUBS 0.019048f
C1304 AVSS.n5 VSUBS 0.135542f
C1305 AVSS.n6 VSUBS 0.013197f
C1306 AVSS.n7 VSUBS 0.013464f
C1307 AVSS.n8 VSUBS 0.013197f
C1308 AVSS.n9 VSUBS 0.013464f
C1309 AVSS.n10 VSUBS 0.013197f
C1310 AVSS.n11 VSUBS 0.019496f
C1311 AVSS.n12 VSUBS 0.013197f
C1312 AVSS.n13 VSUBS 0.013464f
C1313 AVSS.n14 VSUBS 0.33097f
C1314 AVSS.n15 VSUBS 0.218223f
C1315 AVSS.n16 VSUBS 0.013464f
C1316 AVSS.n17 VSUBS 0.013197f
C1317 AVSS.n18 VSUBS 0.013464f
C1318 AVSS.n19 VSUBS 0.144269f
C1319 AVSS.n20 VSUBS 0.205976f
C1320 AVSS.n21 VSUBS 0.205814f
C1321 AVSS.n22 VSUBS 0.046257f
C1322 AVSS.n23 VSUBS 0.090352f
C1323 AVSS.n24 VSUBS 0.033817f
C1324 AVSS.n25 VSUBS 0.090352f
C1325 AVSS.n26 VSUBS 0.205976f
C1326 AVSS.n27 VSUBS 0.051397f
C1327 AVSS.n28 VSUBS 0.090352f
C1328 AVSS.n29 VSUBS 0.067428f
C1329 AVSS.n30 VSUBS 0.045828f
C1330 AVSS.n31 VSUBS 0.109298f
C1331 AVSS.n32 VSUBS 0.043695f
C1332 AVSS.n33 VSUBS 0.084482f
C1333 AVSS.n34 VSUBS 0.036625f
C1334 AVSS.n35 VSUBS 0.046257f
C1335 AVSS.n36 VSUBS 0.183064f
C1336 AVSS.n37 VSUBS 0.144269f
C1337 AVSS.n38 VSUBS 0.205814f
C1338 AVSS.n39 VSUBS 0.031241f
C1339 AVSS.n40 VSUBS 0.0343f
C1340 AVSS.n41 VSUBS 0.045173f
C1341 AVSS.n42 VSUBS 0.033852f
C1342 AVSS.n43 VSUBS 0.165515f
C1343 AVSS.n44 VSUBS 0.048186f
C1344 AVSS.n45 VSUBS 0.052903f
C1345 AVSS.n46 VSUBS 0.089808f
C1346 AVSS.n47 VSUBS 0.165515f
C1347 AVSS.n48 VSUBS 0.048186f
C1348 AVSS.n49 VSUBS 0.052903f
C1349 AVSS.n50 VSUBS 0.089808f
C1350 AVSS.n51 VSUBS 0.165515f
C1351 AVSS.n52 VSUBS 0.048186f
C1352 AVSS.n53 VSUBS 0.052903f
C1353 AVSS.n54 VSUBS 0.117889f
C1354 AVSS.n55 VSUBS 0.01633f
C1355 AVSS.n58 VSUBS 0.015203f
C1356 AVSS.n99 VSUBS 0.010886f
C1357 AVSS.n100 VSUBS 0.010886f
C1358 AVSS.n101 VSUBS 0.013002f
C1359 AVSS.n102 VSUBS 0.013002f
C1360 AVSS.n117 VSUBS 0.013536f
C1361 AVSS.n118 VSUBS 0.013536f
C1362 AVSS.n119 VSUBS 0.014085f
C1363 AVSS.n120 VSUBS 0.014085f
C1364 AVSS.n135 VSUBS 0.014104f
C1365 AVSS.n136 VSUBS 0.014104f
C1366 AVSS.n137 VSUBS 0.015863f
C1367 AVSS.n138 VSUBS 0.015863f
C1368 AVSS.t83 VSUBS 1.58362f
C1369 AVSS.n144 VSUBS 0.014231f
C1370 AVSS.n146 VSUBS 0.011838f
C1371 AVSS.n147 VSUBS 0.025184f
C1372 AVSS.n148 VSUBS 0.01756f
C1373 AVSS.n149 VSUBS 0.013197f
C1374 AVSS.n151 VSUBS 0.863324f
C1375 AVSS.n152 VSUBS 0.013464f
C1376 AVSS.n153 VSUBS 0.013197f
C1377 AVSS.n155 VSUBS 0.013464f
C1378 AVSS.n156 VSUBS 0.013197f
C1379 AVSS.n158 VSUBS 0.017327f
C1380 AVSS.n159 VSUBS 0.013197f
C1381 AVSS.n160 VSUBS 0.013464f
C1382 AVSS.n161 VSUBS 0.030665f
C1383 AVSS.n162 VSUBS 0.027461f
C1384 AVSS.n163 VSUBS 0.013464f
C1385 AVSS.n164 VSUBS 0.013197f
C1386 AVSS.n165 VSUBS 0.013464f
C1387 AVSS.n166 VSUBS 0.135542f
C1388 AVSS.n167 VSUBS 0.212363f
C1389 AVSS.n168 VSUBS 0.167359f
C1390 AVSS.n169 VSUBS 0.027461f
C1391 AVSS.n170 VSUBS 0.013464f
C1392 AVSS.n171 VSUBS 0.013197f
C1393 AVSS.n172 VSUBS 0.013464f
C1394 AVSS.n173 VSUBS 0.028377f
C1395 AVSS.n174 VSUBS 0.014676f
C1396 AVSS.n175 VSUBS 0.013197f
C1397 AVSS.n176 VSUBS 0.013464f
C1398 AVSS.n177 VSUBS 0.253149f
C1399 AVSS.n178 VSUBS 0.013464f
C1400 AVSS.n179 VSUBS 0.013197f
C1401 AVSS.n180 VSUBS 0.013464f
C1402 AVSS.n181 VSUBS 0.013197f
C1403 AVSS.n182 VSUBS 0.013464f
C1404 AVSS.n183 VSUBS 0.253149f
C1405 AVSS.n184 VSUBS 0.013464f
C1406 AVSS.n185 VSUBS 0.020848f
C1407 AVSS.n186 VSUBS 0.021194f
C1408 AVSS.n187 VSUBS 0.205976f
C1409 AVSS.n188 VSUBS 0.045828f
C1410 AVSS.n189 VSUBS 0.205976f
C1411 AVSS.n190 VSUBS 0.045828f
C1412 AVSS.n191 VSUBS 0.205976f
C1413 AVSS.n192 VSUBS 0.045828f
C1414 AVSS.n193 VSUBS 0.205976f
C1415 AVSS.n194 VSUBS 0.045828f
C1416 AVSS.n195 VSUBS 0.205976f
C1417 AVSS.n196 VSUBS 0.045828f
C1418 AVSS.n197 VSUBS 0.135542f
C1419 AVSS.n198 VSUBS 0.383942f
C1420 AVSS.n199 VSUBS 0.302372f
C1421 AVSS.n200 VSUBS 0.135542f
C1422 AVSS.n201 VSUBS 0.135542f
C1423 AVSS.n202 VSUBS 0.302372f
C1424 AVSS.n203 VSUBS 0.135542f
C1425 AVSS.n204 VSUBS 0.135542f
C1426 AVSS.n205 VSUBS 0.302372f
C1427 AVSS.n206 VSUBS 0.383942f
C1428 AVSS.n207 VSUBS 0.135542f
C1429 AVSS.n208 VSUBS 0.135542f
C1430 AVSS.n209 VSUBS 0.302372f
C1431 AVSS.n210 VSUBS 0.253149f
C1432 AVSS.n211 VSUBS 0.021194f
C1433 AVSS.n212 VSUBS 0.013464f
C1434 AVSS.n213 VSUBS 0.020848f
C1435 AVSS.n214 VSUBS 0.013197f
C1436 AVSS.n215 VSUBS 0.013464f
C1437 AVSS.n216 VSUBS 0.212363f
C1438 AVSS.n217 VSUBS 0.013464f
C1439 AVSS.n218 VSUBS 0.013197f
C1440 AVSS.n219 VSUBS 0.013464f
C1441 AVSS.t102 VSUBS 0.243736f
C1442 AVSS.n220 VSUBS 0.253149f
C1443 AVSS.n221 VSUBS 0.013464f
C1444 AVSS.n222 VSUBS 0.013197f
C1445 AVSS.n223 VSUBS 0.014676f
C1446 AVSS.n224 VSUBS 0.013197f
C1447 AVSS.n225 VSUBS 0.013464f
C1448 AVSS.n226 VSUBS 0.013197f
C1449 AVSS.n227 VSUBS 0.013464f
C1450 AVSS.n229 VSUBS 0.017327f
C1451 AVSS.n230 VSUBS 0.017108f
C1452 AVSS.n231 VSUBS 0.075481f
C1453 AVSS.n232 VSUBS 0.017925f
C1454 AVSS.n233 VSUBS 0.013197f
C1455 AVSS.n234 VSUBS 0.013464f
C1456 AVSS.n235 VSUBS 0.013197f
C1457 AVSS.n236 VSUBS 0.013464f
C1458 AVSS.n237 VSUBS 0.013197f
C1459 AVSS.n239 VSUBS 0.013464f
C1460 AVSS.n241 VSUBS 0.013464f
C1461 AVSS.n242 VSUBS 0.013197f
C1462 AVSS.n243 VSUBS 0.013197f
C1463 AVSS.n244 VSUBS 0.013197f
C1464 AVSS.n245 VSUBS 0.013464f
C1465 AVSS.n247 VSUBS 0.013464f
C1466 AVSS.n249 VSUBS 0.013464f
C1467 AVSS.n250 VSUBS 0.013197f
C1468 AVSS.n251 VSUBS 0.013197f
C1469 AVSS.n252 VSUBS 0.013197f
C1470 AVSS.n253 VSUBS 0.013464f
C1471 AVSS.n255 VSUBS 0.013464f
C1472 AVSS.n256 VSUBS 0.019496f
C1473 AVSS.n257 VSUBS 0.021345f
C1474 AVSS.n259 VSUBS 0.013464f
C1475 AVSS.n262 VSUBS 0.018072f
C1476 AVSS.n263 VSUBS 0.192186f
C1477 AVSS.n264 VSUBS 0.058887f
C1478 AVSS.n265 VSUBS 0.077272f
C1479 AVSS.n266 VSUBS 0.030324f
C1480 AVSS.n267 VSUBS 0.04266f
C1481 AVSS.n268 VSUBS 0.205814f
C1482 AVSS.n269 VSUBS 0.211571f
C1483 AVSS.n270 VSUBS 0.067428f
C1484 AVSS.n271 VSUBS 0.051397f
C1485 AVSS.n272 VSUBS 0.051397f
C1486 AVSS.n273 VSUBS 0.046257f
C1487 AVSS.n275 VSUBS 0.053722f
C1488 AVSS.n276 VSUBS 0.068875f
C1489 AVSS.n277 VSUBS 0.084482f
C1490 AVSS.t68 VSUBS 19.7724f
C1491 AVSS.t64 VSUBS 18.4555f
C1492 AVSS.t67 VSUBS 32.52f
C1493 AVSS.t54 VSUBS 18.0884f
C1494 AVSS.n279 VSUBS 1.87162f
C1495 AVSS.t69 VSUBS 17.454802f
C1496 AVSS.t66 VSUBS 18.996801f
C1497 AVSS.t65 VSUBS 17.1225f
C1498 AVSS.n280 VSUBS 15.921201f
C1499 AVSS.t60 VSUBS 18.0884f
C1500 AVSS.n281 VSUBS 1.93621f
C1501 AVSS.t59 VSUBS 17.1225f
C1502 AVSS.n282 VSUBS 15.386299f
C1503 AVSS.t58 VSUBS 18.0884f
C1504 AVSS.n283 VSUBS 1.93431f
C1505 AVSS.t57 VSUBS 17.1225f
C1506 AVSS.n284 VSUBS 15.386299f
C1507 AVSS.t56 VSUBS 18.0884f
C1508 AVSS.t72 VSUBS 18.0884f
C1509 AVSS.n285 VSUBS 1.89159f
C1510 AVSS.n286 VSUBS 1.89841f
C1511 AVSS.t43 VSUBS 0.016087f
C1512 AVSS.t41 VSUBS 0.016087f
C1513 AVSS.n288 VSUBS 0.112879f
C1514 AVSS.n289 VSUBS 0.10409f
C1515 AVSS.t29 VSUBS 0.01689f
C1516 AVSS.n290 VSUBS 0.511197f
C1517 AVSS.n291 VSUBS 0.584938f
C1518 AVSS.n292 VSUBS 0.584938f
C1519 AVSS.n293 VSUBS 1.52709f
C1520 AVSS.n294 VSUBS 1.52163f
C1521 AVSS.t16 VSUBS 22.5751f
C1522 AVSS.n295 VSUBS 3.13518f
C1523 AVSS.n296 VSUBS 0.019986f
C1524 AVSS.n297 VSUBS 0.014646f
C1525 AVSS.n298 VSUBS 6.25128f
C1526 AVSS.n299 VSUBS 0.582149f
C1527 AVSS.n300 VSUBS 0.021345f
C1528 AVSS.n301 VSUBS 0.013464f
C1529 AVSS.n302 VSUBS 0.021004f
C1530 AVSS.n303 VSUBS 0.013197f
C1531 AVSS.n304 VSUBS 0.013464f
C1532 AVSS.n305 VSUBS 0.488358f
C1533 AVSS.n306 VSUBS 0.013464f
C1534 AVSS.n307 VSUBS 0.013197f
C1535 AVSS.n308 VSUBS 0.013464f
C1536 AVSS.t104 VSUBS 0.255169f
C1537 AVSS.n309 VSUBS 0.218223f
C1538 AVSS.n310 VSUBS 0.013464f
C1539 AVSS.n311 VSUBS 0.013197f
C1540 AVSS.n312 VSUBS 0.013464f
C1541 AVSS.n313 VSUBS 0.527322f
C1542 AVSS.n314 VSUBS 0.014835f
C1543 AVSS.n315 VSUBS 0.013197f
C1544 AVSS.n317 VSUBS 0.135542f
C1545 AVSS.n318 VSUBS 0.013464f
C1546 AVSS.n321 VSUBS 0.013464f
C1547 AVSS.n324 VSUBS 0.016888f
C1548 AVSS.n327 VSUBS 0.013464f
C1549 AVSS.t90 VSUBS 0.981716f
C1550 AVSS.n340 VSUBS 0.019048f
C1551 AVSS.n346 VSUBS 0.257281f
C1552 AVSS.n347 VSUBS 0.013464f
C1553 AVSS.n348 VSUBS 0.013197f
C1554 AVSS.n349 VSUBS 0.013464f
C1555 AVSS.n350 VSUBS 0.19582f
C1556 AVSS.n351 VSUBS 0.013464f
C1557 AVSS.n352 VSUBS 0.013197f
C1558 AVSS.n353 VSUBS 0.013464f
C1559 AVSS.n354 VSUBS 0.257281f
C1560 AVSS.n355 VSUBS 0.013464f
C1561 AVSS.n356 VSUBS 0.257281f
C1562 AVSS.n357 VSUBS 0.013464f
C1563 AVSS.n358 VSUBS 0.013197f
C1564 AVSS.n359 VSUBS 0.013197f
C1565 AVSS.n360 VSUBS 0.013197f
C1566 AVSS.n361 VSUBS 0.013464f
C1567 AVSS.n362 VSUBS 0.257281f
C1568 AVSS.n363 VSUBS 0.257281f
C1569 AVSS.n364 VSUBS 0.190102f
C1570 AVSS.n365 VSUBS 0.013464f
C1571 AVSS.n366 VSUBS 0.013197f
C1572 AVSS.n367 VSUBS 0.013197f
C1573 AVSS.n368 VSUBS 0.013197f
C1574 AVSS.n369 VSUBS 0.013464f
C1575 AVSS.n370 VSUBS 0.257281f
C1576 AVSS.n371 VSUBS 0.257281f
C1577 AVSS.n372 VSUBS 0.257281f
C1578 AVSS.n373 VSUBS 0.013464f
C1579 AVSS.n374 VSUBS 0.013197f
C1580 AVSS.n375 VSUBS 0.013197f
C1581 AVSS.n376 VSUBS 0.010705f
C1582 AVSS.n377 VSUBS 0.013197f
C1583 AVSS.n378 VSUBS 0.013464f
C1584 AVSS.n379 VSUBS 0.013464f
C1585 AVSS.n380 VSUBS 0.013197f
C1586 AVSS.n381 VSUBS 0.013197f
C1587 AVSS.n382 VSUBS 0.013464f
C1588 AVSS.n383 VSUBS 0.013464f
C1589 AVSS.n384 VSUBS 0.013197f
C1590 AVSS.n385 VSUBS 0.013197f
C1591 AVSS.n386 VSUBS 0.013464f
C1592 AVSS.n387 VSUBS 0.013464f
C1593 AVSS.n388 VSUBS 0.013197f
C1594 AVSS.n389 VSUBS 0.013197f
C1595 AVSS.n390 VSUBS 0.013464f
C1596 AVSS.n391 VSUBS 0.013464f
C1597 AVSS.n392 VSUBS 0.013197f
C1598 AVSS.n393 VSUBS 0.013464f
C1599 AVSS.n394 VSUBS 0.013197f
C1600 AVSS.n395 VSUBS 0.018889f
C1601 AVSS.n396 VSUBS 0.020848f
C1602 AVSS.n397 VSUBS 0.021194f
C1603 AVSS.n398 VSUBS 0.410221f
C1604 AVSS.n399 VSUBS 1.57993f
C1605 AVSS.n406 VSUBS 0.021194f
C1606 AVSS.n407 VSUBS 0.013464f
C1607 AVSS.n408 VSUBS 0.018062f
C1608 AVSS.n409 VSUBS 0.011763f
C1609 AVSS.n410 VSUBS 0.013464f
C1610 AVSS.n416 VSUBS 0.218223f
C1611 AVSS.n417 VSUBS 0.013464f
C1612 AVSS.n418 VSUBS 0.014835f
C1613 AVSS.n419 VSUBS 0.013197f
C1614 AVSS.n420 VSUBS 0.033817f
C1615 AVSS.n421 VSUBS 0.013197f
C1616 AVSS.n422 VSUBS 0.013464f
C1617 AVSS.n427 VSUBS 0.013464f
C1618 AVSS.n428 VSUBS 0.019496f
C1619 AVSS.n429 VSUBS 0.013197f
C1620 AVSS.n430 VSUBS 0.013464f
C1621 AVSS.n431 VSUBS 0.33097f
C1622 AVSS.n432 VSUBS 0.218223f
C1623 AVSS.n433 VSUBS 0.013464f
C1624 AVSS.n434 VSUBS 0.013197f
C1625 AVSS.n435 VSUBS 0.013464f
C1626 AVSS.n436 VSUBS 0.218223f
C1627 AVSS.n437 VSUBS 0.013464f
C1628 AVSS.n438 VSUBS 0.013197f
C1629 AVSS.n439 VSUBS 0.013464f
C1630 AVSS.n440 VSUBS 0.218223f
C1631 AVSS.n441 VSUBS 0.218223f
C1632 AVSS.n442 VSUBS 0.013464f
C1633 AVSS.n443 VSUBS 0.013197f
C1634 AVSS.n444 VSUBS 0.013197f
C1635 AVSS.n445 VSUBS 0.013197f
C1636 AVSS.n446 VSUBS 0.013464f
C1637 AVSS.n447 VSUBS 0.218223f
C1638 AVSS.n448 VSUBS 0.144269f
C1639 AVSS.n449 VSUBS 0.205976f
C1640 AVSS.n450 VSUBS 0.205814f
C1641 AVSS.n451 VSUBS 0.046257f
C1642 AVSS.n452 VSUBS 0.043547f
C1643 AVSS.n453 VSUBS 0.098567f
C1644 AVSS.n454 VSUBS 0.205814f
C1645 AVSS.n455 VSUBS 0.045828f
C1646 AVSS.n456 VSUBS 0.051397f
C1647 AVSS.n457 VSUBS 0.031136f
C1648 AVSS.n458 VSUBS 0.034184f
C1649 AVSS.n459 VSUBS 0.040019f
C1650 AVSS.n460 VSUBS 0.077272f
C1651 AVSS.n461 VSUBS 0.085645f
C1652 AVSS.n465 VSUBS 0.013536f
C1653 AVSS.n469 VSUBS 0.010886f
C1654 AVSS.n484 VSUBS 0.015863f
C1655 AVSS.n499 VSUBS 0.013002f
C1656 AVSS.n500 VSUBS 0.013002f
C1657 AVSS.n501 VSUBS 0.010886f
C1658 AVSS.n515 VSUBS 0.014231f
C1659 AVSS.n516 VSUBS 0.014231f
C1660 AVSS.n517 VSUBS 0.015203f
C1661 AVSS.n518 VSUBS 0.015203f
C1662 AVSS.n533 VSUBS 0.015863f
C1663 AVSS.n545 VSUBS 0.014104f
C1664 AVSS.n546 VSUBS 0.014104f
C1665 AVSS.t103 VSUBS 1.58362f
C1666 AVSS.n549 VSUBS 0.014085f
C1667 AVSS.n551 VSUBS 0.010932f
C1668 AVSS.n552 VSUBS 0.017999f
C1669 AVSS.n553 VSUBS 0.025256f
C1670 AVSS.n554 VSUBS 0.014516f
C1671 AVSS.n555 VSUBS 0.033888f
C1672 AVSS.n556 VSUBS 0.077272f
C1673 AVSS.n557 VSUBS 0.030324f
C1674 AVSS.n559 VSUBS 0.067428f
C1675 AVSS.n560 VSUBS 0.046257f
C1676 AVSS.n561 VSUBS 0.084482f
C1677 AVSS.n562 VSUBS 0.131596f
C1678 AVSS.n563 VSUBS 0.0905f
C1679 AVSS.n564 VSUBS 0.0905f
C1680 AVSS.n566 VSUBS 0.0905f
C1681 AVSS.n569 VSUBS 0.051397f
C1682 AVSS.n570 VSUBS 0.205976f
C1683 AVSS.n571 VSUBS 0.205976f
C1684 AVSS.n572 VSUBS 0.205814f
C1685 AVSS.n573 VSUBS 0.046257f
C1686 AVSS.n574 VSUBS 0.066046f
C1687 AVSS.n575 VSUBS 0.067394f
C1688 AVSS.n576 VSUBS 0.067394f
C1689 AVSS.n577 VSUBS 0.051397f
C1690 AVSS.n580 VSUBS 0.077272f
C1691 AVSS.n581 VSUBS 0.04266f
C1692 AVSS.n583 VSUBS 0.093787f
C1693 AVSS.n584 VSUBS 0.067428f
C1694 AVSS.n586 VSUBS 0.084482f
C1695 AVSS.n587 VSUBS 0.160158f
C1696 AVSS.n588 VSUBS 0.075481f
C1697 AVSS.n589 VSUBS 0.030324f
C1698 AVSS.n590 VSUBS 0.051397f
C1699 AVSS.n591 VSUBS 0.045828f
C1700 AVSS.n592 VSUBS 0.135542f
C1701 AVSS.n593 VSUBS 0.135542f
C1702 AVSS.n594 VSUBS 0.135542f
C1703 AVSS.n595 VSUBS 0.135542f
C1704 AVSS.n596 VSUBS 0.135542f
C1705 AVSS.n597 VSUBS 0.135542f
C1706 AVSS.n598 VSUBS 0.135542f
C1707 AVSS.n599 VSUBS 0.135542f
C1708 AVSS.n606 VSUBS 0.019496f
C1709 AVSS.n613 VSUBS 0.019496f
C1710 AVSS.n626 VSUBS 0.019496f
C1711 AVSS.n633 VSUBS 0.013464f
C1712 AVSS.n634 VSUBS 0.014835f
C1713 AVSS.n635 VSUBS 0.013197f
C1714 AVSS.n636 VSUBS 0.013197f
C1715 AVSS.n638 VSUBS 0.013464f
C1716 AVSS.n641 VSUBS 0.013464f
C1717 AVSS.n644 VSUBS 0.016888f
C1718 AVSS.n647 VSUBS 0.013464f
C1719 AVSS.t80 VSUBS 2.06361f
C1720 AVSS.n654 VSUBS 0.019048f
C1721 AVSS.n661 VSUBS 0.019048f
C1722 AVSS.n668 VSUBS 0.028377f
C1723 AVSS.n669 VSUBS 0.013464f
C1724 AVSS.n670 VSUBS 0.014676f
C1725 AVSS.n671 VSUBS 0.013197f
C1726 AVSS.n672 VSUBS 0.013197f
C1727 AVSS.n673 VSUBS 0.013464f
C1728 AVSS.n674 VSUBS 0.027461f
C1729 AVSS.n675 VSUBS 0.013464f
C1730 AVSS.n676 VSUBS 0.013197f
C1731 AVSS.n677 VSUBS 0.013464f
C1732 AVSS.n678 VSUBS 0.027461f
C1733 AVSS.n679 VSUBS 0.013464f
C1734 AVSS.n680 VSUBS 0.014713f
C1735 AVSS.n681 VSUBS 0.014835f
C1736 AVSS.n682 VSUBS 0.013464f
C1737 AVSS.n683 VSUBS 0.01756f
C1738 AVSS.n684 VSUBS 0.020848f
C1739 AVSS.n685 VSUBS 0.013464f
C1740 AVSS.n686 VSUBS 0.013197f
C1741 AVSS.n687 VSUBS 0.013464f
C1742 AVSS.n688 VSUBS 0.013197f
C1743 AVSS.n689 VSUBS 0.013464f
C1744 AVSS.n690 VSUBS 0.019496f
C1745 AVSS.n692 VSUBS 0.021345f
C1746 AVSS.n693 VSUBS 0.021004f
C1747 AVSS.n694 VSUBS 0.013197f
C1748 AVSS.n695 VSUBS 0.013197f
C1749 AVSS.n696 VSUBS 0.013464f
C1750 AVSS.n698 VSUBS 0.013464f
C1751 AVSS.n700 VSUBS 0.013464f
C1752 AVSS.n701 VSUBS 0.013197f
C1753 AVSS.n702 VSUBS 0.013197f
C1754 AVSS.n703 VSUBS 0.013197f
C1755 AVSS.n704 VSUBS 0.013464f
C1756 AVSS.n706 VSUBS 0.013464f
C1757 AVSS.n708 VSUBS 0.013464f
C1758 AVSS.n709 VSUBS 0.013197f
C1759 AVSS.n710 VSUBS 0.013197f
C1760 AVSS.n711 VSUBS 0.013197f
C1761 AVSS.n712 VSUBS 0.013464f
C1762 AVSS.n714 VSUBS 0.021194f
C1763 AVSS.n715 VSUBS 0.019048f
C1764 AVSS.n716 VSUBS 0.017129f
C1765 AVSS.n717 VSUBS 0.013197f
C1766 AVSS.n718 VSUBS 0.013464f
C1767 AVSS.n719 VSUBS 0.013464f
C1768 AVSS.n720 VSUBS 0.013197f
C1769 AVSS.n721 VSUBS 0.013197f
C1770 AVSS.n722 VSUBS 0.013464f
C1771 AVSS.n723 VSUBS 0.013464f
C1772 AVSS.n724 VSUBS 0.013197f
C1773 AVSS.n725 VSUBS 0.013197f
C1774 AVSS.n726 VSUBS 0.013464f
C1775 AVSS.n727 VSUBS 0.013464f
C1776 AVSS.n728 VSUBS 0.013197f
C1777 AVSS.n729 VSUBS 0.013197f
C1778 AVSS.n730 VSUBS 0.013464f
C1779 AVSS.n731 VSUBS 0.013464f
C1780 AVSS.n732 VSUBS 0.013197f
C1781 AVSS.n733 VSUBS 0.013197f
C1782 AVSS.n734 VSUBS 0.013464f
C1783 AVSS.n735 VSUBS 0.013464f
C1784 AVSS.n738 VSUBS 0.01633f
C1785 AVSS.n739 VSUBS 0.075481f
C1786 AVSS.n742 VSUBS 0.015203f
C1787 AVSS.n760 VSUBS 0.015863f
C1788 AVSS.n777 VSUBS 0.012104f
C1789 AVSS.n790 VSUBS 0.010886f
C1790 AVSS.n791 VSUBS 0.010886f
C1791 AVSS.n792 VSUBS 0.013002f
C1792 AVSS.n793 VSUBS 0.013002f
C1793 AVSS.n808 VSUBS 0.013536f
C1794 AVSS.n809 VSUBS 0.013536f
C1795 AVSS.n810 VSUBS 0.014085f
C1796 AVSS.n811 VSUBS 0.014085f
C1797 AVSS.n825 VSUBS 0.010825f
C1798 AVSS.n826 VSUBS 0.014104f
C1799 AVSS.t87 VSUBS 1.58362f
C1800 AVSS.n829 VSUBS 0.014231f
C1801 AVSS.n831 VSUBS 0.011838f
C1802 AVSS.n832 VSUBS 0.075408f
C1803 AVSS.n833 VSUBS 0.018072f
C1804 AVSS.n836 VSUBS 0.013464f
C1805 AVSS.n837 VSUBS 0.013464f
C1806 AVSS.n838 VSUBS 0.013197f
C1807 AVSS.n839 VSUBS 0.013197f
C1808 AVSS.n840 VSUBS 0.013464f
C1809 AVSS.n841 VSUBS 0.013464f
C1810 AVSS.n842 VSUBS 0.013197f
C1811 AVSS.n843 VSUBS 0.013197f
C1812 AVSS.n844 VSUBS 0.013464f
C1813 AVSS.n845 VSUBS 0.013464f
C1814 AVSS.n846 VSUBS 0.013197f
C1815 AVSS.n847 VSUBS 0.013197f
C1816 AVSS.n848 VSUBS 0.013464f
C1817 AVSS.n849 VSUBS 0.013464f
C1818 AVSS.n850 VSUBS 0.013197f
C1819 AVSS.n851 VSUBS 0.013197f
C1820 AVSS.n852 VSUBS 0.013464f
C1821 AVSS.n853 VSUBS 0.013464f
C1822 AVSS.n854 VSUBS 0.013197f
C1823 AVSS.n855 VSUBS 0.013197f
C1824 AVSS.n856 VSUBS 0.017108f
C1825 AVSS.n857 VSUBS 0.017327f
C1826 AVSS.n858 VSUBS 0.030665f
C1827 AVSS.n859 VSUBS 0.029139f
C1828 AVSS.n860 VSUBS 0.027461f
C1829 AVSS.n861 VSUBS 0.013464f
C1830 AVSS.n862 VSUBS 0.013197f
C1831 AVSS.n863 VSUBS 0.013197f
C1832 AVSS.n864 VSUBS 0.013197f
C1833 AVSS.n865 VSUBS 0.013197f
C1834 AVSS.n866 VSUBS 0.013464f
C1835 AVSS.n867 VSUBS 0.027461f
C1836 AVSS.n868 VSUBS 0.027461f
C1837 AVSS.n869 VSUBS 0.020291f
C1838 AVSS.n870 VSUBS 0.013464f
C1839 AVSS.n871 VSUBS 0.020901f
C1840 AVSS.n872 VSUBS 0.013464f
C1841 AVSS.n874 VSUBS 0.012464f
C1842 AVSS.n875 VSUBS 0.013197f
C1843 AVSS.n876 VSUBS 0.013464f
C1844 AVSS.n877 VSUBS 0.027461f
C1845 AVSS.n878 VSUBS 0.027461f
C1846 AVSS.n879 VSUBS 0.027461f
C1847 AVSS.n880 VSUBS 0.013464f
C1848 AVSS.n881 VSUBS 0.013197f
C1849 AVSS.n882 VSUBS 0.014549f
C1850 AVSS.n883 VSUBS 0.016685f
C1851 AVSS.n884 VSUBS 0.016888f
C1852 AVSS.n885 VSUBS 0.030055f
C1853 AVSS.n886 VSUBS 1.57993f
C1854 AVSS.n892 VSUBS 0.021194f
C1855 AVSS.n893 VSUBS 0.013464f
C1856 AVSS.n894 VSUBS 0.013197f
C1857 AVSS.n895 VSUBS 0.013464f
C1858 AVSS.n896 VSUBS 0.013197f
C1859 AVSS.n897 VSUBS 0.013464f
C1860 AVSS.n898 VSUBS 0.013197f
C1861 AVSS.n899 VSUBS 0.019496f
C1862 AVSS.n900 VSUBS 0.013197f
C1863 AVSS.n901 VSUBS 0.013464f
C1864 AVSS.n902 VSUBS 0.013464f
C1865 AVSS.n903 VSUBS 0.013197f
C1866 AVSS.n904 VSUBS 0.013197f
C1867 AVSS.n905 VSUBS 0.013464f
C1868 AVSS.n906 VSUBS 0.013464f
C1869 AVSS.n907 VSUBS 0.013197f
C1870 AVSS.n908 VSUBS 0.013197f
C1871 AVSS.n909 VSUBS 0.013464f
C1872 AVSS.n910 VSUBS 0.013464f
C1873 AVSS.n911 VSUBS 0.013197f
C1874 AVSS.n912 VSUBS 0.013197f
C1875 AVSS.n913 VSUBS 0.013464f
C1876 AVSS.n914 VSUBS 0.013464f
C1877 AVSS.n915 VSUBS 0.013197f
C1878 AVSS.n916 VSUBS 0.013197f
C1879 AVSS.n917 VSUBS 0.013464f
C1880 AVSS.n918 VSUBS 0.013464f
C1881 AVSS.n919 VSUBS 0.013197f
C1882 AVSS.n920 VSUBS 0.01932f
C1883 AVSS.n921 VSUBS 0.021004f
C1884 AVSS.n922 VSUBS 0.021345f
C1885 AVSS.n924 VSUBS 0.013464f
C1886 AVSS.n926 VSUBS 0.013464f
C1887 AVSS.n927 VSUBS 0.013197f
C1888 AVSS.n928 VSUBS 0.013197f
C1889 AVSS.n929 VSUBS 0.013197f
C1890 AVSS.n930 VSUBS 0.013464f
C1891 AVSS.n932 VSUBS 0.013464f
C1892 AVSS.n934 VSUBS 0.013464f
C1893 AVSS.n935 VSUBS 0.013197f
C1894 AVSS.n936 VSUBS 0.013197f
C1895 AVSS.n937 VSUBS 0.013197f
C1896 AVSS.n938 VSUBS 0.013464f
C1897 AVSS.n940 VSUBS 0.013464f
C1898 AVSS.n942 VSUBS 0.013464f
C1899 AVSS.n943 VSUBS 0.013197f
C1900 AVSS.n944 VSUBS 0.020848f
C1901 AVSS.n945 VSUBS 0.010705f
C1902 AVSS.n946 VSUBS 0.013197f
C1903 AVSS.n947 VSUBS 0.013464f
C1904 AVSS.n948 VSUBS 0.013464f
C1905 AVSS.n949 VSUBS 0.013197f
C1906 AVSS.n950 VSUBS 0.013197f
C1907 AVSS.n951 VSUBS 0.013464f
C1908 AVSS.n952 VSUBS 0.013464f
C1909 AVSS.n953 VSUBS 0.013197f
C1910 AVSS.n954 VSUBS 0.013197f
C1911 AVSS.n955 VSUBS 0.013464f
C1912 AVSS.n956 VSUBS 0.013464f
C1913 AVSS.n957 VSUBS 0.013197f
C1914 AVSS.n958 VSUBS 0.013197f
C1915 AVSS.n959 VSUBS 0.013464f
C1916 AVSS.n960 VSUBS 0.013464f
C1917 AVSS.n961 VSUBS 0.013197f
C1918 AVSS.n962 VSUBS 0.013197f
C1919 AVSS.n963 VSUBS 0.018889f
C1920 AVSS.n964 VSUBS 0.019048f
C1921 AVSS.n971 VSUBS 0.021194f
C1922 AVSS.n972 VSUBS 0.013464f
C1923 AVSS.n973 VSUBS 0.018062f
C1924 AVSS.n994 VSUBS 0.015203f
C1925 AVSS.n1007 VSUBS 0.014085f
C1926 AVSS.n1008 VSUBS 0.014085f
C1927 AVSS.n1009 VSUBS 0.013536f
C1928 AVSS.n1010 VSUBS 0.013536f
C1929 AVSS.n1025 VSUBS 0.013002f
C1930 AVSS.n1026 VSUBS 0.013002f
C1931 AVSS.n1027 VSUBS 0.010886f
C1932 AVSS.n1028 VSUBS 0.010886f
C1933 AVSS.n1043 VSUBS 0.014231f
C1934 AVSS.n1044 VSUBS 0.014231f
C1935 AVSS.n1045 VSUBS 0.015203f
C1936 AVSS.n1046 VSUBS 0.015863f
C1937 AVSS.t79 VSUBS 1.58362f
C1938 AVSS.n1063 VSUBS 0.014104f
C1939 AVSS.n1064 VSUBS 0.010825f
C1940 AVSS.n1065 VSUBS 0.012104f
C1941 AVSS.n1066 VSUBS 0.024671f
C1942 AVSS.n1067 VSUBS 0.073869f
C1943 AVSS.n1068 VSUBS 0.01756f
C1944 AVSS.n1069 VSUBS 0.013197f
C1945 AVSS.n1070 VSUBS 0.019496f
C1946 AVSS.n1071 VSUBS 0.863324f
C1947 AVSS.n1072 VSUBS 0.013197f
C1948 AVSS.n1073 VSUBS 0.013464f
C1949 AVSS.n1074 VSUBS 0.013197f
C1950 AVSS.n1076 VSUBS 0.013464f
C1951 AVSS.n1077 VSUBS 0.013197f
C1952 AVSS.n1079 VSUBS 0.014835f
C1953 AVSS.n1080 VSUBS 0.013197f
C1954 AVSS.n1082 VSUBS 0.135542f
C1955 AVSS.n1083 VSUBS 0.013464f
C1956 AVSS.n1086 VSUBS 0.013464f
C1957 AVSS.n1087 VSUBS 0.013197f
C1958 AVSS.n1089 VSUBS 0.016888f
C1959 AVSS.n1090 VSUBS 0.013197f
C1960 AVSS.n1091 VSUBS 0.013464f
C1961 AVSS.n1092 VSUBS 0.205976f
C1962 AVSS.n1093 VSUBS 0.205814f
C1963 AVSS.n1094 VSUBS 0.046257f
C1964 AVSS.n1095 VSUBS 0.066046f
C1965 AVSS.n1096 VSUBS 0.067394f
C1966 AVSS.n1097 VSUBS 0.067394f
C1967 AVSS.n1098 VSUBS 0.051397f
C1968 AVSS.n1101 VSUBS 0.077272f
C1969 AVSS.n1102 VSUBS 0.04266f
C1970 AVSS.n1104 VSUBS 0.093787f
C1971 AVSS.n1105 VSUBS 0.067428f
C1972 AVSS.n1107 VSUBS 0.084482f
C1973 AVSS.n1108 VSUBS 0.160158f
C1974 AVSS.n1109 VSUBS 0.075481f
C1975 AVSS.n1110 VSUBS 0.030324f
C1976 AVSS.n1111 VSUBS 0.051397f
C1977 AVSS.n1112 VSUBS 0.045828f
C1978 AVSS.t78 VSUBS 2.06361f
C1979 AVSS.n1119 VSUBS 0.016888f
C1980 AVSS.n1126 VSUBS 0.019048f
C1981 AVSS.n1132 VSUBS 1.57993f
C1982 AVSS.n1139 VSUBS 0.019048f
C1983 AVSS.n1145 VSUBS 0.019048f
C1984 AVSS.n1146 VSUBS 0.013464f
C1985 AVSS.n1148 VSUBS 0.016685f
C1986 AVSS.n1149 VSUBS 0.014676f
C1987 AVSS.n1150 VSUBS 0.027461f
C1988 AVSS.n1151 VSUBS 0.013464f
C1989 AVSS.n1152 VSUBS 0.012464f
C1990 AVSS.n1153 VSUBS 0.013464f
C1991 AVSS.n1154 VSUBS 0.013197f
C1992 AVSS.n1155 VSUBS 0.013464f
C1993 AVSS.n1156 VSUBS 0.027461f
C1994 AVSS.n1157 VSUBS 0.013464f
C1995 AVSS.n1158 VSUBS 0.017108f
C1996 AVSS.n1160 VSUBS 0.013197f
C1997 AVSS.n1161 VSUBS 0.013464f
C1998 AVSS.n1162 VSUBS 0.013197f
C1999 AVSS.n1163 VSUBS 0.013464f
C2000 AVSS.n1165 VSUBS 0.021345f
C2001 AVSS.n1166 VSUBS 0.013197f
C2002 AVSS.n1167 VSUBS 0.013464f
C2003 AVSS.n1172 VSUBS 0.013464f
C2004 AVSS.n1173 VSUBS 0.017129f
C2005 AVSS.n1174 VSUBS 0.021194f
C2006 AVSS.n1175 VSUBS 0.020848f
C2007 AVSS.n1176 VSUBS 0.013197f
C2008 AVSS.n1177 VSUBS 0.013464f
C2009 AVSS.n1178 VSUBS 0.013464f
C2010 AVSS.n1179 VSUBS 0.013197f
C2011 AVSS.n1180 VSUBS 0.013197f
C2012 AVSS.n1181 VSUBS 0.013464f
C2013 AVSS.n1182 VSUBS 0.013464f
C2014 AVSS.n1183 VSUBS 0.013197f
C2015 AVSS.n1184 VSUBS 0.013197f
C2016 AVSS.n1185 VSUBS 0.013464f
C2017 AVSS.n1186 VSUBS 0.013464f
C2018 AVSS.n1187 VSUBS 0.013197f
C2019 AVSS.n1188 VSUBS 0.013197f
C2020 AVSS.n1189 VSUBS 0.013197f
C2021 AVSS.n1190 VSUBS 0.013464f
C2022 AVSS.n1192 VSUBS 0.135542f
C2023 AVSS.n1194 VSUBS 0.013464f
C2024 AVSS.n1195 VSUBS 0.013197f
C2025 AVSS.n1196 VSUBS 0.021004f
C2026 AVSS.n1197 VSUBS 0.01633f
C2027 AVSS.n1198 VSUBS 0.075481f
C2028 AVSS.n1201 VSUBS 0.015203f
C2029 AVSS.n1219 VSUBS 0.015863f
C2030 AVSS.n1236 VSUBS 0.012104f
C2031 AVSS.n1249 VSUBS 0.010886f
C2032 AVSS.n1250 VSUBS 0.010886f
C2033 AVSS.n1251 VSUBS 0.013002f
C2034 AVSS.n1252 VSUBS 0.013002f
C2035 AVSS.n1267 VSUBS 0.013536f
C2036 AVSS.n1268 VSUBS 0.013536f
C2037 AVSS.n1269 VSUBS 0.014085f
C2038 AVSS.n1270 VSUBS 0.014085f
C2039 AVSS.n1284 VSUBS 0.010825f
C2040 AVSS.n1285 VSUBS 0.014104f
C2041 AVSS.t96 VSUBS 1.58362f
C2042 AVSS.n1288 VSUBS 0.014231f
C2043 AVSS.n1290 VSUBS 0.011838f
C2044 AVSS.n1291 VSUBS 0.075408f
C2045 AVSS.n1292 VSUBS 0.01633f
C2046 AVSS.n1294 VSUBS 0.01756f
C2047 AVSS.n1295 VSUBS 0.019496f
C2048 AVSS.n1297 VSUBS 0.013464f
C2049 AVSS.n1299 VSUBS 0.013464f
C2050 AVSS.n1300 VSUBS 0.013197f
C2051 AVSS.n1301 VSUBS 0.013197f
C2052 AVSS.n1302 VSUBS 0.013197f
C2053 AVSS.n1303 VSUBS 0.013464f
C2054 AVSS.n1305 VSUBS 0.013464f
C2055 AVSS.n1307 VSUBS 0.013464f
C2056 AVSS.n1308 VSUBS 0.013197f
C2057 AVSS.n1309 VSUBS 0.013197f
C2058 AVSS.n1310 VSUBS 0.013197f
C2059 AVSS.n1311 VSUBS 0.013464f
C2060 AVSS.n1313 VSUBS 0.013464f
C2061 AVSS.n1314 VSUBS 0.013464f
C2062 AVSS.n1315 VSUBS 0.013197f
C2063 AVSS.n1316 VSUBS 0.013197f
C2064 AVSS.n1317 VSUBS 0.013464f
C2065 AVSS.n1318 VSUBS 0.017327f
C2066 AVSS.n1319 VSUBS 0.030665f
C2067 AVSS.n1320 VSUBS 0.029139f
C2068 AVSS.n1321 VSUBS 0.014835f
C2069 AVSS.n1322 VSUBS 0.014713f
C2070 AVSS.n1323 VSUBS 0.013197f
C2071 AVSS.n1324 VSUBS 0.013197f
C2072 AVSS.n1325 VSUBS 0.013464f
C2073 AVSS.n1326 VSUBS 0.027461f
C2074 AVSS.n1327 VSUBS 0.027461f
C2075 AVSS.n1328 VSUBS 0.020291f
C2076 AVSS.n1329 VSUBS 0.027461f
C2077 AVSS.n1330 VSUBS 0.013464f
C2078 AVSS.n1331 VSUBS 0.013197f
C2079 AVSS.n1332 VSUBS 0.013197f
C2080 AVSS.n1334 VSUBS 0.013464f
C2081 AVSS.n1335 VSUBS 0.013464f
C2082 AVSS.n1336 VSUBS 0.027461f
C2083 AVSS.n1337 VSUBS 0.013464f
C2084 AVSS.n1338 VSUBS 0.013197f
C2085 AVSS.n1339 VSUBS 0.013197f
C2086 AVSS.n1340 VSUBS 0.014549f
C2087 AVSS.n1341 VSUBS 0.013197f
C2088 AVSS.n1342 VSUBS 0.013464f
C2089 AVSS.n1343 VSUBS 0.027461f
C2090 AVSS.n1344 VSUBS 0.028377f
C2091 AVSS.n1345 VSUBS 0.030055f
C2092 AVSS.n1346 VSUBS 0.016888f
C2093 AVSS.n1347 VSUBS 0.013464f
C2094 AVSS.n1348 VSUBS 0.013197f
C2095 AVSS.n1349 VSUBS 0.013197f
C2096 AVSS.n1350 VSUBS 0.013464f
C2097 AVSS.n1351 VSUBS 0.013464f
C2098 AVSS.n1352 VSUBS 0.013197f
C2099 AVSS.n1353 VSUBS 0.013197f
C2100 AVSS.n1354 VSUBS 0.013464f
C2101 AVSS.n1355 VSUBS 0.013464f
C2102 AVSS.n1356 VSUBS 0.013197f
C2103 AVSS.n1357 VSUBS 0.013197f
C2104 AVSS.n1358 VSUBS 0.013464f
C2105 AVSS.n1359 VSUBS 0.013464f
C2106 AVSS.n1360 VSUBS 0.013197f
C2107 AVSS.n1361 VSUBS 0.013197f
C2108 AVSS.n1362 VSUBS 0.013464f
C2109 AVSS.n1363 VSUBS 0.013464f
C2110 AVSS.n1364 VSUBS 0.013197f
C2111 AVSS.n1365 VSUBS 0.013197f
C2112 AVSS.n1367 VSUBS 0.013464f
C2113 AVSS.n1369 VSUBS 0.013464f
C2114 AVSS.n1370 VSUBS 0.014676f
C2115 AVSS.n1372 VSUBS 0.013197f
C2116 AVSS.n1373 VSUBS 0.013464f
C2117 AVSS.n1378 VSUBS 0.013464f
C2118 AVSS.n1379 VSUBS 0.017108f
C2119 AVSS.n1380 VSUBS 0.013464f
C2120 AVSS.n1381 VSUBS 0.010705f
C2121 AVSS.n1382 VSUBS 0.075481f
C2122 AVSS.n1383 VSUBS 0.010705f
C2123 AVSS.n1384 VSUBS 0.014549f
C2124 AVSS.n1385 VSUBS 0.013464f
C2125 AVSS.n1386 VSUBS 0.012464f
C2126 AVSS.n1387 VSUBS 0.013464f
C2127 AVSS.n1388 VSUBS 0.013197f
C2128 AVSS.n1389 VSUBS 0.013464f
C2129 AVSS.n1393 VSUBS 0.013002f
C2130 AVSS.n1412 VSUBS 0.015863f
C2131 AVSS.n1424 VSUBS 0.014231f
C2132 AVSS.n1425 VSUBS 0.014231f
C2133 AVSS.n1426 VSUBS 0.015203f
C2134 AVSS.n1427 VSUBS 0.015203f
C2135 AVSS.n1442 VSUBS 0.015863f
C2136 AVSS.n1457 VSUBS 0.013536f
C2137 AVSS.n1459 VSUBS 0.010931f
C2138 AVSS.n1461 VSUBS 0.014085f
C2139 AVSS.n1475 VSUBS 0.014104f
C2140 AVSS.n1476 VSUBS 0.014104f
C2141 AVSS.t86 VSUBS 1.58362f
C2142 AVSS.n1478 VSUBS 0.010886f
C2143 AVSS.n1481 VSUBS 0.075408f
C2144 AVSS.n1482 VSUBS 0.018072f
C2145 AVSS.n1484 VSUBS 0.013197f
C2146 AVSS.n1485 VSUBS 0.013464f
C2147 AVSS.n1486 VSUBS 0.257281f
C2148 AVSS.n1487 VSUBS 0.013464f
C2149 AVSS.n1488 VSUBS 0.013197f
C2150 AVSS.n1489 VSUBS 0.013464f
C2151 AVSS.n1490 VSUBS 0.013197f
C2152 AVSS.n1491 VSUBS 0.257281f
C2153 AVSS.n1492 VSUBS 0.013464f
C2154 AVSS.n1493 VSUBS 0.013197f
C2155 AVSS.n1494 VSUBS 0.013197f
C2156 AVSS.n1495 VSUBS 0.013464f
C2157 AVSS.n1496 VSUBS 0.013464f
C2158 AVSS.n1497 VSUBS 0.013197f
C2159 AVSS.n1498 VSUBS 0.013197f
C2160 AVSS.n1499 VSUBS 0.013464f
C2161 AVSS.n1500 VSUBS 0.013464f
C2162 AVSS.n1501 VSUBS 0.013197f
C2163 AVSS.n1502 VSUBS 0.013197f
C2164 AVSS.n1503 VSUBS 0.013464f
C2165 AVSS.n1504 VSUBS 0.013464f
C2166 AVSS.n1505 VSUBS 0.013197f
C2167 AVSS.n1506 VSUBS 0.013197f
C2168 AVSS.n1507 VSUBS 0.013464f
C2169 AVSS.n1508 VSUBS 0.013464f
C2170 AVSS.n1509 VSUBS 0.013197f
C2171 AVSS.n1510 VSUBS 0.013464f
C2172 AVSS.n1511 VSUBS 0.013197f
C2173 AVSS.n1512 VSUBS 0.018889f
C2174 AVSS.n1513 VSUBS 0.020848f
C2175 AVSS.n1514 VSUBS 0.021194f
C2176 AVSS.n1515 VSUBS 0.410221f
C2177 AVSS.n1516 VSUBS 0.257281f
C2178 AVSS.n1517 VSUBS 0.013464f
C2179 AVSS.n1518 VSUBS 0.013197f
C2180 AVSS.n1519 VSUBS 0.013197f
C2181 AVSS.n1520 VSUBS 0.013197f
C2182 AVSS.n1521 VSUBS 0.013464f
C2183 AVSS.n1522 VSUBS 0.257281f
C2184 AVSS.n1523 VSUBS 0.257281f
C2185 AVSS.n1524 VSUBS 0.19582f
C2186 AVSS.n1525 VSUBS 0.013464f
C2187 AVSS.n1526 VSUBS 0.013464f
C2188 AVSS.n1527 VSUBS 0.190102f
C2189 AVSS.n1528 VSUBS 0.257281f
C2190 AVSS.n1529 VSUBS 0.013464f
C2191 AVSS.n1530 VSUBS 0.013197f
C2192 AVSS.n1531 VSUBS 0.013197f
C2193 AVSS.n1532 VSUBS 0.013197f
C2194 AVSS.n1533 VSUBS 0.013464f
C2195 AVSS.n1534 VSUBS 0.257281f
C2196 AVSS.n1535 VSUBS 0.257281f
C2197 AVSS.n1536 VSUBS 0.415938f
C2198 AVSS.n1537 VSUBS 0.021345f
C2199 AVSS.n1538 VSUBS 0.021004f
C2200 AVSS.n1539 VSUBS 0.01932f
C2201 AVSS.n1540 VSUBS 0.013464f
C2202 AVSS.n1541 VSUBS 0.013197f
C2203 AVSS.n1542 VSUBS 0.013197f
C2204 AVSS.n1543 VSUBS 0.013464f
C2205 AVSS.n1544 VSUBS 0.013464f
C2206 AVSS.n1545 VSUBS 0.013197f
C2207 AVSS.n1546 VSUBS 0.013197f
C2208 AVSS.n1547 VSUBS 0.013464f
C2209 AVSS.n1548 VSUBS 0.013464f
C2210 AVSS.n1549 VSUBS 0.013197f
C2211 AVSS.n1550 VSUBS 0.013197f
C2212 AVSS.n1551 VSUBS 0.013464f
C2213 AVSS.n1552 VSUBS 0.013464f
C2214 AVSS.n1553 VSUBS 0.013197f
C2215 AVSS.n1554 VSUBS 0.013197f
C2216 AVSS.n1555 VSUBS 0.013464f
C2217 AVSS.n1556 VSUBS 0.013464f
C2218 AVSS.n1557 VSUBS 0.013197f
C2219 AVSS.n1558 VSUBS 0.010705f
C2220 AVSS.n1559 VSUBS 0.013464f
C2221 AVSS.n1560 VSUBS 0.013464f
C2222 AVSS.n1562 VSUBS 0.017108f
C2223 AVSS.n1563 VSUBS 0.017327f
C2224 AVSS.n1565 VSUBS 0.014835f
C2225 AVSS.n1566 VSUBS 0.014713f
C2226 AVSS.n1567 VSUBS 0.013197f
C2227 AVSS.n1568 VSUBS 0.013197f
C2228 AVSS.n1569 VSUBS 0.013464f
C2229 AVSS.n1571 VSUBS 0.013464f
C2230 AVSS.n1573 VSUBS 0.013464f
C2231 AVSS.n1574 VSUBS 0.013197f
C2232 AVSS.n1575 VSUBS 0.013197f
C2233 AVSS.n1577 VSUBS 0.013464f
C2234 AVSS.n1579 VSUBS 0.013464f
C2235 AVSS.n1581 VSUBS 0.013464f
C2236 AVSS.n1582 VSUBS 0.013197f
C2237 AVSS.n1583 VSUBS 0.013197f
C2238 AVSS.n1584 VSUBS 0.013197f
C2239 AVSS.n1585 VSUBS 0.013464f
C2240 AVSS.n1587 VSUBS 0.014676f
C2241 AVSS.n1588 VSUBS 0.016888f
C2242 AVSS.n1589 VSUBS 0.016685f
C2243 AVSS.n1590 VSUBS 0.013464f
C2244 AVSS.n1591 VSUBS 0.013464f
C2245 AVSS.n1594 VSUBS 0.018072f
C2246 AVSS.n1595 VSUBS 0.088342f
C2247 AVSS.n1597 VSUBS 0.077272f
C2248 AVSS.n1598 VSUBS 0.030324f
C2249 AVSS.n1599 VSUBS 0.067428f
C2250 AVSS.n1600 VSUBS 0.046257f
C2251 AVSS.n1601 VSUBS 0.051397f
C2252 AVSS.n1602 VSUBS 0.205976f
C2253 AVSS.n1603 VSUBS 0.084482f
C2254 AVSS.n1604 VSUBS 0.0905f
C2255 AVSS.n1605 VSUBS 0.0905f
C2256 AVSS.n1607 VSUBS 0.0905f
C2257 AVSS.n1609 VSUBS 0.0905f
C2258 AVSS.n1610 VSUBS 0.114219f
C2259 AVSS.n1612 VSUBS 0.051397f
C2260 AVSS.n1613 VSUBS 0.045828f
C2261 AVSS.n1614 VSUBS 0.04266f
C2262 AVSS.n1615 VSUBS 0.205814f
C2263 AVSS.n1616 VSUBS 0.093787f
C2264 AVSS.n1617 VSUBS 0.165515f
C2265 AVSS.n1619 VSUBS 0.143448f
C2266 AVSS.n1620 VSUBS 0.160158f
C2267 AVSS.n1621 VSUBS 0.131596f
C2268 AVSS.n1622 VSUBS 0.114219f
C2269 AVSS.n1623 VSUBS 0.018072f
C2270 AVSS.n1624 VSUBS 0.017703f
C2271 AVSS.n1627 VSUBS 0.013002f
C2272 AVSS.t113 VSUBS 1.58362f
C2273 AVSS.n1631 VSUBS 0.014231f
C2274 AVSS.n1636 VSUBS 0.015863f
C2275 AVSS.n1660 VSUBS 0.013536f
C2276 AVSS.n1661 VSUBS 0.013536f
C2277 AVSS.n1662 VSUBS 0.014085f
C2278 AVSS.n1663 VSUBS 0.014085f
C2279 AVSS.n1677 VSUBS 0.014104f
C2280 AVSS.n1678 VSUBS 0.014104f
C2281 AVSS.n1680 VSUBS 0.015863f
C2282 AVSS.n1695 VSUBS 0.015203f
C2283 AVSS.n1696 VSUBS 0.015203f
C2284 AVSS.n1697 VSUBS 0.014231f
C2285 AVSS.n1712 VSUBS 0.010886f
C2286 AVSS.n1715 VSUBS 0.024671f
C2287 AVSS.n1716 VSUBS 0.010705f
C2288 AVSS.n1717 VSUBS 0.017108f
C2289 AVSS.n1718 VSUBS 0.013464f
C2290 AVSS.n1719 VSUBS 0.863324f
C2291 AVSS.n1722 VSUBS 0.092461f
C2292 AVSS.n1723 VSUBS 0.017925f
C2293 AVSS.n1724 VSUBS 0.013197f
C2294 AVSS.n1725 VSUBS 0.013464f
C2295 AVSS.n1726 VSUBS 0.135542f
C2296 AVSS.n1727 VSUBS 0.013464f
C2297 AVSS.n1728 VSUBS 0.013197f
C2298 AVSS.n1730 VSUBS 0.013464f
C2299 AVSS.n1731 VSUBS 0.013197f
C2300 AVSS.n1733 VSUBS 0.013464f
C2301 AVSS.n1734 VSUBS 0.013197f
C2302 AVSS.n1736 VSUBS 0.014835f
C2303 AVSS.n1738 VSUBS 0.138076f
C2304 AVSS.n1739 VSUBS 0.010705f
C2305 AVSS.n1741 VSUBS 0.013464f
C2306 AVSS.n1746 VSUBS 0.013464f
C2307 AVSS.n1747 VSUBS 0.011633f
C2308 AVSS.n1748 VSUBS 0.025381f
C2309 AVSS.n1749 VSUBS 0.138021f
C2310 AVSS.n1753 VSUBS 0.013002f
C2311 AVSS.n1770 VSUBS 0.015203f
C2312 AVSS.n1784 VSUBS 0.014231f
C2313 AVSS.n1786 VSUBS 0.011838f
C2314 AVSS.n1788 VSUBS 0.010931f
C2315 AVSS.n1804 VSUBS 0.013536f
C2316 AVSS.n1805 VSUBS 0.014085f
C2317 AVSS.n1821 VSUBS 0.014104f
C2318 AVSS.n1822 VSUBS 0.010825f
C2319 AVSS.n1823 VSUBS 0.025381f
C2320 AVSS.n1825 VSUBS 0.013464f
C2321 AVSS.n1826 VSUBS 0.013464f
C2322 AVSS.n1827 VSUBS 0.013197f
C2323 AVSS.n1828 VSUBS 0.013197f
C2324 AVSS.n1829 VSUBS 0.013464f
C2325 AVSS.n1830 VSUBS 0.013464f
C2326 AVSS.n1831 VSUBS 0.013197f
C2327 AVSS.n1832 VSUBS 0.013197f
C2328 AVSS.n1833 VSUBS 0.013464f
C2329 AVSS.n1834 VSUBS 0.013464f
C2330 AVSS.n1835 VSUBS 0.013197f
C2331 AVSS.n1836 VSUBS 0.013197f
C2332 AVSS.n1837 VSUBS 0.013464f
C2333 AVSS.n1838 VSUBS 0.013464f
C2334 AVSS.n1839 VSUBS 0.013197f
C2335 AVSS.n1840 VSUBS 0.013197f
C2336 AVSS.n1841 VSUBS 0.013464f
C2337 AVSS.n1842 VSUBS 0.013464f
C2338 AVSS.n1845 VSUBS 0.017129f
C2339 AVSS.n1846 VSUBS 0.019048f
C2340 AVSS.n1847 VSUBS 0.135542f
C2341 AVSS.n1848 VSUBS 0.013197f
C2342 AVSS.n1849 VSUBS 0.013464f
C2343 AVSS.n1850 VSUBS 0.013197f
C2344 AVSS.n1851 VSUBS 0.013464f
C2345 AVSS.n1853 VSUBS 0.019496f
C2346 AVSS.n1854 VSUBS 0.013197f
C2347 AVSS.n1855 VSUBS 0.013464f
C2348 AVSS.n1856 VSUBS 0.013197f
C2349 AVSS.n1857 VSUBS 0.013464f
C2350 AVSS.n1858 VSUBS 0.010705f
C2351 AVSS.n1859 VSUBS 0.014835f
C2352 AVSS.n1860 VSUBS 0.017327f
C2353 AVSS.n1862 VSUBS 0.017108f
C2354 AVSS.n1864 VSUBS 0.013464f
C2355 AVSS.n1866 VSUBS 0.013464f
C2356 AVSS.n1868 VSUBS 0.013464f
C2357 AVSS.n1869 VSUBS 0.013197f
C2358 AVSS.n1870 VSUBS 0.013197f
C2359 AVSS.n1871 VSUBS 0.013197f
C2360 AVSS.n1872 VSUBS 0.013464f
C2361 AVSS.n1874 VSUBS 0.013464f
C2362 AVSS.n1876 VSUBS 0.013464f
C2363 AVSS.n1877 VSUBS 0.013197f
C2364 AVSS.n1878 VSUBS 0.013197f
C2365 AVSS.n1879 VSUBS 0.013197f
C2366 AVSS.n1880 VSUBS 0.013464f
C2367 AVSS.n1882 VSUBS 0.013464f
C2368 AVSS.n1884 VSUBS 0.013464f
C2369 AVSS.n1889 VSUBS 0.013536f
C2370 AVSS.n1893 VSUBS 0.010886f
C2371 AVSS.n1908 VSUBS 0.015863f
C2372 AVSS.n1923 VSUBS 0.013002f
C2373 AVSS.n1924 VSUBS 0.013002f
C2374 AVSS.n1925 VSUBS 0.010886f
C2375 AVSS.n1939 VSUBS 0.014231f
C2376 AVSS.n1940 VSUBS 0.014231f
C2377 AVSS.n1941 VSUBS 0.015203f
C2378 AVSS.n1942 VSUBS 0.015203f
C2379 AVSS.n1957 VSUBS 0.015863f
C2380 AVSS.n1969 VSUBS 0.014104f
C2381 AVSS.n1970 VSUBS 0.014104f
C2382 AVSS.t81 VSUBS 1.58362f
C2383 AVSS.n1973 VSUBS 0.014085f
C2384 AVSS.n1975 VSUBS 0.010931f
C2385 AVSS.n1976 VSUBS 0.073941f
C2386 AVSS.n1980 VSUBS 0.013002f
C2387 AVSS.n1999 VSUBS 0.015863f
C2388 AVSS.n2011 VSUBS 0.014231f
C2389 AVSS.n2012 VSUBS 0.014231f
C2390 AVSS.n2013 VSUBS 0.015203f
C2391 AVSS.n2014 VSUBS 0.015203f
C2392 AVSS.n2029 VSUBS 0.015863f
C2393 AVSS.n2044 VSUBS 0.013536f
C2394 AVSS.n2046 VSUBS 0.010931f
C2395 AVSS.n2048 VSUBS 0.014085f
C2396 AVSS.n2062 VSUBS 0.014104f
C2397 AVSS.n2063 VSUBS 0.014104f
C2398 AVSS.t77 VSUBS 1.58362f
C2399 AVSS.n2065 VSUBS 0.010886f
C2400 AVSS.n2068 VSUBS 0.073869f
C2401 AVSS.n2069 VSUBS 0.010705f
C2402 AVSS.n2070 VSUBS 0.017108f
C2403 AVSS.n2071 VSUBS 0.013464f
C2404 AVSS.n2072 VSUBS 0.014713f
C2405 AVSS.n2073 VSUBS 0.135542f
C2406 AVSS.n2074 VSUBS 0.013464f
C2407 AVSS.n2075 VSUBS 0.013197f
C2408 AVSS.n2077 VSUBS 0.013464f
C2409 AVSS.n2078 VSUBS 0.013197f
C2410 AVSS.n2080 VSUBS 0.013464f
C2411 AVSS.n2082 VSUBS 0.013197f
C2412 AVSS.n2083 VSUBS 0.135542f
C2413 AVSS.n2084 VSUBS 0.013197f
C2414 AVSS.n2085 VSUBS 0.013464f
C2415 AVSS.n2086 VSUBS 0.013197f
C2416 AVSS.n2087 VSUBS 0.013464f
C2417 AVSS.n2088 VSUBS 0.013197f
C2418 AVSS.n2089 VSUBS 0.019496f
C2419 AVSS.n2090 VSUBS 0.013197f
C2420 AVSS.n2091 VSUBS 0.013197f
C2421 AVSS.n2092 VSUBS 0.013464f
C2422 AVSS.n2093 VSUBS 0.013197f
C2423 AVSS.n2096 VSUBS 0.013464f
C2424 AVSS.n2097 VSUBS 0.013197f
C2425 AVSS.n2098 VSUBS 0.013197f
C2426 AVSS.n2099 VSUBS 0.013464f
C2427 AVSS.n2101 VSUBS 0.013464f
C2428 AVSS.n2102 VSUBS 0.013464f
C2429 AVSS.n2103 VSUBS 0.013197f
C2430 AVSS.n2104 VSUBS 0.013197f
C2431 AVSS.n2105 VSUBS 0.013197f
C2432 AVSS.n2106 VSUBS 0.013464f
C2433 AVSS.n2108 VSUBS 0.013464f
C2434 AVSS.n2109 VSUBS 0.013464f
C2435 AVSS.n2111 VSUBS 0.013464f
C2436 AVSS.n2112 VSUBS 0.013197f
C2437 AVSS.n2113 VSUBS 0.01932f
C2438 AVSS.n2114 VSUBS 0.021004f
C2439 AVSS.n2115 VSUBS 0.021345f
C2440 AVSS.n2117 VSUBS 0.013464f
C2441 AVSS.n2119 VSUBS 0.013464f
C2442 AVSS.n2120 VSUBS 0.013197f
C2443 AVSS.n2121 VSUBS 0.013197f
C2444 AVSS.n2122 VSUBS 0.013197f
C2445 AVSS.n2123 VSUBS 0.013464f
C2446 AVSS.n2125 VSUBS 0.013464f
C2447 AVSS.n2127 VSUBS 0.013464f
C2448 AVSS.n2128 VSUBS 0.013197f
C2449 AVSS.n2129 VSUBS 0.013197f
C2450 AVSS.n2130 VSUBS 0.013197f
C2451 AVSS.n2131 VSUBS 0.013464f
C2452 AVSS.n2133 VSUBS 0.013464f
C2453 AVSS.n2134 VSUBS 0.013464f
C2454 AVSS.n2136 VSUBS 0.021194f
C2455 AVSS.n2137 VSUBS 0.020848f
C2456 AVSS.n2138 VSUBS 0.018889f
C2457 AVSS.n2139 VSUBS 0.013464f
C2458 AVSS.n2140 VSUBS 0.013197f
C2459 AVSS.n2141 VSUBS 0.013197f
C2460 AVSS.n2142 VSUBS 0.013464f
C2461 AVSS.n2143 VSUBS 0.013464f
C2462 AVSS.n2144 VSUBS 0.013197f
C2463 AVSS.n2145 VSUBS 0.013197f
C2464 AVSS.n2146 VSUBS 0.013464f
C2465 AVSS.n2147 VSUBS 0.013464f
C2466 AVSS.n2148 VSUBS 0.013197f
C2467 AVSS.n2149 VSUBS 0.013197f
C2468 AVSS.n2150 VSUBS 0.013464f
C2469 AVSS.n2151 VSUBS 0.013464f
C2470 AVSS.n2152 VSUBS 0.013197f
C2471 AVSS.n2153 VSUBS 0.013197f
C2472 AVSS.n2154 VSUBS 0.013464f
C2473 AVSS.n2155 VSUBS 0.013464f
C2474 AVSS.n2156 VSUBS 0.013197f
C2475 AVSS.n2157 VSUBS 0.010705f
C2476 AVSS.n2158 VSUBS 0.013464f
C2477 AVSS.n2159 VSUBS 0.013464f
C2478 AVSS.n2161 VSUBS 0.016685f
C2479 AVSS.n2163 VSUBS 0.016888f
C2480 AVSS.n2164 VSUBS 0.014676f
C2481 AVSS.n2165 VSUBS 0.014549f
C2482 AVSS.n2166 VSUBS 0.013197f
C2483 AVSS.n2167 VSUBS 0.013197f
C2484 AVSS.n2168 VSUBS 0.013464f
C2485 AVSS.n2170 VSUBS 0.013464f
C2486 AVSS.n2171 VSUBS 0.013464f
C2487 AVSS.n2172 VSUBS 0.012464f
C2488 AVSS.n2174 VSUBS 0.013197f
C2489 AVSS.n2175 VSUBS 0.013464f
C2490 AVSS.n2177 VSUBS 0.013464f
C2491 AVSS.n2178 VSUBS 0.013464f
C2492 AVSS.n2179 VSUBS 0.013197f
C2493 AVSS.n2180 VSUBS 0.013197f
C2494 AVSS.n2181 VSUBS 0.013197f
C2495 AVSS.n2182 VSUBS 0.013464f
C2496 AVSS.n2184 VSUBS 0.014835f
C2497 AVSS.n2185 VSUBS 0.017327f
C2498 AVSS.n2187 VSUBS 0.013464f
C2499 AVSS.n2190 VSUBS 0.017703f
C2500 AVSS.n2191 VSUBS 0.068602f
C2501 AVSS.n2192 VSUBS 0.01429f
C2502 AVSS.n2193 VSUBS 0.024742f
C2503 AVSS.n2194 VSUBS 0.024813f
C2504 AVSS.n2195 VSUBS 0.024742f
C2505 AVSS.n2196 VSUBS 0.013197f
C2506 AVSS.n2197 VSUBS 0.013464f
C2507 AVSS.n2198 VSUBS 0.013197f
C2508 AVSS.n2199 VSUBS 0.013464f
C2509 AVSS.n2200 VSUBS 0.013197f
C2510 AVSS.n2201 VSUBS 0.014713f
C2511 AVSS.n2202 VSUBS 0.013464f
C2512 AVSS.n2203 VSUBS 0.013197f
C2513 AVSS.n2205 VSUBS 0.013464f
C2514 AVSS.n2206 VSUBS 0.013197f
C2515 AVSS.n2208 VSUBS 0.013464f
C2516 AVSS.n2209 VSUBS 0.013197f
C2517 AVSS.n2210 VSUBS 0.013464f
C2518 AVSS.n2211 VSUBS 0.013464f
C2519 AVSS.n2212 VSUBS 0.013197f
C2520 AVSS.n2213 VSUBS 0.013197f
C2521 AVSS.n2214 VSUBS 0.013464f
C2522 AVSS.n2215 VSUBS 0.013464f
C2523 AVSS.n2216 VSUBS 0.013197f
C2524 AVSS.n2217 VSUBS 0.013197f
C2525 AVSS.n2218 VSUBS 0.013464f
C2526 AVSS.n2219 VSUBS 0.013464f
C2527 AVSS.n2220 VSUBS 0.013197f
C2528 AVSS.n2221 VSUBS 0.013197f
C2529 AVSS.n2222 VSUBS 0.013464f
C2530 AVSS.n2223 VSUBS 0.013464f
C2531 AVSS.n2224 VSUBS 0.013197f
C2532 AVSS.n2225 VSUBS 0.013197f
C2533 AVSS.n2226 VSUBS 0.013464f
C2534 AVSS.n2227 VSUBS 0.013464f
C2535 AVSS.n2228 VSUBS 0.013197f
C2536 AVSS.n2229 VSUBS 0.016685f
C2537 AVSS.n2231 VSUBS 0.016888f
C2538 AVSS.n2232 VSUBS 0.014676f
C2539 AVSS.n2233 VSUBS 0.014549f
C2540 AVSS.n2234 VSUBS 0.013197f
C2541 AVSS.n2235 VSUBS 0.013197f
C2542 AVSS.n2236 VSUBS 0.013464f
C2543 AVSS.n2238 VSUBS 0.013464f
C2544 AVSS.n2239 VSUBS 0.013464f
C2545 AVSS.n2240 VSUBS 0.012464f
C2546 AVSS.n2242 VSUBS 0.013197f
C2547 AVSS.n2243 VSUBS 0.013464f
C2548 AVSS.n2245 VSUBS 0.013464f
C2549 AVSS.n2246 VSUBS 0.013464f
C2550 AVSS.n2247 VSUBS 0.013197f
C2551 AVSS.n2248 VSUBS 0.013197f
C2552 AVSS.n2249 VSUBS 0.013197f
C2553 AVSS.n2250 VSUBS 0.013464f
C2554 AVSS.n2252 VSUBS 0.014835f
C2555 AVSS.n2253 VSUBS 0.017327f
C2556 AVSS.n2254 VSUBS 0.017108f
C2557 AVSS.n2255 VSUBS 0.013197f
C2558 AVSS.n2256 VSUBS 0.013464f
C2559 AVSS.n2257 VSUBS 0.013464f
C2560 AVSS.n2258 VSUBS 0.013197f
C2561 AVSS.n2259 VSUBS 0.013197f
C2562 AVSS.n2260 VSUBS 0.013464f
C2563 AVSS.n2261 VSUBS 0.013464f
C2564 AVSS.n2262 VSUBS 0.013197f
C2565 AVSS.n2263 VSUBS 0.013197f
C2566 AVSS.n2264 VSUBS 0.013464f
C2567 AVSS.n2265 VSUBS 0.013464f
C2568 AVSS.n2266 VSUBS 0.013197f
C2569 AVSS.n2267 VSUBS 0.013197f
C2570 AVSS.n2268 VSUBS 0.013464f
C2571 AVSS.n2269 VSUBS 0.013464f
C2572 AVSS.n2270 VSUBS 0.013197f
C2573 AVSS.n2271 VSUBS 0.013197f
C2574 AVSS.n2272 VSUBS 0.013464f
C2575 AVSS.n2273 VSUBS 0.013464f
C2576 AVSS.n2274 VSUBS 0.013197f
C2577 AVSS.n2275 VSUBS 0.013464f
C2578 AVSS.n2276 VSUBS 0.013197f
C2579 AVSS.n2277 VSUBS 0.01932f
C2580 AVSS.n2278 VSUBS 0.021004f
C2581 AVSS.n2279 VSUBS 0.021345f
C2582 AVSS.n2281 VSUBS 0.013464f
C2583 AVSS.n2283 VSUBS 0.013464f
C2584 AVSS.n2284 VSUBS 0.013197f
C2585 AVSS.n2285 VSUBS 0.013197f
C2586 AVSS.n2286 VSUBS 0.013197f
C2587 AVSS.n2287 VSUBS 0.013464f
C2588 AVSS.n2289 VSUBS 0.013464f
C2589 AVSS.n2291 VSUBS 0.013464f
C2590 AVSS.n2292 VSUBS 0.013197f
C2591 AVSS.n2293 VSUBS 0.013197f
C2592 AVSS.n2294 VSUBS 0.013197f
C2593 AVSS.n2295 VSUBS 0.013464f
C2594 AVSS.n2297 VSUBS 0.013464f
C2595 AVSS.n2299 VSUBS 0.013464f
C2596 AVSS.n2302 VSUBS 0.024742f
C2597 AVSS.n2304 VSUBS 0.016685f
C2598 AVSS.n2306 VSUBS 0.012464f
C2599 AVSS.n2307 VSUBS 0.013464f
C2600 AVSS.n2308 VSUBS 0.013197f
C2601 AVSS.n2309 VSUBS 0.013464f
C2602 AVSS.n2310 VSUBS 0.013197f
C2603 AVSS.n2312 VSUBS 0.013197f
C2604 AVSS.n2313 VSUBS 0.013464f
C2605 AVSS.n2314 VSUBS 0.013197f
C2606 AVSS.n2315 VSUBS 0.013464f
C2607 AVSS.n2316 VSUBS 0.013197f
C2608 AVSS.n2317 VSUBS 0.013464f
C2609 AVSS.n2318 VSUBS 0.013464f
C2610 AVSS.n2319 VSUBS 0.013197f
C2611 AVSS.n2320 VSUBS 0.013197f
C2612 AVSS.n2321 VSUBS 0.013464f
C2613 AVSS.n2322 VSUBS 0.013464f
C2614 AVSS.n2323 VSUBS 0.013197f
C2615 AVSS.n2324 VSUBS 0.013197f
C2616 AVSS.n2325 VSUBS 0.013464f
C2617 AVSS.n2326 VSUBS 0.013464f
C2618 AVSS.n2327 VSUBS 0.013197f
C2619 AVSS.n2328 VSUBS 0.013197f
C2620 AVSS.n2329 VSUBS 0.013464f
C2621 AVSS.n2330 VSUBS 0.013464f
C2622 AVSS.n2331 VSUBS 0.013197f
C2623 AVSS.n2332 VSUBS 0.013197f
C2624 AVSS.n2333 VSUBS 0.013464f
C2625 AVSS.n2334 VSUBS 0.013464f
C2626 AVSS.n2335 VSUBS 0.013197f
C2627 AVSS.n2336 VSUBS 0.013464f
C2628 AVSS.n2337 VSUBS 0.013197f
C2629 AVSS.n2338 VSUBS 0.018889f
C2630 AVSS.n2340 VSUBS 0.021194f
C2631 AVSS.n2341 VSUBS 0.018062f
C2632 AVSS.n2344 VSUBS 0.013197f
C2633 AVSS.n2345 VSUBS 0.013464f
C2634 AVSS.n2347 VSUBS 0.013464f
C2635 AVSS.n2349 VSUBS 0.013464f
C2636 AVSS.n2350 VSUBS 0.013197f
C2637 AVSS.n2351 VSUBS 0.013197f
C2638 AVSS.n2352 VSUBS 0.013197f
C2639 AVSS.n2353 VSUBS 0.013464f
C2640 AVSS.n2355 VSUBS 0.013464f
C2641 AVSS.n2356 VSUBS 0.013464f
C2642 AVSS.n2357 VSUBS 0.013197f
C2643 AVSS.n2358 VSUBS 0.013197f
C2644 AVSS.n2359 VSUBS 0.013464f
C2645 AVSS.n2360 VSUBS 0.013464f
C2646 AVSS.n2362 VSUBS 0.021345f
C2647 AVSS.n2363 VSUBS 0.021004f
C2648 AVSS.n2364 VSUBS 0.01932f
C2649 AVSS.n2365 VSUBS 0.013464f
C2650 AVSS.n2366 VSUBS 0.013197f
C2651 AVSS.n2367 VSUBS 0.013197f
C2652 AVSS.n2368 VSUBS 0.013464f
C2653 AVSS.n2369 VSUBS 0.013464f
C2654 AVSS.n2370 VSUBS 0.013197f
C2655 AVSS.n2371 VSUBS 0.013197f
C2656 AVSS.n2372 VSUBS 0.013464f
C2657 AVSS.n2373 VSUBS 0.013464f
C2658 AVSS.n2374 VSUBS 0.013197f
C2659 AVSS.n2375 VSUBS 0.013197f
C2660 AVSS.n2376 VSUBS 0.013464f
C2661 AVSS.n2377 VSUBS 0.013464f
C2662 AVSS.n2378 VSUBS 0.013197f
C2663 AVSS.n2379 VSUBS 0.013197f
C2664 AVSS.n2380 VSUBS 0.013464f
C2665 AVSS.n2381 VSUBS 0.013464f
C2666 AVSS.n2382 VSUBS 0.013197f
C2667 AVSS.n2383 VSUBS 0.013197f
C2668 AVSS.n2384 VSUBS 0.013464f
C2669 AVSS.n2385 VSUBS 0.013464f
C2670 AVSS.n2386 VSUBS 0.013197f
C2671 AVSS.n2387 VSUBS 0.017108f
C2672 AVSS.n2388 VSUBS 0.017327f
C2673 AVSS.n2390 VSUBS 0.014835f
C2674 AVSS.n2391 VSUBS 0.014713f
C2675 AVSS.n2392 VSUBS 0.013197f
C2676 AVSS.n2393 VSUBS 0.013197f
C2677 AVSS.n2394 VSUBS 0.013464f
C2678 AVSS.n2396 VSUBS 0.013464f
C2679 AVSS.n2398 VSUBS 0.013464f
C2680 AVSS.n2399 VSUBS 0.013197f
C2681 AVSS.n2400 VSUBS 0.013197f
C2682 AVSS.n2402 VSUBS 0.013464f
C2683 AVSS.n2404 VSUBS 0.013464f
C2684 AVSS.n2405 VSUBS 0.013464f
C2685 AVSS.n2406 VSUBS 0.013197f
C2686 AVSS.n2407 VSUBS 0.013197f
C2687 AVSS.n2408 VSUBS 0.013464f
C2688 AVSS.n2409 VSUBS 0.013464f
C2689 AVSS.n2411 VSUBS 0.016888f
C2690 AVSS.n2412 VSUBS 0.014676f
C2691 AVSS.n2413 VSUBS 0.011763f
C2692 AVSS.n2415 VSUBS 0.024813f
C2693 AVSS.n2416 VSUBS 0.092666f
C2694 AVSS.t114 VSUBS 1.58362f
C2695 AVSS.n2424 VSUBS 0.014231f
C2696 AVSS.n2428 VSUBS 0.010886f
C2697 AVSS.n2435 VSUBS 0.014085f
C2698 AVSS.n2453 VSUBS 0.010931f
C2699 AVSS.n2455 VSUBS 0.013536f
C2700 AVSS.n2468 VSUBS 0.013002f
C2701 AVSS.n2469 VSUBS 0.013002f
C2702 AVSS.n2471 VSUBS 0.010886f
C2703 AVSS.n2487 VSUBS 0.014231f
C2704 AVSS.n2489 VSUBS 0.015203f
C2705 AVSS.n2490 VSUBS 0.015203f
C2706 AVSS.n2504 VSUBS 0.015863f
C2707 AVSS.n2506 VSUBS 0.014104f
C2708 AVSS.n2507 VSUBS 0.010825f
C2709 AVSS.n2508 VSUBS 0.012104f
C2710 AVSS.n2509 VSUBS 0.092595f
C2711 AVSS.n2510 VSUBS 0.025381f
C2712 AVSS.n2512 VSUBS 0.01756f
C2713 AVSS.n2514 VSUBS 0.017925f
C2714 AVSS.n2515 VSUBS 0.021345f
C2715 AVSS.n2517 VSUBS 0.013464f
C2716 AVSS.n2519 VSUBS 0.013464f
C2717 AVSS.n2520 VSUBS 0.013197f
C2718 AVSS.n2521 VSUBS 0.013197f
C2719 AVSS.n2522 VSUBS 0.013197f
C2720 AVSS.n2523 VSUBS 0.013464f
C2721 AVSS.n2525 VSUBS 0.013464f
C2722 AVSS.n2527 VSUBS 0.013464f
C2723 AVSS.n2528 VSUBS 0.013197f
C2724 AVSS.n2529 VSUBS 0.013197f
C2725 AVSS.n2530 VSUBS 0.013197f
C2726 AVSS.n2531 VSUBS 0.013464f
C2727 AVSS.n2533 VSUBS 0.013464f
C2728 AVSS.n2534 VSUBS 0.013464f
C2729 AVSS.n2536 VSUBS 0.021194f
C2730 AVSS.n2537 VSUBS 0.018062f
C2731 AVSS.n2539 VSUBS 0.138083f
C2732 AVSS.n2540 VSUBS 0.012104f
C2733 AVSS.n2542 VSUBS 0.015863f
C2734 AVSS.t82 VSUBS 1.58362f
C2735 AVSS.n2558 VSUBS 0.010886f
C2736 AVSS.n2561 VSUBS 0.13802f
C2737 AVSS.n2564 VSUBS 0.013464f
C2738 AVSS.n2565 VSUBS 0.013464f
C2739 AVSS.n2566 VSUBS 0.013197f
C2740 AVSS.n2567 VSUBS 0.013197f
C2741 AVSS.n2568 VSUBS 0.013464f
C2742 AVSS.n2569 VSUBS 0.013464f
C2743 AVSS.n2570 VSUBS 0.013197f
C2744 AVSS.n2571 VSUBS 0.013197f
C2745 AVSS.n2572 VSUBS 0.013464f
C2746 AVSS.n2573 VSUBS 0.013464f
C2747 AVSS.n2575 VSUBS 0.013464f
C2748 AVSS.n2576 VSUBS 0.012464f
C2749 AVSS.n2577 VSUBS 0.013197f
C2750 AVSS.n2579 VSUBS 0.013197f
C2751 AVSS.n2580 VSUBS 0.013464f
C2752 AVSS.n2582 VSUBS 0.135542f
C2753 AVSS.n2584 VSUBS 0.014676f
C2754 AVSS.n2585 VSUBS 0.011763f
C2755 AVSS.n2586 VSUBS 0.016685f
C2756 AVSS.n2587 VSUBS 0.013464f
C2757 AVSS.n2590 VSUBS 0.025568f
C2758 AVSS.n2591 VSUBS 0.081912f
C2759 AVSS.n2594 VSUBS 0.013002f
C2760 AVSS.t111 VSUBS 1.58362f
C2761 AVSS.n2598 VSUBS 0.014231f
C2762 AVSS.n2603 VSUBS 0.015863f
C2763 AVSS.n2627 VSUBS 0.013536f
C2764 AVSS.n2628 VSUBS 0.013536f
C2765 AVSS.n2629 VSUBS 0.014085f
C2766 AVSS.n2630 VSUBS 0.014085f
C2767 AVSS.n2644 VSUBS 0.014104f
C2768 AVSS.n2645 VSUBS 0.014104f
C2769 AVSS.n2647 VSUBS 0.015863f
C2770 AVSS.n2662 VSUBS 0.015203f
C2771 AVSS.n2664 VSUBS 0.011838f
C2772 AVSS.n2680 VSUBS 0.010886f
C2773 AVSS.n2683 VSUBS 0.010736f
C2774 AVSS.n2686 VSUBS 0.015203f
C2775 AVSS.n2727 VSUBS 0.010886f
C2776 AVSS.n2728 VSUBS 0.010886f
C2777 AVSS.n2729 VSUBS 0.013002f
C2778 AVSS.n2730 VSUBS 0.013002f
C2779 AVSS.n2745 VSUBS 0.013536f
C2780 AVSS.n2746 VSUBS 0.013536f
C2781 AVSS.n2747 VSUBS 0.014085f
C2782 AVSS.n2748 VSUBS 0.014085f
C2783 AVSS.n2763 VSUBS 0.014104f
C2784 AVSS.n2764 VSUBS 0.014104f
C2785 AVSS.n2765 VSUBS 0.015863f
C2786 AVSS.n2766 VSUBS 0.015863f
C2787 AVSS.t75 VSUBS 1.58362f
C2788 AVSS.n2772 VSUBS 0.014231f
C2789 AVSS.n2774 VSUBS 0.011838f
C2790 AVSS.n2775 VSUBS 0.0246f
C2791 AVSS.n2776 VSUBS 0.017925f
C2792 AVSS.n2777 VSUBS 0.013197f
C2793 AVSS.n2778 VSUBS 0.013464f
C2794 AVSS.n2779 VSUBS 0.135542f
C2795 AVSS.n2780 VSUBS 0.013464f
C2796 AVSS.n2781 VSUBS 0.013197f
C2797 AVSS.n2783 VSUBS 0.013464f
C2798 AVSS.n2784 VSUBS 0.013197f
C2799 AVSS.n2786 VSUBS 0.013464f
C2800 AVSS.n2787 VSUBS 0.013197f
C2801 AVSS.n2789 VSUBS 0.014835f
C2802 AVSS.n2790 VSUBS 0.013197f
C2803 AVSS.n2791 VSUBS 0.013464f
C2804 AVSS.t76 VSUBS 2.06361f
C2805 AVSS.n2797 VSUBS 0.205976f
C2806 AVSS.n2798 VSUBS 0.045828f
C2807 AVSS.n2799 VSUBS 0.135542f
C2808 AVSS.n2800 VSUBS 0.135542f
C2809 AVSS.n2801 VSUBS 0.135542f
C2810 AVSS.n2802 VSUBS 0.135542f
C2811 AVSS.n2807 VSUBS 0.013464f
C2812 AVSS.n2808 VSUBS 0.016888f
C2813 AVSS.n2809 VSUBS 0.013464f
C2814 AVSS.n2810 VSUBS 0.013464f
C2815 AVSS.n2811 VSUBS 0.013197f
C2816 AVSS.n2812 VSUBS 0.013197f
C2817 AVSS.n2813 VSUBS 0.013464f
C2818 AVSS.n2814 VSUBS 0.013464f
C2819 AVSS.n2815 VSUBS 0.013197f
C2820 AVSS.n2816 VSUBS 0.013197f
C2821 AVSS.n2817 VSUBS 0.013464f
C2822 AVSS.n2818 VSUBS 0.013464f
C2823 AVSS.n2820 VSUBS 0.012464f
C2824 AVSS.n2821 VSUBS 0.013464f
C2825 AVSS.n2822 VSUBS 0.013464f
C2826 AVSS.n2823 VSUBS 0.013197f
C2827 AVSS.n2824 VSUBS 0.013464f
C2828 AVSS.n2825 VSUBS 0.013197f
C2829 AVSS.n2826 VSUBS 0.013197f
C2830 AVSS.n2827 VSUBS 0.013197f
C2831 AVSS.n2828 VSUBS 0.013464f
C2832 AVSS.n2829 VSUBS 0.019048f
C2833 AVSS.n2835 VSUBS 0.013464f
C2834 AVSS.n2836 VSUBS 0.014676f
C2835 AVSS.n2837 VSUBS 0.013197f
C2836 AVSS.n2838 VSUBS 0.013197f
C2837 AVSS.n2839 VSUBS 0.013464f
C2838 AVSS.n2840 VSUBS 0.013197f
C2839 AVSS.n2842 VSUBS 0.013464f
C2840 AVSS.n2843 VSUBS 0.013197f
C2841 AVSS.n2844 VSUBS 0.013197f
C2842 AVSS.n2845 VSUBS 0.013464f
C2843 AVSS.n2847 VSUBS 0.013464f
C2844 AVSS.n2849 VSUBS 0.013464f
C2845 AVSS.n2850 VSUBS 0.013197f
C2846 AVSS.n2851 VSUBS 0.013197f
C2847 AVSS.n2852 VSUBS 0.013197f
C2848 AVSS.n2853 VSUBS 0.013464f
C2849 AVSS.n2855 VSUBS 0.013464f
C2850 AVSS.n2856 VSUBS 0.013464f
C2851 AVSS.n2858 VSUBS 0.021194f
C2852 AVSS.n2859 VSUBS 0.020848f
C2853 AVSS.n2860 VSUBS 0.018889f
C2854 AVSS.n2861 VSUBS 0.013464f
C2855 AVSS.n2862 VSUBS 0.013197f
C2856 AVSS.n2863 VSUBS 0.013197f
C2857 AVSS.n2864 VSUBS 0.013464f
C2858 AVSS.n2865 VSUBS 0.013464f
C2859 AVSS.n2866 VSUBS 0.013197f
C2860 AVSS.n2867 VSUBS 0.013197f
C2861 AVSS.n2868 VSUBS 0.013464f
C2862 AVSS.n2869 VSUBS 0.013464f
C2863 AVSS.n2870 VSUBS 0.013197f
C2864 AVSS.n2871 VSUBS 0.013197f
C2865 AVSS.n2872 VSUBS 0.013464f
C2866 AVSS.n2873 VSUBS 0.013464f
C2867 AVSS.n2874 VSUBS 0.013197f
C2868 AVSS.n2875 VSUBS 0.013197f
C2869 AVSS.n2876 VSUBS 0.013464f
C2870 AVSS.n2877 VSUBS 0.013464f
C2871 AVSS.n2878 VSUBS 0.013197f
C2872 AVSS.n2879 VSUBS 0.013464f
C2873 AVSS.n2880 VSUBS 0.013197f
C2874 AVSS.n2881 VSUBS 0.013197f
C2875 AVSS.n2882 VSUBS 0.013197f
C2876 AVSS.n2883 VSUBS 0.013464f
C2877 AVSS.n2884 VSUBS 0.013464f
C2878 AVSS.n2885 VSUBS 0.013197f
C2879 AVSS.n2886 VSUBS 0.013197f
C2880 AVSS.n2887 VSUBS 0.013464f
C2881 AVSS.n2888 VSUBS 0.013464f
C2882 AVSS.n2890 VSUBS 0.012464f
C2883 AVSS.n2891 VSUBS 0.013464f
C2884 AVSS.n2892 VSUBS 0.013464f
C2885 AVSS.n2893 VSUBS 0.013197f
C2886 AVSS.n2894 VSUBS 0.013197f
C2887 AVSS.n2895 VSUBS 0.013464f
C2888 AVSS.n2896 VSUBS 0.013464f
C2889 AVSS.n2897 VSUBS 0.013197f
C2890 AVSS.n2898 VSUBS 0.014549f
C2891 AVSS.n2899 VSUBS 0.016685f
C2892 AVSS.n2900 VSUBS 0.016888f
C2893 AVSS.n2902 VSUBS 0.019048f
C2894 AVSS.n2907 VSUBS 0.013464f
C2895 AVSS.n2908 VSUBS 0.013197f
C2896 AVSS.n2910 VSUBS 0.013197f
C2897 AVSS.n2911 VSUBS 0.013464f
C2898 AVSS.n2912 VSUBS 0.013197f
C2899 AVSS.n2913 VSUBS 0.013464f
C2900 AVSS.n2914 VSUBS 0.01932f
C2901 AVSS.n2915 VSUBS 0.013197f
C2902 AVSS.n2916 VSUBS 0.013464f
C2903 AVSS.n2917 VSUBS 0.013197f
C2904 AVSS.n2919 VSUBS 0.013464f
C2905 AVSS.n2920 VSUBS 0.013197f
C2906 AVSS.n2923 VSUBS 0.013464f
C2907 AVSS.n2924 VSUBS 0.013464f
C2908 AVSS.n2925 VSUBS 0.013197f
C2909 AVSS.n2926 VSUBS 0.013197f
C2910 AVSS.n2927 VSUBS 0.013197f
C2911 AVSS.n2928 VSUBS 0.013464f
C2912 AVSS.n2930 VSUBS 0.013464f
C2913 AVSS.n2931 VSUBS 0.013464f
C2914 AVSS.n2932 VSUBS 0.013197f
C2915 AVSS.n2933 VSUBS 0.013197f
C2916 AVSS.n2934 VSUBS 0.013197f
C2917 AVSS.n2935 VSUBS 0.013464f
C2918 AVSS.n2937 VSUBS 0.013464f
C2919 AVSS.n2938 VSUBS 0.019496f
C2920 AVSS.n2940 VSUBS 0.021345f
C2921 AVSS.n2941 VSUBS 0.021004f
C2922 AVSS.n2942 VSUBS 0.013197f
C2923 AVSS.n2943 VSUBS 0.013197f
C2924 AVSS.n2944 VSUBS 0.013464f
C2925 AVSS.n2946 VSUBS 0.013464f
C2926 AVSS.n2948 VSUBS 0.013464f
C2927 AVSS.n2949 VSUBS 0.013197f
C2928 AVSS.n2950 VSUBS 0.013197f
C2929 AVSS.n2951 VSUBS 0.013197f
C2930 AVSS.n2952 VSUBS 0.013464f
C2931 AVSS.n2954 VSUBS 0.013464f
C2932 AVSS.n2955 VSUBS 0.013464f
C2933 AVSS.n2956 VSUBS 0.013197f
C2934 AVSS.n2957 VSUBS 0.013197f
C2935 AVSS.n2958 VSUBS 0.013464f
C2936 AVSS.n2959 VSUBS 0.013464f
C2937 AVSS.n2961 VSUBS 0.021194f
C2938 AVSS.n2962 VSUBS 0.020848f
C2939 AVSS.n2963 VSUBS 0.018889f
C2940 AVSS.n2964 VSUBS 0.013464f
C2941 AVSS.n2965 VSUBS 0.013197f
C2942 AVSS.n2966 VSUBS 0.013197f
C2943 AVSS.n2967 VSUBS 0.013464f
C2944 AVSS.n2968 VSUBS 0.013464f
C2945 AVSS.n2969 VSUBS 0.013197f
C2946 AVSS.n2970 VSUBS 0.013197f
C2947 AVSS.n2971 VSUBS 0.013464f
C2948 AVSS.n2972 VSUBS 0.013464f
C2949 AVSS.n2973 VSUBS 0.013197f
C2950 AVSS.n2974 VSUBS 0.013197f
C2951 AVSS.n2975 VSUBS 0.013464f
C2952 AVSS.n2976 VSUBS 0.013464f
C2953 AVSS.n2977 VSUBS 0.013197f
C2954 AVSS.n2978 VSUBS 0.013197f
C2955 AVSS.n2979 VSUBS 0.013197f
C2956 AVSS.n2980 VSUBS 0.013464f
C2957 AVSS.n2982 VSUBS 1.57993f
C2958 AVSS.n2989 VSUBS 0.021194f
C2959 AVSS.n2990 VSUBS 0.013464f
C2960 AVSS.n2991 VSUBS 0.013197f
C2961 AVSS.n2992 VSUBS 0.013464f
C2962 AVSS.n2993 VSUBS 0.013197f
C2963 AVSS.n2995 VSUBS 0.013464f
C2964 AVSS.n2996 VSUBS 0.013197f
C2965 AVSS.n2997 VSUBS 0.013197f
C2966 AVSS.n2998 VSUBS 0.013464f
C2967 AVSS.n3000 VSUBS 0.013464f
C2968 AVSS.n3002 VSUBS 0.013464f
C2969 AVSS.n3003 VSUBS 0.013197f
C2970 AVSS.n3004 VSUBS 0.013197f
C2971 AVSS.n3005 VSUBS 0.013197f
C2972 AVSS.n3006 VSUBS 0.013464f
C2973 AVSS.n3008 VSUBS 0.013464f
C2974 AVSS.n3010 VSUBS 0.013464f
C2975 AVSS.n3011 VSUBS 0.013197f
C2976 AVSS.n3012 VSUBS 0.020848f
C2977 AVSS.n3013 VSUBS 0.014549f
C2978 AVSS.n3014 VSUBS 0.013464f
C2979 AVSS.n3015 VSUBS 0.012464f
C2980 AVSS.n3016 VSUBS 0.013464f
C2981 AVSS.n3017 VSUBS 0.013197f
C2982 AVSS.n3019 VSUBS 0.013464f
C2983 AVSS.n3020 VSUBS 0.013197f
C2984 AVSS.n3021 VSUBS 0.013464f
C2985 AVSS.n3023 VSUBS 0.013464f
C2986 AVSS.n3025 VSUBS 0.013464f
C2987 AVSS.n3026 VSUBS 0.013197f
C2988 AVSS.n3027 VSUBS 0.013197f
C2989 AVSS.n3029 VSUBS 0.013464f
C2990 AVSS.n3031 VSUBS 0.013464f
C2991 AVSS.n3033 VSUBS 0.013464f
C2992 AVSS.n3034 VSUBS 0.013197f
C2993 AVSS.n3035 VSUBS 0.013197f
C2994 AVSS.n3036 VSUBS 0.013197f
C2995 AVSS.n3037 VSUBS 0.013464f
C2996 AVSS.n3039 VSUBS 0.014676f
C2997 AVSS.n3040 VSUBS 0.016888f
C2998 AVSS.n3041 VSUBS 0.016685f
C2999 AVSS.n3042 VSUBS 0.013197f
C3000 AVSS.n3043 VSUBS 0.013464f
C3001 AVSS.n3044 VSUBS 0.013464f
C3002 AVSS.n3045 VSUBS 0.013197f
C3003 AVSS.n3046 VSUBS 0.013197f
C3004 AVSS.n3047 VSUBS 0.013464f
C3005 AVSS.n3048 VSUBS 0.013464f
C3006 AVSS.n3049 VSUBS 0.013197f
C3007 AVSS.n3050 VSUBS 0.013197f
C3008 AVSS.n3051 VSUBS 0.013464f
C3009 AVSS.n3052 VSUBS 0.013464f
C3010 AVSS.n3053 VSUBS 0.013197f
C3011 AVSS.n3054 VSUBS 0.013197f
C3012 AVSS.n3055 VSUBS 0.013464f
C3013 AVSS.n3056 VSUBS 0.013464f
C3014 AVSS.n3057 VSUBS 0.013197f
C3015 AVSS.n3058 VSUBS 0.013197f
C3016 AVSS.n3059 VSUBS 0.013464f
C3017 AVSS.n3060 VSUBS 0.013464f
C3018 AVSS.n3061 VSUBS 0.013197f
C3019 AVSS.n3062 VSUBS 0.013197f
C3020 AVSS.n3063 VSUBS 0.018889f
C3021 AVSS.n3064 VSUBS 0.019048f
C3022 AVSS.n3070 VSUBS 0.019048f
C3023 AVSS.n3071 VSUBS 0.013464f
C3024 AVSS.n3073 VSUBS 0.016685f
C3025 AVSS.n3074 VSUBS 0.014676f
C3026 AVSS.n3075 VSUBS 0.027461f
C3027 AVSS.n3076 VSUBS 0.013464f
C3028 AVSS.n3077 VSUBS 0.012464f
C3029 AVSS.n3078 VSUBS 0.013464f
C3030 AVSS.n3079 VSUBS 0.013464f
C3031 AVSS.n3080 VSUBS 0.013197f
C3032 AVSS.n3081 VSUBS 0.013464f
C3033 AVSS.n3082 VSUBS 0.027461f
C3034 AVSS.n3083 VSUBS 0.013464f
C3035 AVSS.n3084 VSUBS 0.017108f
C3036 AVSS.n3086 VSUBS 0.013197f
C3037 AVSS.n3087 VSUBS 0.013464f
C3038 AVSS.n3088 VSUBS 0.013197f
C3039 AVSS.n3089 VSUBS 0.013464f
C3040 AVSS.n3091 VSUBS 0.021345f
C3041 AVSS.n3092 VSUBS 0.013197f
C3042 AVSS.n3093 VSUBS 0.013464f
C3043 AVSS.n3094 VSUBS 0.013197f
C3044 AVSS.n3095 VSUBS 0.013464f
C3045 AVSS.n3096 VSUBS 0.013197f
C3046 AVSS.n3097 VSUBS 0.017129f
C3047 AVSS.n3098 VSUBS 0.020848f
C3048 AVSS.n3099 VSUBS 0.021194f
C3049 AVSS.n3101 VSUBS 0.013464f
C3050 AVSS.n3103 VSUBS 0.013464f
C3051 AVSS.n3104 VSUBS 0.013197f
C3052 AVSS.n3105 VSUBS 0.013197f
C3053 AVSS.n3106 VSUBS 0.013197f
C3054 AVSS.n3107 VSUBS 0.013464f
C3055 AVSS.n3109 VSUBS 0.013464f
C3056 AVSS.n3111 VSUBS 0.013464f
C3057 AVSS.n3112 VSUBS 0.013197f
C3058 AVSS.n3113 VSUBS 0.013197f
C3059 AVSS.n3114 VSUBS 0.013197f
C3060 AVSS.n3115 VSUBS 0.013464f
C3061 AVSS.n3117 VSUBS 0.013464f
C3062 AVSS.n3119 VSUBS 0.013464f
C3063 AVSS.n3120 VSUBS 0.013197f
C3064 AVSS.n3121 VSUBS 0.021004f
C3065 AVSS.n3122 VSUBS 0.075481f
C3066 AVSS.n3125 VSUBS 0.015203f
C3067 AVSS.n3143 VSUBS 0.015863f
C3068 AVSS.n3160 VSUBS 0.012104f
C3069 AVSS.n3173 VSUBS 0.010886f
C3070 AVSS.n3174 VSUBS 0.010886f
C3071 AVSS.n3175 VSUBS 0.013002f
C3072 AVSS.n3176 VSUBS 0.013002f
C3073 AVSS.n3191 VSUBS 0.013536f
C3074 AVSS.n3192 VSUBS 0.013536f
C3075 AVSS.n3193 VSUBS 0.014085f
C3076 AVSS.n3194 VSUBS 0.014085f
C3077 AVSS.n3208 VSUBS 0.010825f
C3078 AVSS.n3209 VSUBS 0.014104f
C3079 AVSS.t100 VSUBS 1.58362f
C3080 AVSS.n3212 VSUBS 0.014231f
C3081 AVSS.n3214 VSUBS 0.011838f
C3082 AVSS.n3215 VSUBS 0.075408f
C3083 AVSS.n3216 VSUBS 0.01633f
C3084 AVSS.n3218 VSUBS 0.01756f
C3085 AVSS.n3219 VSUBS 0.019496f
C3086 AVSS.n3221 VSUBS 0.013464f
C3087 AVSS.n3223 VSUBS 0.013464f
C3088 AVSS.n3224 VSUBS 0.013197f
C3089 AVSS.n3225 VSUBS 0.013197f
C3090 AVSS.n3226 VSUBS 0.013197f
C3091 AVSS.n3227 VSUBS 0.013464f
C3092 AVSS.n3229 VSUBS 0.013464f
C3093 AVSS.n3231 VSUBS 0.013464f
C3094 AVSS.n3232 VSUBS 0.013197f
C3095 AVSS.n3233 VSUBS 0.013197f
C3096 AVSS.n3234 VSUBS 0.013197f
C3097 AVSS.n3235 VSUBS 0.013464f
C3098 AVSS.n3237 VSUBS 0.013464f
C3099 AVSS.n3238 VSUBS 0.013464f
C3100 AVSS.n3239 VSUBS 0.013197f
C3101 AVSS.n3240 VSUBS 0.013197f
C3102 AVSS.n3241 VSUBS 0.013464f
C3103 AVSS.n3242 VSUBS 0.017327f
C3104 AVSS.n3243 VSUBS 0.030665f
C3105 AVSS.n3244 VSUBS 0.029139f
C3106 AVSS.n3245 VSUBS 0.014835f
C3107 AVSS.n3246 VSUBS 0.014713f
C3108 AVSS.n3247 VSUBS 0.013197f
C3109 AVSS.n3248 VSUBS 0.013197f
C3110 AVSS.n3249 VSUBS 0.013464f
C3111 AVSS.n3250 VSUBS 0.027461f
C3112 AVSS.n3251 VSUBS 0.027461f
C3113 AVSS.n3252 VSUBS 0.020291f
C3114 AVSS.n3253 VSUBS 0.027461f
C3115 AVSS.n3254 VSUBS 0.013464f
C3116 AVSS.n3255 VSUBS 0.013197f
C3117 AVSS.n3256 VSUBS 0.013197f
C3118 AVSS.n3258 VSUBS 0.013464f
C3119 AVSS.n3259 VSUBS 0.020901f
C3120 AVSS.n3260 VSUBS 0.027461f
C3121 AVSS.n3261 VSUBS 0.027461f
C3122 AVSS.n3262 VSUBS 0.013464f
C3123 AVSS.n3263 VSUBS 0.013197f
C3124 AVSS.n3264 VSUBS 0.013197f
C3125 AVSS.n3265 VSUBS 0.014549f
C3126 AVSS.n3266 VSUBS 0.013197f
C3127 AVSS.n3267 VSUBS 0.013464f
C3128 AVSS.n3268 VSUBS 0.027461f
C3129 AVSS.n3269 VSUBS 0.028377f
C3130 AVSS.n3270 VSUBS 0.030055f
C3131 AVSS.n3271 VSUBS 0.016888f
C3132 AVSS.n3272 VSUBS 0.013464f
C3133 AVSS.n3273 VSUBS 0.013197f
C3134 AVSS.n3274 VSUBS 0.013197f
C3135 AVSS.n3275 VSUBS 0.013464f
C3136 AVSS.n3276 VSUBS 0.013464f
C3137 AVSS.n3277 VSUBS 0.013197f
C3138 AVSS.n3278 VSUBS 0.013197f
C3139 AVSS.n3279 VSUBS 0.013464f
C3140 AVSS.n3280 VSUBS 0.013464f
C3141 AVSS.n3281 VSUBS 0.013197f
C3142 AVSS.n3282 VSUBS 0.013197f
C3143 AVSS.n3283 VSUBS 0.013464f
C3144 AVSS.n3284 VSUBS 0.013464f
C3145 AVSS.n3285 VSUBS 0.013197f
C3146 AVSS.n3286 VSUBS 0.013197f
C3147 AVSS.n3287 VSUBS 0.013464f
C3148 AVSS.n3288 VSUBS 0.013464f
C3149 AVSS.n3289 VSUBS 0.013197f
C3150 AVSS.n3290 VSUBS 0.013197f
C3151 AVSS.n3292 VSUBS 0.013464f
C3152 AVSS.n3300 VSUBS 0.021194f
C3153 AVSS.n3301 VSUBS 0.013464f
C3154 AVSS.n3302 VSUBS 0.020848f
C3155 AVSS.n3303 VSUBS 0.075408f
C3156 AVSS.n3307 VSUBS 0.013536f
C3157 AVSS.n3311 VSUBS 0.010886f
C3158 AVSS.n3326 VSUBS 0.015863f
C3159 AVSS.n3341 VSUBS 0.013002f
C3160 AVSS.n3358 VSUBS 0.014231f
C3161 AVSS.n3359 VSUBS 0.014231f
C3162 AVSS.n3360 VSUBS 0.015203f
C3163 AVSS.n3361 VSUBS 0.015203f
C3164 AVSS.n3376 VSUBS 0.015863f
C3165 AVSS.n3388 VSUBS 0.014104f
C3166 AVSS.n3389 VSUBS 0.014104f
C3167 AVSS.t97 VSUBS 1.58362f
C3168 AVSS.n3392 VSUBS 0.014085f
C3169 AVSS.n3394 VSUBS 0.010931f
C3170 AVSS.n3395 VSUBS 0.075481f
C3171 AVSS.n3397 VSUBS 0.077272f
C3172 AVSS.n3398 VSUBS 0.030324f
C3173 AVSS.n3399 VSUBS 0.067428f
C3174 AVSS.n3400 VSUBS 0.051397f
C3175 AVSS.n3401 VSUBS 0.051397f
C3176 AVSS.n3402 VSUBS 0.046257f
C3177 AVSS.n3403 VSUBS 0.084482f
C3178 AVSS.n3404 VSUBS 0.0905f
C3179 AVSS.n3405 VSUBS 0.0905f
C3180 AVSS.n3407 VSUBS 0.0905f
C3181 AVSS.n3409 VSUBS 0.0905f
C3182 AVSS.n3411 VSUBS 0.04266f
C3183 AVSS.n3412 VSUBS 0.205814f
C3184 AVSS.n3413 VSUBS 0.093787f
C3185 AVSS.n3414 VSUBS 0.165515f
C3186 AVSS.n3416 VSUBS 0.143448f
C3187 AVSS.n3417 VSUBS 0.160158f
C3188 AVSS.n3418 VSUBS 0.131596f
C3189 AVSS.n3419 VSUBS 0.111365f
C3190 AVSS.n3422 VSUBS 0.013002f
C3191 AVSS.t109 VSUBS 1.58362f
C3192 AVSS.n3426 VSUBS 0.014231f
C3193 AVSS.n3431 VSUBS 0.015863f
C3194 AVSS.n3455 VSUBS 0.013536f
C3195 AVSS.n3456 VSUBS 0.013536f
C3196 AVSS.n3457 VSUBS 0.014085f
C3197 AVSS.n3458 VSUBS 0.014085f
C3198 AVSS.n3472 VSUBS 0.014104f
C3199 AVSS.n3473 VSUBS 0.014104f
C3200 AVSS.n3475 VSUBS 0.015863f
C3201 AVSS.n3490 VSUBS 0.015203f
C3202 AVSS.n3491 VSUBS 0.015203f
C3203 AVSS.n3492 VSUBS 0.014231f
C3204 AVSS.n3507 VSUBS 0.010886f
C3205 AVSS.n3510 VSUBS 0.02533f
C3206 AVSS.n3511 VSUBS 0.010777f
C3207 AVSS.n3512 VSUBS 0.017108f
C3208 AVSS.n3513 VSUBS 0.013464f
C3209 AVSS.n3515 VSUBS 0.013197f
C3210 AVSS.n3516 VSUBS 0.013464f
C3211 AVSS.n3518 VSUBS 0.013464f
C3212 AVSS.n3519 VSUBS 0.013197f
C3213 AVSS.n3520 VSUBS 0.016888f
C3214 AVSS.n3521 VSUBS 0.013197f
C3215 AVSS.n3522 VSUBS 0.013464f
C3216 AVSS.n3523 VSUBS 0.253149f
C3217 AVSS.n3524 VSUBS 0.013464f
C3218 AVSS.n3525 VSUBS 0.013197f
C3219 AVSS.n3526 VSUBS 0.013464f
C3220 AVSS.n3527 VSUBS 0.212363f
C3221 AVSS.n3528 VSUBS 0.190102f
C3222 AVSS.n3529 VSUBS 0.257281f
C3223 AVSS.n3530 VSUBS 0.013464f
C3224 AVSS.n3531 VSUBS 0.013464f
C3225 AVSS.n3532 VSUBS 0.013197f
C3226 AVSS.n3533 VSUBS 0.013464f
C3227 AVSS.n3534 VSUBS 0.257281f
C3228 AVSS.n3535 VSUBS 0.013464f
C3229 AVSS.n3536 VSUBS 0.01932f
C3230 AVSS.n3537 VSUBS 0.013197f
C3231 AVSS.n3538 VSUBS 0.013464f
C3232 AVSS.n3539 VSUBS 0.013197f
C3233 AVSS.n3541 VSUBS 0.013464f
C3234 AVSS.n3542 VSUBS 0.013197f
C3235 AVSS.n3545 VSUBS 0.013464f
C3236 AVSS.n3546 VSUBS 0.013464f
C3237 AVSS.n3547 VSUBS 0.013197f
C3238 AVSS.n3548 VSUBS 0.013197f
C3239 AVSS.n3549 VSUBS 0.013197f
C3240 AVSS.n3550 VSUBS 0.013464f
C3241 AVSS.n3552 VSUBS 0.013464f
C3242 AVSS.n3553 VSUBS 0.013464f
C3243 AVSS.n3554 VSUBS 0.013197f
C3244 AVSS.n3555 VSUBS 0.013197f
C3245 AVSS.n3556 VSUBS 0.013197f
C3246 AVSS.n3557 VSUBS 0.013464f
C3247 AVSS.n3559 VSUBS 0.013464f
C3248 AVSS.n3560 VSUBS 0.019496f
C3249 AVSS.n3561 VSUBS 0.415938f
C3250 AVSS.n3562 VSUBS 0.021345f
C3251 AVSS.n3563 VSUBS 0.021004f
C3252 AVSS.n3564 VSUBS 0.013197f
C3253 AVSS.n3565 VSUBS 0.013197f
C3254 AVSS.n3566 VSUBS 0.013464f
C3255 AVSS.n3567 VSUBS 0.257281f
C3256 AVSS.n3568 VSUBS 0.257281f
C3257 AVSS.n3569 VSUBS 0.257281f
C3258 AVSS.n3570 VSUBS 0.013464f
C3259 AVSS.n3571 VSUBS 0.013197f
C3260 AVSS.n3572 VSUBS 0.013197f
C3261 AVSS.n3573 VSUBS 0.013197f
C3262 AVSS.n3574 VSUBS 0.013464f
C3263 AVSS.n3575 VSUBS 1.54076f
C3264 AVSS.n3576 VSUBS 0.021194f
C3265 AVSS.n3577 VSUBS 0.013197f
C3266 AVSS.n3578 VSUBS 0.013464f
C3267 AVSS.n3579 VSUBS 0.253149f
C3268 AVSS.n3580 VSUBS 0.013464f
C3269 AVSS.n3581 VSUBS 0.013197f
C3270 AVSS.n3582 VSUBS 0.013464f
C3271 AVSS.n3583 VSUBS 0.253149f
C3272 AVSS.n3584 VSUBS 0.013464f
C3273 AVSS.n3585 VSUBS 0.013197f
C3274 AVSS.n3586 VSUBS 0.013197f
C3275 AVSS.n3587 VSUBS 0.013197f
C3276 AVSS.n3588 VSUBS 0.013464f
C3277 AVSS.n3589 VSUBS 0.253149f
C3278 AVSS.n3590 VSUBS 0.253149f
C3279 AVSS.n3591 VSUBS 4.21714f
C3280 AVSS.n3592 VSUBS 0.019048f
C3281 AVSS.n3593 VSUBS 0.018889f
C3282 AVSS.n3594 VSUBS 0.020848f
C3283 AVSS.n3595 VSUBS 0.013197f
C3284 AVSS.n3596 VSUBS 0.013464f
C3285 AVSS.n3597 VSUBS 0.257281f
C3286 AVSS.n3598 VSUBS 0.257281f
C3287 AVSS.n3599 VSUBS 0.257281f
C3288 AVSS.n3600 VSUBS 0.013464f
C3289 AVSS.n3601 VSUBS 0.013197f
C3290 AVSS.n3602 VSUBS 0.013197f
C3291 AVSS.n3603 VSUBS 0.013197f
C3292 AVSS.n3604 VSUBS 0.013464f
C3293 AVSS.n3605 VSUBS 0.19582f
C3294 AVSS.t110 VSUBS 0.312647f
C3295 AVSS.n3606 VSUBS 0.167359f
C3296 AVSS.n3607 VSUBS 0.253149f
C3297 AVSS.n3608 VSUBS 0.013464f
C3298 AVSS.n3609 VSUBS 0.013197f
C3299 AVSS.n3610 VSUBS 0.013197f
C3300 AVSS.n3611 VSUBS 0.013197f
C3301 AVSS.n3612 VSUBS 0.013464f
C3302 AVSS.n3613 VSUBS 0.253149f
C3303 AVSS.n3614 VSUBS 0.253149f
C3304 AVSS.n3615 VSUBS 0.253149f
C3305 AVSS.n3616 VSUBS 0.013464f
C3306 AVSS.n3617 VSUBS 0.013197f
C3307 AVSS.n3618 VSUBS 0.016685f
C3308 AVSS.n3619 VSUBS 0.014549f
C3309 AVSS.n3620 VSUBS 0.014676f
C3310 AVSS.n3622 VSUBS 0.013464f
C3311 AVSS.n3624 VSUBS 0.013464f
C3312 AVSS.n3625 VSUBS 0.013197f
C3313 AVSS.n3626 VSUBS 0.013197f
C3314 AVSS.n3627 VSUBS 0.012464f
C3315 AVSS.n3628 VSUBS 0.013464f
C3316 AVSS.n3630 VSUBS 0.013464f
C3317 AVSS.n3632 VSUBS 0.013464f
C3318 AVSS.n3633 VSUBS 0.013197f
C3319 AVSS.n3634 VSUBS 0.013197f
C3320 AVSS.n3635 VSUBS 0.013197f
C3321 AVSS.n3636 VSUBS 0.013464f
C3322 AVSS.n3638 VSUBS 0.013464f
C3323 AVSS.n3639 VSUBS 0.013464f
C3324 AVSS.n3641 VSUBS 0.043818f
C3325 AVSS.n3642 VSUBS 0.067428f
C3326 AVSS.n3643 VSUBS 0.165515f
C3327 AVSS.n3644 VSUBS 0.051397f
C3328 AVSS.n3646 VSUBS 0.027674f
C3329 AVSS.n3647 VSUBS 0.051249f
C3330 AVSS.n3648 VSUBS 0.093787f
C3331 AVSS.n3649 VSUBS 0.205814f
C3332 AVSS.n3650 VSUBS 0.04266f
C3333 AVSS.n3652 VSUBS 0.049199f
C3334 AVSS.n3654 VSUBS 0.051397f
C3335 AVSS.n3656 VSUBS 0.021116f
C3336 AVSS.n3657 VSUBS 0.045176f
C3337 AVSS.n3658 VSUBS 0.037539f
C3338 AVSS.n3659 VSUBS 0.017666f
C3339 AVSS.n3660 VSUBS 0.077272f
C3340 AVSS.n3662 VSUBS 0.039103f
C3341 AVSS.n3663 VSUBS 0.06022f
C3342 AVSS.n3664 VSUBS 0.084482f
C3343 AVSS.n3665 VSUBS 0.038321f
C3344 AVSS.n3666 VSUBS 0.160194f
C3345 AVSS.n3667 VSUBS 0.032065f
C3346 AVSS.n3669 VSUBS 0.046257f
C3347 AVSS.n3670 VSUBS 0.013957f
C3348 AVSS.n3672 VSUBS 0.053022f
C3349 AVSS.n3673 VSUBS 0.030324f
C3350 AVSS.n3674 VSUBS 0.032543f
C3351 AVSS.n3675 VSUBS 0.070566f
C3352 AVSS.n3676 VSUBS 0.11133f
C3353 AVSS.n3677 VSUBS 0.075408f
C3354 AVSS.n3678 VSUBS 0.017925f
C3355 AVSS.n3679 VSUBS 0.013197f
C3356 AVSS.n3680 VSUBS 0.013464f
C3357 AVSS.n3681 VSUBS 0.013464f
C3358 AVSS.n3682 VSUBS 0.013197f
C3359 AVSS.n3684 VSUBS 0.013464f
C3360 AVSS.n3685 VSUBS 0.013197f
C3361 AVSS.n3687 VSUBS 0.013464f
C3362 AVSS.n3688 VSUBS 0.013197f
C3363 AVSS.n3690 VSUBS 0.014835f
C3364 AVSS.n3691 VSUBS 0.013197f
C3365 AVSS.n3692 VSUBS 0.013464f
C3366 AVSS.n3694 VSUBS 0.013464f
C3367 AVSS.n3695 VSUBS 0.013197f
C3368 AVSS.n3696 VSUBS 0.016888f
C3369 AVSS.n3697 VSUBS 0.013197f
C3370 AVSS.n3698 VSUBS 0.013464f
C3371 AVSS.n3699 VSUBS 0.253149f
C3372 AVSS.n3700 VSUBS 0.013464f
C3373 AVSS.n3701 VSUBS 0.013197f
C3374 AVSS.n3702 VSUBS 0.013464f
C3375 AVSS.n3703 VSUBS 0.253149f
C3376 AVSS.n3704 VSUBS 0.013464f
C3377 AVSS.n3705 VSUBS 0.013197f
C3378 AVSS.n3706 VSUBS 0.013464f
C3379 AVSS.n3707 VSUBS 0.019048f
C3380 AVSS.n3708 VSUBS 0.013197f
C3381 AVSS.n3709 VSUBS 0.013197f
C3382 AVSS.n3710 VSUBS 0.013464f
C3383 AVSS.n3711 VSUBS 0.013197f
C3384 AVSS.n3713 VSUBS 0.013464f
C3385 AVSS.n3714 VSUBS 0.013197f
C3386 AVSS.n3715 VSUBS 0.013197f
C3387 AVSS.n3716 VSUBS 0.013464f
C3388 AVSS.n3718 VSUBS 0.013464f
C3389 AVSS.n3720 VSUBS 0.013464f
C3390 AVSS.n3721 VSUBS 0.013197f
C3391 AVSS.n3722 VSUBS 0.013197f
C3392 AVSS.n3723 VSUBS 0.013197f
C3393 AVSS.n3724 VSUBS 0.013464f
C3394 AVSS.n3726 VSUBS 0.013464f
C3395 AVSS.n3727 VSUBS 0.013464f
C3396 AVSS.n3729 VSUBS 0.021194f
C3397 AVSS.n3730 VSUBS 0.020848f
C3398 AVSS.n3731 VSUBS 0.018889f
C3399 AVSS.n3732 VSUBS 0.013197f
C3400 AVSS.n3733 VSUBS 0.013464f
C3401 AVSS.n3734 VSUBS 0.253149f
C3402 AVSS.n3735 VSUBS 0.253149f
C3403 AVSS.n3736 VSUBS 0.253149f
C3404 AVSS.n3737 VSUBS 0.013464f
C3405 AVSS.n3738 VSUBS 0.013197f
C3406 AVSS.n3739 VSUBS 0.013197f
C3407 AVSS.n3740 VSUBS 0.013197f
C3408 AVSS.n3741 VSUBS 0.013464f
C3409 AVSS.n3742 VSUBS 0.212363f
C3410 AVSS.t108 VSUBS 0.243736f
C3411 AVSS.n3743 VSUBS 0.167359f
C3412 AVSS.n3744 VSUBS 0.253149f
C3413 AVSS.n3745 VSUBS 0.013464f
C3414 AVSS.n3746 VSUBS 0.013197f
C3415 AVSS.n3747 VSUBS 0.013197f
C3416 AVSS.n3748 VSUBS 0.013197f
C3417 AVSS.n3749 VSUBS 0.013464f
C3418 AVSS.n3750 VSUBS 0.253149f
C3419 AVSS.n3751 VSUBS 0.253149f
C3420 AVSS.n3752 VSUBS 0.253149f
C3421 AVSS.n3753 VSUBS 0.013464f
C3422 AVSS.n3754 VSUBS 0.013197f
C3423 AVSS.n3755 VSUBS 0.016685f
C3424 AVSS.n3756 VSUBS 0.014549f
C3425 AVSS.n3757 VSUBS 0.014676f
C3426 AVSS.n3759 VSUBS 0.013464f
C3427 AVSS.n3761 VSUBS 0.013464f
C3428 AVSS.n3762 VSUBS 0.013197f
C3429 AVSS.n3763 VSUBS 0.013197f
C3430 AVSS.n3764 VSUBS 0.012464f
C3431 AVSS.n3765 VSUBS 0.013464f
C3432 AVSS.n3767 VSUBS 0.013464f
C3433 AVSS.n3769 VSUBS 0.013464f
C3434 AVSS.n3770 VSUBS 0.013197f
C3435 AVSS.n3771 VSUBS 0.013197f
C3436 AVSS.n3772 VSUBS 0.013197f
C3437 AVSS.n3773 VSUBS 0.013464f
C3438 AVSS.n3775 VSUBS 0.013464f
C3439 AVSS.n3777 VSUBS 0.013464f
C3440 AVSS.n3781 VSUBS 0.013002f
C3441 AVSS.t107 VSUBS 1.58362f
C3442 AVSS.n3785 VSUBS 0.014231f
C3443 AVSS.n3790 VSUBS 0.015863f
C3444 AVSS.n3814 VSUBS 0.013536f
C3445 AVSS.n3815 VSUBS 0.013536f
C3446 AVSS.n3816 VSUBS 0.014085f
C3447 AVSS.n3817 VSUBS 0.014085f
C3448 AVSS.n3831 VSUBS 0.014104f
C3449 AVSS.n3832 VSUBS 0.014104f
C3450 AVSS.n3834 VSUBS 0.015863f
C3451 AVSS.n3849 VSUBS 0.015203f
C3452 AVSS.n3851 VSUBS 0.011838f
C3453 AVSS.n3867 VSUBS 0.010886f
C3454 AVSS.n3870 VSUBS 0.075481f
C3455 AVSS.n3871 VSUBS 0.0905f
C3456 AVSS.n3872 VSUBS 0.205814f
C3457 AVSS.n3873 VSUBS 0.051397f
C3458 AVSS.n3874 VSUBS 0.0905f
C3459 AVSS.n3875 VSUBS 0.186635f
C3460 AVSS.n3876 VSUBS 0.189601f
C3461 AVSS.n3877 VSUBS 0.077272f
C3462 AVSS.n3878 VSUBS 0.051397f
C3463 AVSS.n3879 VSUBS 0.046257f
C3464 AVSS.n3880 VSUBS 0.0905f
C3465 AVSS.n3881 VSUBS 0.0905f
C3466 AVSS.n3882 VSUBS 0.030324f
C3467 AVSS.n3883 VSUBS 0.04266f
C3468 AVSS.n3884 VSUBS 0.067428f
C3469 AVSS.n3885 VSUBS 0.210564f
C3470 AVSS.n3886 VSUBS 0.192186f
C3471 AVSS.n3887 VSUBS 0.114184f
C3472 AVSS.n3888 VSUBS 0.075408f
C3473 AVSS.n3889 VSUBS 0.017925f
C3474 AVSS.n3890 VSUBS 0.013197f
C3475 AVSS.n3891 VSUBS 0.013464f
C3476 AVSS.n3892 VSUBS 0.013464f
C3477 AVSS.n3893 VSUBS 0.013197f
C3478 AVSS.n3895 VSUBS 0.013464f
C3479 AVSS.n3896 VSUBS 0.013197f
C3480 AVSS.n3898 VSUBS 0.013464f
C3481 AVSS.n3899 VSUBS 0.013197f
C3482 AVSS.n3901 VSUBS 0.014835f
C3483 AVSS.n3902 VSUBS 0.013197f
C3484 AVSS.n3903 VSUBS 0.013464f
C3485 AVSS.n3905 VSUBS 0.013464f
C3486 AVSS.n3906 VSUBS 0.013197f
C3487 AVSS.n3907 VSUBS 0.016888f
C3488 AVSS.n3908 VSUBS 0.013197f
C3489 AVSS.n3909 VSUBS 0.013464f
C3490 AVSS.n3910 VSUBS 0.253149f
C3491 AVSS.n3911 VSUBS 0.013464f
C3492 AVSS.n3912 VSUBS 0.013197f
C3493 AVSS.n3913 VSUBS 0.013464f
C3494 AVSS.n3914 VSUBS 0.253149f
C3495 AVSS.n3915 VSUBS 0.013464f
C3496 AVSS.n3916 VSUBS 0.013197f
C3497 AVSS.n3917 VSUBS 0.013464f
C3498 AVSS.n3918 VSUBS 0.019048f
C3499 AVSS.n3919 VSUBS 0.013197f
C3500 AVSS.n3920 VSUBS 0.013197f
C3501 AVSS.n3921 VSUBS 0.013464f
C3502 AVSS.n3922 VSUBS 0.013197f
C3503 AVSS.n3924 VSUBS 0.013464f
C3504 AVSS.n3925 VSUBS 0.013197f
C3505 AVSS.n3926 VSUBS 0.013197f
C3506 AVSS.n3927 VSUBS 0.013464f
C3507 AVSS.n3929 VSUBS 0.013464f
C3508 AVSS.n3931 VSUBS 0.013464f
C3509 AVSS.n3932 VSUBS 0.013197f
C3510 AVSS.n3933 VSUBS 0.013197f
C3511 AVSS.n3934 VSUBS 0.013197f
C3512 AVSS.n3935 VSUBS 0.013464f
C3513 AVSS.n3937 VSUBS 0.013464f
C3514 AVSS.n3938 VSUBS 0.013464f
C3515 AVSS.n3940 VSUBS 0.021194f
C3516 AVSS.n3941 VSUBS 0.020848f
C3517 AVSS.n3942 VSUBS 0.018889f
C3518 AVSS.n3943 VSUBS 0.013197f
C3519 AVSS.n3944 VSUBS 0.013464f
C3520 AVSS.n3945 VSUBS 0.253149f
C3521 AVSS.n3946 VSUBS 0.253149f
C3522 AVSS.n3947 VSUBS 0.253149f
C3523 AVSS.n3948 VSUBS 0.013464f
C3524 AVSS.n3949 VSUBS 0.013197f
C3525 AVSS.n3950 VSUBS 0.013197f
C3526 AVSS.n3951 VSUBS 0.013197f
C3527 AVSS.n3952 VSUBS 0.013464f
C3528 AVSS.n3953 VSUBS 0.212363f
C3529 AVSS.t95 VSUBS 0.243736f
C3530 AVSS.n3954 VSUBS 0.167359f
C3531 AVSS.n3955 VSUBS 0.253149f
C3532 AVSS.n3956 VSUBS 0.013464f
C3533 AVSS.n3957 VSUBS 0.013197f
C3534 AVSS.n3958 VSUBS 0.013197f
C3535 AVSS.n3959 VSUBS 0.013197f
C3536 AVSS.n3960 VSUBS 0.013464f
C3537 AVSS.n3961 VSUBS 0.253149f
C3538 AVSS.n3962 VSUBS 0.253149f
C3539 AVSS.n3963 VSUBS 0.253149f
C3540 AVSS.n3964 VSUBS 0.013464f
C3541 AVSS.n3965 VSUBS 0.013197f
C3542 AVSS.n3966 VSUBS 0.016685f
C3543 AVSS.n3967 VSUBS 0.014549f
C3544 AVSS.n3968 VSUBS 0.014676f
C3545 AVSS.n3970 VSUBS 0.013464f
C3546 AVSS.n3972 VSUBS 0.013464f
C3547 AVSS.n3973 VSUBS 0.013197f
C3548 AVSS.n3974 VSUBS 0.013197f
C3549 AVSS.n3975 VSUBS 0.012464f
C3550 AVSS.n3976 VSUBS 0.013464f
C3551 AVSS.n3978 VSUBS 0.013464f
C3552 AVSS.n3980 VSUBS 0.013464f
C3553 AVSS.n3981 VSUBS 0.013197f
C3554 AVSS.n3982 VSUBS 0.013197f
C3555 AVSS.n3983 VSUBS 0.013197f
C3556 AVSS.n3984 VSUBS 0.013464f
C3557 AVSS.n3986 VSUBS 0.013464f
C3558 AVSS.n3988 VSUBS 0.013464f
C3559 AVSS.n3992 VSUBS 0.013002f
C3560 AVSS.t94 VSUBS 1.58362f
C3561 AVSS.n3996 VSUBS 0.014231f
C3562 AVSS.n4001 VSUBS 0.015863f
C3563 AVSS.n4025 VSUBS 0.013536f
C3564 AVSS.n4026 VSUBS 0.013536f
C3565 AVSS.n4027 VSUBS 0.014085f
C3566 AVSS.n4028 VSUBS 0.014085f
C3567 AVSS.n4042 VSUBS 0.014104f
C3568 AVSS.n4043 VSUBS 0.014104f
C3569 AVSS.n4045 VSUBS 0.015863f
C3570 AVSS.n4060 VSUBS 0.015203f
C3571 AVSS.n4062 VSUBS 0.011838f
C3572 AVSS.n4078 VSUBS 0.010886f
C3573 AVSS.n4081 VSUBS 0.075481f
C3574 AVSS.n4082 VSUBS 0.0905f
C3575 AVSS.n4083 VSUBS 0.205814f
C3576 AVSS.n4084 VSUBS 0.051397f
C3577 AVSS.n4085 VSUBS 0.0905f
C3578 AVSS.n4086 VSUBS 0.186635f
C3579 AVSS.n4087 VSUBS 0.189601f
C3580 AVSS.n4088 VSUBS 0.077272f
C3581 AVSS.n4089 VSUBS 0.051397f
C3582 AVSS.n4090 VSUBS 0.046257f
C3583 AVSS.n4091 VSUBS 0.0905f
C3584 AVSS.n4092 VSUBS 0.0905f
C3585 AVSS.n4093 VSUBS 0.030324f
C3586 AVSS.n4094 VSUBS 0.04266f
C3587 AVSS.n4095 VSUBS 0.067428f
C3588 AVSS.n4096 VSUBS 0.210564f
C3589 AVSS.n4097 VSUBS 0.192186f
C3590 AVSS.n4098 VSUBS 0.0905f
C3591 AVSS.n4099 VSUBS 0.051397f
C3592 AVSS.n4100 VSUBS 0.0905f
C3593 AVSS.n4101 VSUBS 0.067428f
C3594 AVSS.n4102 VSUBS 0.210564f
C3595 AVSS.n4103 VSUBS 0.205814f
C3596 AVSS.n4104 VSUBS 0.04266f
C3597 AVSS.n4105 VSUBS 0.030324f
C3598 AVSS.n4106 VSUBS 0.0905f
C3599 AVSS.n4107 VSUBS 0.0905f
C3600 AVSS.n4108 VSUBS 0.046257f
C3601 AVSS.n4109 VSUBS 0.051397f
C3602 AVSS.n4110 VSUBS 0.077272f
C3603 AVSS.n4111 VSUBS 0.189601f
C3604 AVSS.n4112 VSUBS 0.186635f
C3605 AVSS.n4113 VSUBS 0.114184f
C3606 AVSS.n4116 VSUBS 0.015203f
C3607 AVSS.n4150 VSUBS 0.010886f
C3608 AVSS.n4151 VSUBS 0.013002f
C3609 AVSS.n4167 VSUBS 0.013536f
C3610 AVSS.n4168 VSUBS 0.013536f
C3611 AVSS.n4169 VSUBS 0.014085f
C3612 AVSS.n4170 VSUBS 0.014085f
C3613 AVSS.n4184 VSUBS 0.014104f
C3614 AVSS.n4185 VSUBS 0.014104f
C3615 AVSS.n4186 VSUBS 0.015863f
C3616 AVSS.n4187 VSUBS 0.015863f
C3617 AVSS.t101 VSUBS 1.58362f
C3618 AVSS.n4202 VSUBS 0.014231f
C3619 AVSS.n4204 VSUBS 0.011838f
C3620 AVSS.n4205 VSUBS 0.075408f
C3621 AVSS.n4206 VSUBS 0.017925f
C3622 AVSS.n4207 VSUBS 0.013197f
C3623 AVSS.n4208 VSUBS 0.013464f
C3624 AVSS.n4209 VSUBS 0.013197f
C3625 AVSS.n4210 VSUBS 0.013464f
C3626 AVSS.n4211 VSUBS 0.013197f
C3627 AVSS.n4213 VSUBS 0.013464f
C3628 AVSS.n4215 VSUBS 0.013464f
C3629 AVSS.n4216 VSUBS 0.013197f
C3630 AVSS.n4217 VSUBS 0.013197f
C3631 AVSS.n4218 VSUBS 0.013197f
C3632 AVSS.n4219 VSUBS 0.013464f
C3633 AVSS.n4221 VSUBS 0.013464f
C3634 AVSS.n4223 VSUBS 0.013464f
C3635 AVSS.n4224 VSUBS 0.013197f
C3636 AVSS.n4225 VSUBS 0.013197f
C3637 AVSS.n4226 VSUBS 0.013197f
C3638 AVSS.n4227 VSUBS 0.013464f
C3639 AVSS.n4229 VSUBS 0.013464f
C3640 AVSS.n4231 VSUBS 0.013197f
C3641 AVSS.n4232 VSUBS 0.013464f
C3642 AVSS.n4233 VSUBS 0.013197f
C3643 AVSS.n4234 VSUBS 0.013464f
C3644 AVSS.n4235 VSUBS 0.013197f
C3645 AVSS.n4236 VSUBS 0.013197f
C3646 AVSS.n4237 VSUBS 0.013464f
C3647 AVSS.n4239 VSUBS 0.013464f
C3648 AVSS.n4241 VSUBS 0.013464f
C3649 AVSS.n4242 VSUBS 0.013197f
C3650 AVSS.n4243 VSUBS 0.013197f
C3651 AVSS.n4244 VSUBS 0.013197f
C3652 AVSS.n4245 VSUBS 0.013464f
C3653 AVSS.n4247 VSUBS 0.013464f
C3654 AVSS.n4249 VSUBS 0.013464f
C3655 AVSS.n4250 VSUBS 0.013197f
C3656 AVSS.n4251 VSUBS 0.013197f
C3657 AVSS.n4252 VSUBS 0.013197f
C3658 AVSS.n4253 VSUBS 0.013464f
C3659 AVSS.n4255 VSUBS 0.013464f
C3660 AVSS.n4256 VSUBS 0.013464f
C3661 AVSS.n4257 VSUBS 0.013197f
C3662 AVSS.n4258 VSUBS 0.01932f
C3663 AVSS.n4259 VSUBS 0.019496f
C3664 AVSS.n4260 VSUBS 0.021345f
C3665 AVSS.n4262 VSUBS 0.013464f
C3666 AVSS.n4265 VSUBS 0.018072f
C3667 AVSS.n4266 VSUBS 0.033852f
C3668 AVSS.n4267 VSUBS 0.018072f
C3669 AVSS.n4269 VSUBS 0.011633f
C3670 AVSS.n4270 VSUBS 0.017108f
C3671 AVSS.n4271 VSUBS 0.017327f
C3672 AVSS.n4273 VSUBS 0.013464f
C3673 AVSS.n4274 VSUBS 0.013464f
C3674 AVSS.n4275 VSUBS 0.013197f
C3675 AVSS.n4276 VSUBS 0.013197f
C3676 AVSS.n4277 VSUBS 0.013197f
C3677 AVSS.n4278 VSUBS 0.013464f
C3678 AVSS.n4280 VSUBS 0.013464f
C3679 AVSS.n4281 VSUBS 0.013464f
C3680 AVSS.n4282 VSUBS 0.013197f
C3681 AVSS.n4283 VSUBS 0.013197f
C3682 AVSS.n4284 VSUBS 0.013197f
C3683 AVSS.n4285 VSUBS 0.013464f
C3684 AVSS.n4287 VSUBS 0.013464f
C3685 AVSS.n4288 VSUBS 0.013464f
C3686 AVSS.n4289 VSUBS 0.013197f
C3687 AVSS.n4290 VSUBS 0.013197f
C3688 AVSS.n4291 VSUBS 0.01932f
C3689 AVSS.n4292 VSUBS 0.019496f
C3690 AVSS.n4293 VSUBS 0.021345f
C3691 AVSS.n4295 VSUBS 0.013464f
C3692 AVSS.n4298 VSUBS 0.018072f
C3693 AVSS.n4299 VSUBS 0.033852f
C3694 AVSS.n4300 VSUBS 0.018072f
C3695 AVSS.n4302 VSUBS 0.011633f
C3696 AVSS.n4303 VSUBS 0.017108f
C3697 AVSS.n4304 VSUBS 0.017327f
C3698 AVSS.n4306 VSUBS 0.013464f
C3699 AVSS.n4307 VSUBS 0.013464f
C3700 AVSS.n4308 VSUBS 0.013197f
C3701 AVSS.n4309 VSUBS 0.013197f
C3702 AVSS.n4310 VSUBS 0.013197f
C3703 AVSS.n4311 VSUBS 0.013464f
C3704 AVSS.n4313 VSUBS 0.013464f
C3705 AVSS.n4314 VSUBS 0.013464f
C3706 AVSS.n4315 VSUBS 0.013197f
C3707 AVSS.n4316 VSUBS 0.013197f
C3708 AVSS.n4317 VSUBS 0.013197f
C3709 AVSS.n4318 VSUBS 0.013464f
C3710 AVSS.n4320 VSUBS 0.013464f
C3711 AVSS.n4321 VSUBS 0.013464f
C3712 AVSS.n4322 VSUBS 0.013197f
C3713 AVSS.n4323 VSUBS 0.013197f
C3714 AVSS.n4324 VSUBS 0.01932f
C3715 AVSS.n4325 VSUBS 0.019496f
C3716 AVSS.n4326 VSUBS 0.021345f
C3717 AVSS.n4328 VSUBS 0.013464f
C3718 AVSS.n4331 VSUBS 0.018072f
C3719 AVSS.n4332 VSUBS 0.03378f
C3720 AVSS.n4333 VSUBS 0.017999f
C3721 AVSS.n4335 VSUBS 0.011633f
C3722 AVSS.n4336 VSUBS 0.014835f
C3723 AVSS.n4337 VSUBS 0.017327f
C3724 AVSS.n4339 VSUBS 0.013464f
C3725 AVSS.n4342 VSUBS 0.014516f
C3726 AVSS.n4343 VSUBS 0.033888f
C3727 AVSS.n4344 VSUBS 0.018072f
C3728 AVSS.n4346 VSUBS 0.014549f
C3729 AVSS.n4347 VSUBS 0.013464f
C3730 AVSS.n4348 VSUBS 0.012464f
C3731 AVSS.n4349 VSUBS 0.013464f
C3732 AVSS.n4350 VSUBS 0.013197f
C3733 AVSS.n4351 VSUBS 0.013464f
C3734 AVSS.n4352 VSUBS 0.017108f
C3735 AVSS.n4353 VSUBS 0.013464f
C3736 AVSS.n4354 VSUBS 0.013197f
C3737 AVSS.n4355 VSUBS 0.013464f
C3738 AVSS.n4356 VSUBS 0.013197f
C3739 AVSS.n4357 VSUBS 0.013464f
C3740 AVSS.n4358 VSUBS 0.01932f
C3741 AVSS.n4359 VSUBS 0.013464f
C3742 AVSS.n4360 VSUBS 0.021004f
C3743 AVSS.n4361 VSUBS 0.257281f
C3744 AVSS.n4362 VSUBS 0.013464f
C3745 AVSS.n4363 VSUBS 0.013197f
C3746 AVSS.n4364 VSUBS 0.013197f
C3747 AVSS.n4365 VSUBS 0.013464f
C3748 AVSS.n4366 VSUBS 0.013197f
C3749 AVSS.n4367 VSUBS 0.257281f
C3750 AVSS.n4368 VSUBS 0.013464f
C3751 AVSS.n4369 VSUBS 0.013197f
C3752 AVSS.n4370 VSUBS 0.410221f
C3753 AVSS.n4371 VSUBS 0.257281f
C3754 AVSS.n4372 VSUBS 0.013464f
C3755 AVSS.n4373 VSUBS 0.013197f
C3756 AVSS.n4374 VSUBS 0.013197f
C3757 AVSS.n4375 VSUBS 0.013197f
C3758 AVSS.n4376 VSUBS 0.013464f
C3759 AVSS.n4377 VSUBS 0.257281f
C3760 AVSS.n4378 VSUBS 0.257281f
C3761 AVSS.n4379 VSUBS 0.19582f
C3762 AVSS.n4380 VSUBS 0.013464f
C3763 AVSS.n4381 VSUBS 0.013464f
C3764 AVSS.n4382 VSUBS 0.190102f
C3765 AVSS.n4383 VSUBS 0.257281f
C3766 AVSS.n4384 VSUBS 0.013464f
C3767 AVSS.n4385 VSUBS 0.013197f
C3768 AVSS.n4386 VSUBS 0.013197f
C3769 AVSS.n4387 VSUBS 0.013197f
C3770 AVSS.n4388 VSUBS 0.013464f
C3771 AVSS.n4389 VSUBS 0.257281f
C3772 AVSS.n4390 VSUBS 0.257281f
C3773 AVSS.n4391 VSUBS 0.415938f
C3774 AVSS.n4392 VSUBS 0.021345f
C3775 AVSS.n4393 VSUBS 0.019496f
C3776 AVSS.n4395 VSUBS 0.013464f
C3777 AVSS.n4396 VSUBS 0.013197f
C3778 AVSS.n4397 VSUBS 0.013197f
C3779 AVSS.n4398 VSUBS 0.013197f
C3780 AVSS.n4399 VSUBS 0.013464f
C3781 AVSS.n4401 VSUBS 0.013464f
C3782 AVSS.n4403 VSUBS 0.013464f
C3783 AVSS.n4404 VSUBS 0.013197f
C3784 AVSS.n4405 VSUBS 0.013197f
C3785 AVSS.n4406 VSUBS 0.013197f
C3786 AVSS.n4407 VSUBS 0.013464f
C3787 AVSS.n4409 VSUBS 0.013464f
C3788 AVSS.n4411 VSUBS 0.013464f
C3789 AVSS.n4412 VSUBS 0.013197f
C3790 AVSS.n4413 VSUBS 0.010705f
C3791 AVSS.n4416 VSUBS 0.013464f
C3792 AVSS.n4418 VSUBS 0.017327f
C3793 AVSS.n4420 VSUBS 0.014835f
C3794 AVSS.n4421 VSUBS 0.014713f
C3795 AVSS.n4422 VSUBS 0.013197f
C3796 AVSS.n4423 VSUBS 0.013197f
C3797 AVSS.n4424 VSUBS 0.013464f
C3798 AVSS.n4426 VSUBS 0.013464f
C3799 AVSS.n4428 VSUBS 0.013464f
C3800 AVSS.n4429 VSUBS 0.013197f
C3801 AVSS.n4430 VSUBS 0.013197f
C3802 AVSS.n4432 VSUBS 0.013464f
C3803 AVSS.n4434 VSUBS 0.013464f
C3804 AVSS.n4436 VSUBS 0.013464f
C3805 AVSS.n4437 VSUBS 0.013197f
C3806 AVSS.n4438 VSUBS 0.013197f
C3807 AVSS.n4439 VSUBS 0.013197f
C3808 AVSS.n4440 VSUBS 0.013464f
C3809 AVSS.n4442 VSUBS 0.014676f
C3810 AVSS.n4443 VSUBS 0.016888f
C3811 AVSS.n4444 VSUBS 0.016685f
C3812 AVSS.n4446 VSUBS 0.013464f
C3813 AVSS.n4447 VSUBS 0.013464f
C3814 AVSS.n4448 VSUBS 0.010705f
C3815 AVSS.n4449 VSUBS 0.013197f
C3816 AVSS.n4450 VSUBS 0.013464f
C3817 AVSS.n4451 VSUBS 0.013464f
C3818 AVSS.n4452 VSUBS 0.013197f
C3819 AVSS.n4453 VSUBS 0.013197f
C3820 AVSS.n4454 VSUBS 0.013464f
C3821 AVSS.n4455 VSUBS 0.013464f
C3822 AVSS.n4456 VSUBS 0.013197f
C3823 AVSS.n4457 VSUBS 0.013197f
C3824 AVSS.n4458 VSUBS 0.013464f
C3825 AVSS.n4459 VSUBS 0.013464f
C3826 AVSS.n4460 VSUBS 0.013197f
C3827 AVSS.n4461 VSUBS 0.013197f
C3828 AVSS.n4462 VSUBS 0.013464f
C3829 AVSS.n4463 VSUBS 0.013464f
C3830 AVSS.n4464 VSUBS 0.013197f
C3831 AVSS.n4465 VSUBS 0.013197f
C3832 AVSS.n4466 VSUBS 0.018889f
C3833 AVSS.n4467 VSUBS 0.019048f
C3834 AVSS.n4468 VSUBS 0.863324f
C3835 AVSS.n4470 VSUBS 0.013464f
C3836 AVSS.n4471 VSUBS 0.013197f
C3837 AVSS.n4472 VSUBS 0.016685f
C3838 AVSS.n4473 VSUBS 0.014549f
C3839 AVSS.n4474 VSUBS 0.014676f
C3840 AVSS.n4476 VSUBS 0.135542f
C3841 AVSS.n4477 VSUBS 0.205976f
C3842 AVSS.n4478 VSUBS 0.205814f
C3843 AVSS.n4479 VSUBS 0.046257f
C3844 AVSS.n4480 VSUBS 0.066046f
C3845 AVSS.n4481 VSUBS 0.067394f
C3846 AVSS.n4482 VSUBS 0.067394f
C3847 AVSS.n4483 VSUBS 0.051397f
C3848 AVSS.n4486 VSUBS 0.077272f
C3849 AVSS.n4487 VSUBS 0.04266f
C3850 AVSS.n4489 VSUBS 0.093787f
C3851 AVSS.n4490 VSUBS 0.067428f
C3852 AVSS.n4492 VSUBS 0.084482f
C3853 AVSS.n4493 VSUBS 0.160158f
C3854 AVSS.n4494 VSUBS 0.075481f
C3855 AVSS.n4495 VSUBS 0.030324f
C3856 AVSS.n4496 VSUBS 0.051397f
C3857 AVSS.n4497 VSUBS 0.045828f
C3858 AVSS.n4498 VSUBS 0.135542f
C3859 AVSS.n4500 VSUBS 0.013464f
C3860 AVSS.n4501 VSUBS 0.013197f
C3861 AVSS.n4502 VSUBS 0.014713f
C3862 AVSS.n4503 VSUBS 0.017108f
C3863 AVSS.n4504 VSUBS 0.017327f
C3864 AVSS.n4506 VSUBS 0.013464f
C3865 AVSS.n4507 VSUBS 0.013464f
C3866 AVSS.n4508 VSUBS 0.013197f
C3867 AVSS.n4509 VSUBS 0.013197f
C3868 AVSS.n4510 VSUBS 0.013197f
C3869 AVSS.n4511 VSUBS 0.013464f
C3870 AVSS.n4513 VSUBS 0.013464f
C3871 AVSS.n4514 VSUBS 0.013464f
C3872 AVSS.n4515 VSUBS 0.013197f
C3873 AVSS.n4516 VSUBS 0.013197f
C3874 AVSS.n4517 VSUBS 0.013197f
C3875 AVSS.n4518 VSUBS 0.013464f
C3876 AVSS.n4520 VSUBS 0.013464f
C3877 AVSS.n4521 VSUBS 0.013464f
C3878 AVSS.n4522 VSUBS 0.013197f
C3879 AVSS.n4543 VSUBS 0.015203f
C3880 AVSS.n4556 VSUBS 0.014085f
C3881 AVSS.n4557 VSUBS 0.014085f
C3882 AVSS.n4558 VSUBS 0.013536f
C3883 AVSS.n4559 VSUBS 0.013536f
C3884 AVSS.n4574 VSUBS 0.013002f
C3885 AVSS.n4575 VSUBS 0.013002f
C3886 AVSS.n4576 VSUBS 0.010886f
C3887 AVSS.n4577 VSUBS 0.010886f
C3888 AVSS.n4592 VSUBS 0.014231f
C3889 AVSS.n4594 VSUBS 0.011838f
C3890 AVSS.n4596 VSUBS 0.015863f
C3891 AVSS.t112 VSUBS 1.58362f
C3892 AVSS.n4613 VSUBS 0.014104f
C3893 AVSS.n4614 VSUBS 0.010825f
C3894 AVSS.n4615 VSUBS 0.012104f
C3895 AVSS.n4616 VSUBS 0.073941f
C3896 AVSS.n4617 VSUBS 0.013197f
C3897 AVSS.n4618 VSUBS 0.135542f
C3898 AVSS.n4619 VSUBS 0.013197f
C3899 AVSS.n4620 VSUBS 0.013464f
C3900 AVSS.n4621 VSUBS 0.013197f
C3901 AVSS.n4622 VSUBS 0.013464f
C3902 AVSS.n4623 VSUBS 0.013197f
C3903 AVSS.n4624 VSUBS 0.021004f
C3904 AVSS.n4625 VSUBS 0.021345f
C3905 AVSS.n4627 VSUBS 0.013464f
C3906 AVSS.n4629 VSUBS 0.013464f
C3907 AVSS.n4630 VSUBS 0.013197f
C3908 AVSS.n4631 VSUBS 0.013197f
C3909 AVSS.n4632 VSUBS 0.013197f
C3910 AVSS.n4633 VSUBS 0.013464f
C3911 AVSS.n4635 VSUBS 0.013464f
C3912 AVSS.n4637 VSUBS 0.013464f
C3913 AVSS.n4638 VSUBS 0.013197f
C3914 AVSS.n4639 VSUBS 0.013197f
C3915 AVSS.n4640 VSUBS 0.013197f
C3916 AVSS.n4641 VSUBS 0.013464f
C3917 AVSS.n4643 VSUBS 0.013464f
C3918 AVSS.n4644 VSUBS 0.013464f
C3919 AVSS.n4646 VSUBS 0.021194f
C3920 AVSS.n4647 VSUBS 0.020848f
C3921 AVSS.n4648 VSUBS 0.017129f
C3922 AVSS.n4649 VSUBS 0.013197f
C3923 AVSS.n4650 VSUBS 0.013464f
C3924 AVSS.n4651 VSUBS 0.013464f
C3925 AVSS.n4652 VSUBS 0.013197f
C3926 AVSS.n4653 VSUBS 0.013197f
C3927 AVSS.n4654 VSUBS 0.013464f
C3928 AVSS.n4655 VSUBS 0.013464f
C3929 AVSS.n4656 VSUBS 0.013197f
C3930 AVSS.n4657 VSUBS 0.013197f
C3931 AVSS.n4658 VSUBS 0.013464f
C3932 AVSS.n4659 VSUBS 0.013464f
C3933 AVSS.n4660 VSUBS 0.013197f
C3934 AVSS.n4661 VSUBS 0.013197f
C3935 AVSS.n4662 VSUBS 0.013464f
C3936 AVSS.n4663 VSUBS 0.013464f
C3937 AVSS.n4664 VSUBS 0.013197f
C3938 AVSS.n4665 VSUBS 0.013464f
C3939 AVSS.n4668 VSUBS 0.017703f
C3940 AVSS.n4669 VSUBS 0.06892f
C3941 AVSS.n4670 VSUBS 0.01429f
C3942 AVSS.n4672 VSUBS 0.01756f
C3943 AVSS.n4673 VSUBS 0.019496f
C3944 AVSS.n4674 VSUBS 0.021345f
C3945 AVSS.n4676 VSUBS 0.013464f
C3946 AVSS.n4679 VSUBS 0.024742f
C3947 AVSS.n4680 VSUBS 0.024813f
C3948 AVSS.n4682 VSUBS 0.011633f
C3949 AVSS.n4683 VSUBS 0.017108f
C3950 AVSS.n4684 VSUBS 0.017327f
C3951 AVSS.n4686 VSUBS 0.013464f
C3952 AVSS.n4687 VSUBS 0.013464f
C3953 AVSS.n4688 VSUBS 0.013197f
C3954 AVSS.n4689 VSUBS 0.013197f
C3955 AVSS.n4690 VSUBS 0.013197f
C3956 AVSS.n4691 VSUBS 0.013464f
C3957 AVSS.n4693 VSUBS 0.013464f
C3958 AVSS.n4694 VSUBS 0.013464f
C3959 AVSS.n4695 VSUBS 0.013197f
C3960 AVSS.n4696 VSUBS 0.013197f
C3961 AVSS.n4697 VSUBS 0.013197f
C3962 AVSS.n4698 VSUBS 0.013464f
C3963 AVSS.n4700 VSUBS 0.013464f
C3964 AVSS.n4701 VSUBS 0.013464f
C3965 AVSS.n4702 VSUBS 0.013197f
C3966 AVSS.n4703 VSUBS 0.013197f
C3967 AVSS.n4704 VSUBS 0.01932f
C3968 AVSS.n4705 VSUBS 0.019496f
C3969 AVSS.n4706 VSUBS 0.021345f
C3970 AVSS.n4708 VSUBS 0.013464f
C3971 AVSS.n4711 VSUBS 0.024742f
C3972 AVSS.n4712 VSUBS 0.024813f
C3973 AVSS.n4714 VSUBS 0.011633f
C3974 AVSS.n4715 VSUBS 0.014835f
C3975 AVSS.n4716 VSUBS 0.017327f
C3976 AVSS.n4718 VSUBS 0.013464f
C3977 AVSS.n4721 VSUBS 0.01429f
C3978 AVSS.n4722 VSUBS 0.068602f
C3979 AVSS.n4723 VSUBS 0.088342f
C3980 AVSS.n4724 VSUBS 0.020848f
C3981 AVSS.n4725 VSUBS 0.013464f
C3982 AVSS.n4726 VSUBS 0.257281f
C3983 AVSS.n4727 VSUBS 0.013464f
C3984 AVSS.n4728 VSUBS 0.013197f
C3985 AVSS.n4729 VSUBS 0.013464f
C3986 AVSS.n4730 VSUBS 0.013197f
C3987 AVSS.n4731 VSUBS 0.257281f
C3988 AVSS.n4732 VSUBS 0.013464f
C3989 AVSS.n4733 VSUBS 0.021004f
C3990 AVSS.n4734 VSUBS 0.013464f
C3991 AVSS.n4735 VSUBS 0.013197f
C3992 AVSS.n4737 VSUBS 0.013464f
C3993 AVSS.n4738 VSUBS 0.013197f
C3994 AVSS.n4741 VSUBS 0.013464f
C3995 AVSS.n4742 VSUBS 0.013197f
C3996 AVSS.n4743 VSUBS 0.013197f
C3997 AVSS.n4744 VSUBS 0.013464f
C3998 AVSS.n4746 VSUBS 0.013464f
C3999 AVSS.n4747 VSUBS 0.013464f
C4000 AVSS.n4748 VSUBS 0.013197f
C4001 AVSS.n4749 VSUBS 0.013197f
C4002 AVSS.n4750 VSUBS 0.013197f
C4003 AVSS.n4751 VSUBS 0.013464f
C4004 AVSS.n4753 VSUBS 0.013464f
C4005 AVSS.n4754 VSUBS 0.013464f
C4006 AVSS.n4755 VSUBS 0.013197f
C4007 AVSS.n4756 VSUBS 0.013197f
C4008 AVSS.n4757 VSUBS 0.01932f
C4009 AVSS.n4758 VSUBS 0.019496f
C4010 AVSS.n4759 VSUBS 0.021345f
C4011 AVSS.n4760 VSUBS 0.415938f
C4012 AVSS.n4761 VSUBS 0.257281f
C4013 AVSS.n4762 VSUBS 0.013464f
C4014 AVSS.n4763 VSUBS 0.013197f
C4015 AVSS.n4764 VSUBS 0.013197f
C4016 AVSS.n4765 VSUBS 0.013197f
C4017 AVSS.n4766 VSUBS 0.013197f
C4018 AVSS.n4767 VSUBS 0.013464f
C4019 AVSS.n4768 VSUBS 0.257281f
C4020 AVSS.n4769 VSUBS 0.257281f
C4021 AVSS.n4770 VSUBS 0.190102f
C4022 AVSS.n4771 VSUBS 0.013464f
C4023 AVSS.n4772 VSUBS 0.013464f
C4024 AVSS.n4773 VSUBS 0.19582f
C4025 AVSS.n4774 VSUBS 0.257281f
C4026 AVSS.n4775 VSUBS 0.013464f
C4027 AVSS.n4776 VSUBS 0.013197f
C4028 AVSS.n4777 VSUBS 0.013197f
C4029 AVSS.n4778 VSUBS 0.013197f
C4030 AVSS.n4779 VSUBS 0.013197f
C4031 AVSS.n4780 VSUBS 0.013464f
C4032 AVSS.n4781 VSUBS 0.257281f
C4033 AVSS.n4782 VSUBS 0.257281f
C4034 AVSS.n4783 VSUBS 0.410221f
C4035 AVSS.n4784 VSUBS 0.021194f
C4036 AVSS.n4785 VSUBS 0.019048f
C4037 AVSS.n4786 VSUBS 0.018889f
C4038 AVSS.n4787 VSUBS 0.013197f
C4039 AVSS.n4788 VSUBS 0.013464f
C4040 AVSS.n4789 VSUBS 0.013464f
C4041 AVSS.n4790 VSUBS 0.013197f
C4042 AVSS.n4791 VSUBS 0.013197f
C4043 AVSS.n4792 VSUBS 0.013464f
C4044 AVSS.n4793 VSUBS 0.013464f
C4045 AVSS.n4794 VSUBS 0.013197f
C4046 AVSS.n4795 VSUBS 0.013197f
C4047 AVSS.n4796 VSUBS 0.013464f
C4048 AVSS.n4797 VSUBS 0.013464f
C4049 AVSS.n4798 VSUBS 0.013197f
C4050 AVSS.n4799 VSUBS 0.013197f
C4051 AVSS.n4800 VSUBS 0.013464f
C4052 AVSS.n4801 VSUBS 0.013464f
C4053 AVSS.n4802 VSUBS 0.013197f
C4054 AVSS.n4803 VSUBS 0.013197f
C4055 AVSS.n4804 VSUBS 0.013464f
C4056 AVSS.n4805 VSUBS 0.013464f
C4057 AVSS.n4806 VSUBS 0.010705f
C4058 AVSS.n4808 VSUBS 0.018072f
C4059 AVSS.n4809 VSUBS 0.075481f
C4060 AVSS.n4813 VSUBS 0.013002f
C4061 AVSS.n4832 VSUBS 0.015863f
C4062 AVSS.n4844 VSUBS 0.014231f
C4063 AVSS.n4845 VSUBS 0.014231f
C4064 AVSS.n4846 VSUBS 0.015203f
C4065 AVSS.n4847 VSUBS 0.015203f
C4066 AVSS.n4862 VSUBS 0.015863f
C4067 AVSS.n4877 VSUBS 0.013536f
C4068 AVSS.n4879 VSUBS 0.010931f
C4069 AVSS.n4881 VSUBS 0.014085f
C4070 AVSS.n4895 VSUBS 0.014104f
C4071 AVSS.n4896 VSUBS 0.014104f
C4072 AVSS.t93 VSUBS 1.58362f
C4073 AVSS.n4898 VSUBS 0.010886f
C4074 AVSS.n4901 VSUBS 0.075408f
C4075 AVSS.n4902 VSUBS 0.018072f
C4076 AVSS.n4905 VSUBS 0.013464f
C4077 AVSS.n4907 VSUBS 0.017327f
C4078 AVSS.n4908 VSUBS 0.014835f
C4079 AVSS.n4909 VSUBS 0.014713f
C4080 AVSS.n4910 VSUBS 0.013197f
C4081 AVSS.n4911 VSUBS 0.013464f
C4082 AVSS.n4912 VSUBS 0.013464f
C4083 AVSS.n4913 VSUBS 0.013197f
C4084 AVSS.n4914 VSUBS 0.013197f
C4085 AVSS.n4915 VSUBS 0.013464f
C4086 AVSS.n4916 VSUBS 0.013464f
C4087 AVSS.n4917 VSUBS 0.013197f
C4088 AVSS.n4918 VSUBS 0.013197f
C4089 AVSS.n4919 VSUBS 0.013464f
C4090 AVSS.n4920 VSUBS 0.013464f
C4091 AVSS.n4922 VSUBS 0.012464f
C4092 AVSS.n4923 VSUBS 0.013197f
C4093 AVSS.n4924 VSUBS 0.013464f
C4094 AVSS.n4926 VSUBS 0.135542f
C4095 AVSS.n4928 VSUBS 0.013464f
C4096 AVSS.n4929 VSUBS 0.013197f
C4097 AVSS.n4930 VSUBS 0.014549f
C4098 AVSS.n4931 VSUBS 0.016685f
C4099 AVSS.n4932 VSUBS 0.016888f
C4100 AVSS.n4933 VSUBS 0.863324f
C4101 AVSS.n4935 VSUBS 0.013464f
C4102 AVSS.n4936 VSUBS 0.013197f
C4103 AVSS.n4937 VSUBS 0.016685f
C4104 AVSS.n4938 VSUBS 0.014549f
C4105 AVSS.n4939 VSUBS 0.014676f
C4106 AVSS.n4941 VSUBS 0.013464f
C4107 AVSS.n4942 VSUBS 0.013464f
C4108 AVSS.n4943 VSUBS 0.013197f
C4109 AVSS.n4944 VSUBS 0.013197f
C4110 AVSS.n4945 VSUBS 0.012464f
C4111 AVSS.n4946 VSUBS 0.013464f
C4112 AVSS.n4948 VSUBS 0.013464f
C4113 AVSS.n4949 VSUBS 0.013464f
C4114 AVSS.n4950 VSUBS 0.013197f
C4115 AVSS.n4951 VSUBS 0.013197f
C4116 AVSS.n4952 VSUBS 0.013197f
C4117 AVSS.n4953 VSUBS 0.013464f
C4118 AVSS.n4955 VSUBS 0.013464f
C4119 AVSS.n4956 VSUBS 0.013464f
C4120 AVSS.n4957 VSUBS 0.013197f
C4121 AVSS.n4958 VSUBS 0.014713f
C4122 AVSS.n4959 VSUBS 0.017108f
C4123 AVSS.n4960 VSUBS 0.017327f
C4124 AVSS.n4962 VSUBS 0.013464f
C4125 AVSS.n4963 VSUBS 0.013464f
C4126 AVSS.n4964 VSUBS 0.013197f
C4127 AVSS.n4965 VSUBS 0.013197f
C4128 AVSS.n4966 VSUBS 0.013197f
C4129 AVSS.n4967 VSUBS 0.013464f
C4130 AVSS.n4969 VSUBS 0.013464f
C4131 AVSS.n4970 VSUBS 0.013464f
C4132 AVSS.n4971 VSUBS 0.013197f
C4133 AVSS.n4972 VSUBS 0.013197f
C4134 AVSS.n4973 VSUBS 0.013197f
C4135 AVSS.n4974 VSUBS 0.013464f
C4136 AVSS.n4976 VSUBS 0.013464f
C4137 AVSS.n4977 VSUBS 0.013464f
C4138 AVSS.n4979 VSUBS 0.013464f
C4139 AVSS.n4982 VSUBS 0.017703f
C4140 AVSS.n4983 VSUBS 0.06892f
C4141 AVSS.n4984 VSUBS 0.01429f
C4142 AVSS.n4986 VSUBS 0.017129f
C4143 AVSS.n4987 VSUBS 0.019048f
C4144 AVSS.n4988 VSUBS 0.863324f
C4145 AVSS.n4990 VSUBS 0.013464f
C4146 AVSS.n4992 VSUBS 0.016685f
C4147 AVSS.n4993 VSUBS 0.011763f
C4148 AVSS.n4994 VSUBS 0.014676f
C4149 AVSS.n4996 VSUBS 0.013464f
C4150 AVSS.n4997 VSUBS 0.013464f
C4151 AVSS.n4998 VSUBS 0.013197f
C4152 AVSS.n4999 VSUBS 0.013197f
C4153 AVSS.n5000 VSUBS 0.012464f
C4154 AVSS.n5001 VSUBS 0.013464f
C4155 AVSS.n5003 VSUBS 0.013464f
C4156 AVSS.n5004 VSUBS 0.013464f
C4157 AVSS.n5005 VSUBS 0.013197f
C4158 AVSS.n5006 VSUBS 0.013197f
C4159 AVSS.n5007 VSUBS 0.013197f
C4160 AVSS.n5008 VSUBS 0.013464f
C4161 AVSS.n5010 VSUBS 0.013464f
C4162 AVSS.n5011 VSUBS 0.013464f
C4163 AVSS.n5012 VSUBS 0.013197f
C4164 AVSS.n5013 VSUBS 0.014713f
C4165 AVSS.n5014 VSUBS 0.017108f
C4166 AVSS.n5015 VSUBS 0.017327f
C4167 AVSS.n5016 VSUBS 0.863324f
C4168 AVSS.n5017 VSUBS 0.051397f
C4169 AVSS.n5018 VSUBS 0.045828f
C4170 AVSS.n5019 VSUBS 0.04266f
C4171 AVSS.n5020 VSUBS 0.205814f
C4172 AVSS.n5021 VSUBS 0.093787f
C4173 AVSS.n5022 VSUBS 0.165515f
C4174 AVSS.n5024 VSUBS 0.0905f
C4175 AVSS.n5025 VSUBS 0.160158f
C4176 AVSS.n5026 VSUBS 0.143448f
C4177 AVSS.n5027 VSUBS 0.112183f
C4178 AVSS.n5028 VSUBS 0.097957f
C4179 AVSS.n5029 VSUBS 0.160845f
C4180 AVSS.n5030 VSUBS 0.084482f
C4181 AVSS.n5031 VSUBS 0.205976f
C4182 AVSS.n5032 VSUBS 0.051397f
C4183 AVSS.n5033 VSUBS 0.046257f
C4184 AVSS.n5034 VSUBS 0.036742f
C4185 AVSS.n5035 VSUBS 0.045176f
C4186 AVSS.n5036 VSUBS 0.033466f
C4187 AVSS.n5037 VSUBS 0.030324f
C4188 AVSS.n5038 VSUBS 0.04266f
C4189 AVSS.n5039 VSUBS 0.067428f
C4190 AVSS.n5040 VSUBS 0.093787f
C4191 AVSS.n5041 VSUBS 0.166175f
C4192 AVSS.n5042 VSUBS 0.089157f
C4193 AVSS.n5043 VSUBS 0.115853f
C4194 AVSS.n5044 VSUBS 0.186488f
C4195 AVSS.n5045 VSUBS 0.189601f
C4196 AVSS.n5046 VSUBS 0.051397f
C4197 AVSS.n5047 VSUBS 0.077272f
C4198 AVSS.n5048 VSUBS 0.090352f
C4199 AVSS.n5049 VSUBS 0.090352f
C4200 AVSS.n5050 VSUBS 0.090352f
C4201 AVSS.n5051 VSUBS 0.051397f
C4202 AVSS.n5052 VSUBS 0.077272f
C4203 AVSS.n5053 VSUBS 0.189601f
C4204 AVSS.n5054 VSUBS 0.186488f
C4205 AVSS.n5055 VSUBS 0.114153f
C4206 AVSS.n5056 VSUBS 0.192018f
C4207 AVSS.n5057 VSUBS 0.04266f
C4208 AVSS.n5058 VSUBS 0.210564f
C4209 AVSS.n5059 VSUBS 0.067428f
C4210 AVSS.n5060 VSUBS 0.090352f
C4211 AVSS.n5061 VSUBS 0.090352f
C4212 AVSS.n5062 VSUBS 0.030324f
C4213 AVSS.n5063 VSUBS 0.051397f
C4214 AVSS.n5064 VSUBS 0.045828f
C4215 AVSS.t99 VSUBS 0.154434f
C4216 AVSS.n5065 VSUBS 0.183064f
C4217 AVSS.n5066 VSUBS 0.013464f
C4218 AVSS.n5067 VSUBS 0.013197f
C4219 AVSS.n5068 VSUBS 0.013197f
C4220 AVSS.n5069 VSUBS 0.013197f
C4221 AVSS.n5070 VSUBS 0.013464f
C4222 AVSS.n5071 VSUBS 0.218223f
C4223 AVSS.n5072 VSUBS 0.218223f
C4224 AVSS.n5073 VSUBS 0.218223f
C4225 AVSS.n5074 VSUBS 0.013464f
C4226 AVSS.n5075 VSUBS 0.013197f
C4227 AVSS.n5076 VSUBS 0.01932f
C4228 AVSS.n5077 VSUBS 0.013197f
C4229 AVSS.n5078 VSUBS 0.013464f
C4230 AVSS.n5079 VSUBS 0.013464f
C4231 AVSS.n5080 VSUBS 0.013197f
C4232 AVSS.n5081 VSUBS 0.013197f
C4233 AVSS.n5082 VSUBS 0.013464f
C4234 AVSS.n5083 VSUBS 0.013464f
C4235 AVSS.n5084 VSUBS 0.013197f
C4236 AVSS.n5085 VSUBS 0.013197f
C4237 AVSS.n5086 VSUBS 0.013464f
C4238 AVSS.n5087 VSUBS 0.013464f
C4239 AVSS.n5088 VSUBS 0.013197f
C4240 AVSS.n5089 VSUBS 0.013464f
C4241 AVSS.n5090 VSUBS 0.013197f
C4242 AVSS.n5091 VSUBS 0.013197f
C4243 AVSS.n5092 VSUBS 0.021004f
C4244 AVSS.n5093 VSUBS 0.021345f
C4245 AVSS.n5095 VSUBS 0.135542f
C4246 AVSS.n5097 VSUBS 0.013464f
C4247 AVSS.n5100 VSUBS 0.018072f
C4248 AVSS.n5101 VSUBS 0.075408f
C4249 AVSS.n5104 VSUBS 0.013536f
C4250 AVSS.t98 VSUBS 1.58362f
C4251 AVSS.n5108 VSUBS 0.014104f
C4252 AVSS.n5113 VSUBS 0.014231f
C4253 AVSS.n5117 VSUBS 0.010886f
C4254 AVSS.n5136 VSUBS 0.013002f
C4255 AVSS.n5137 VSUBS 0.013002f
C4256 AVSS.n5139 VSUBS 0.010886f
C4257 AVSS.n5155 VSUBS 0.014231f
C4258 AVSS.n5157 VSUBS 0.015203f
C4259 AVSS.n5158 VSUBS 0.015203f
C4260 AVSS.n5173 VSUBS 0.015863f
C4261 AVSS.n5175 VSUBS 0.012104f
C4262 AVSS.n5176 VSUBS 0.010825f
C4263 AVSS.n5191 VSUBS 0.014085f
C4264 AVSS.n5193 VSUBS 0.010931f
C4265 AVSS.n5194 VSUBS 0.075481f
C4266 AVSS.n5195 VSUBS 0.018072f
C4267 AVSS.n5198 VSUBS 0.013464f
C4268 AVSS.n5199 VSUBS 0.013197f
C4269 AVSS.n5200 VSUBS 0.013197f
C4270 AVSS.n5201 VSUBS 0.013464f
C4271 AVSS.n5202 VSUBS 0.013464f
C4272 AVSS.n5203 VSUBS 0.012464f
C4273 AVSS.n5205 VSUBS 0.013464f
C4274 AVSS.n5206 VSUBS 0.013464f
C4275 AVSS.n5207 VSUBS 0.013197f
C4276 AVSS.n5208 VSUBS 0.013197f
C4277 AVSS.n5209 VSUBS 0.013464f
C4278 AVSS.n5210 VSUBS 0.013464f
C4279 AVSS.n5211 VSUBS 0.013197f
C4280 AVSS.n5212 VSUBS 0.013197f
C4281 AVSS.n5213 VSUBS 0.013464f
C4282 AVSS.n5214 VSUBS 0.013464f
C4283 AVSS.n5215 VSUBS 0.013197f
C4284 AVSS.n5216 VSUBS 0.014713f
C4285 AVSS.n5217 VSUBS 0.017108f
C4286 AVSS.n5218 VSUBS 0.017327f
C4287 AVSS.n5219 VSUBS 0.260654f
C4288 AVSS.n5220 VSUBS 0.527322f
C4289 AVSS.n5221 VSUBS 0.135542f
C4290 AVSS.n5223 VSUBS 0.014676f
C4291 AVSS.n5224 VSUBS 0.016888f
C4292 AVSS.n5225 VSUBS 0.016685f
C4293 AVSS.n5226 VSUBS 0.013197f
C4294 AVSS.n5227 VSUBS 0.013464f
C4295 AVSS.n5228 VSUBS 0.013464f
C4296 AVSS.n5229 VSUBS 0.013197f
C4297 AVSS.n5230 VSUBS 0.013197f
C4298 AVSS.n5231 VSUBS 0.013464f
C4299 AVSS.n5232 VSUBS 0.013464f
C4300 AVSS.n5233 VSUBS 0.013197f
C4301 AVSS.n5234 VSUBS 0.013197f
C4302 AVSS.n5235 VSUBS 0.013464f
C4303 AVSS.n5236 VSUBS 0.013464f
C4304 AVSS.n5237 VSUBS 0.013197f
C4305 AVSS.n5238 VSUBS 0.013197f
C4306 AVSS.n5239 VSUBS 0.013464f
C4307 AVSS.n5240 VSUBS 0.013464f
C4308 AVSS.n5241 VSUBS 0.013197f
C4309 AVSS.n5242 VSUBS 0.013197f
C4310 AVSS.n5243 VSUBS 0.013464f
C4311 AVSS.n5244 VSUBS 0.013464f
C4312 AVSS.n5245 VSUBS 0.013197f
C4313 AVSS.n5246 VSUBS 0.013197f
C4314 AVSS.n5247 VSUBS 0.018889f
C4315 AVSS.n5248 VSUBS 0.019048f
C4316 AVSS.n5255 VSUBS 0.021194f
C4317 AVSS.n5256 VSUBS 0.013464f
C4318 AVSS.n5257 VSUBS 0.018062f
C4319 AVSS.n5258 VSUBS 0.014549f
C4320 AVSS.n5259 VSUBS 0.013464f
C4321 AVSS.n5265 VSUBS 0.218223f
C4322 AVSS.n5266 VSUBS 0.013464f
C4323 AVSS.n5267 VSUBS 0.014835f
C4324 AVSS.n5268 VSUBS 0.013197f
C4325 AVSS.n5269 VSUBS 0.013464f
C4326 AVSS.n5270 VSUBS 0.218223f
C4327 AVSS.n5271 VSUBS 0.013464f
C4328 AVSS.n5272 VSUBS 0.013197f
C4329 AVSS.n5273 VSUBS 0.013464f
C4330 AVSS.n5274 VSUBS 0.218223f
C4331 AVSS.n5275 VSUBS 0.013464f
C4332 AVSS.n5276 VSUBS 0.013197f
C4333 AVSS.n5277 VSUBS 0.013464f
C4334 AVSS.n5278 VSUBS 0.135542f
C4335 AVSS.n5279 VSUBS 0.218223f
C4336 AVSS.n5280 VSUBS 0.013464f
C4337 AVSS.n5281 VSUBS 0.014835f
C4338 AVSS.n5282 VSUBS 0.013197f
C4339 AVSS.n5283 VSUBS 0.013464f
C4340 AVSS.n5284 VSUBS 0.218223f
C4341 AVSS.n5285 VSUBS 0.013464f
C4342 AVSS.n5286 VSUBS 0.013197f
C4343 AVSS.n5287 VSUBS 0.013197f
C4344 AVSS.n5288 VSUBS 0.013464f
C4345 AVSS.n5289 VSUBS 0.218223f
C4346 AVSS.n5290 VSUBS 0.218223f
C4347 AVSS.n5291 VSUBS 0.218223f
C4348 AVSS.n5292 VSUBS 0.013464f
C4349 AVSS.n5293 VSUBS 0.013197f
C4350 AVSS.n5294 VSUBS 0.013197f
C4351 AVSS.n5295 VSUBS 0.013197f
C4352 AVSS.n5296 VSUBS 0.013464f
C4353 AVSS.n5298 VSUBS 0.013464f
C4354 AVSS.n5300 VSUBS 0.016888f
C4355 AVSS.n5303 VSUBS 0.013536f
C4356 AVSS.t88 VSUBS 1.58362f
C4357 AVSS.n5307 VSUBS 0.014104f
C4358 AVSS.n5312 VSUBS 0.014231f
C4359 AVSS.n5316 VSUBS 0.010886f
C4360 AVSS.n5335 VSUBS 0.013002f
C4361 AVSS.n5336 VSUBS 0.013002f
C4362 AVSS.n5338 VSUBS 0.010886f
C4363 AVSS.n5354 VSUBS 0.014231f
C4364 AVSS.n5356 VSUBS 0.015203f
C4365 AVSS.n5357 VSUBS 0.015203f
C4366 AVSS.n5372 VSUBS 0.015863f
C4367 AVSS.n5374 VSUBS 0.012104f
C4368 AVSS.n5375 VSUBS 0.010825f
C4369 AVSS.n5390 VSUBS 0.014085f
C4370 AVSS.n5392 VSUBS 0.010931f
C4371 AVSS.n5393 VSUBS 0.075481f
C4372 AVSS.n5394 VSUBS 0.018072f
C4373 AVSS.n5396 VSUBS 0.013464f
C4374 AVSS.n5397 VSUBS 0.013197f
C4375 AVSS.n5398 VSUBS 0.013197f
C4376 AVSS.n5399 VSUBS 0.013464f
C4377 AVSS.n5400 VSUBS 0.013464f
C4378 AVSS.n5401 VSUBS 0.013197f
C4379 AVSS.n5402 VSUBS 0.013197f
C4380 AVSS.n5403 VSUBS 0.013464f
C4381 AVSS.n5404 VSUBS 0.013464f
C4382 AVSS.n5405 VSUBS 0.013197f
C4383 AVSS.n5406 VSUBS 0.013197f
C4384 AVSS.n5407 VSUBS 0.013464f
C4385 AVSS.n5408 VSUBS 0.013464f
C4386 AVSS.n5409 VSUBS 0.013197f
C4387 AVSS.n5410 VSUBS 0.013197f
C4388 AVSS.n5411 VSUBS 0.013464f
C4389 AVSS.n5412 VSUBS 0.013464f
C4390 AVSS.n5413 VSUBS 0.013197f
C4391 AVSS.n5414 VSUBS 0.013197f
C4392 AVSS.n5415 VSUBS 0.013464f
C4393 AVSS.n5416 VSUBS 0.013464f
C4394 AVSS.n5417 VSUBS 0.013197f
C4395 AVSS.n5418 VSUBS 0.016685f
C4396 AVSS.n5419 VSUBS 0.011763f
C4397 AVSS.n5420 VSUBS 0.014676f
C4398 AVSS.n5422 VSUBS 0.013464f
C4399 AVSS.n5424 VSUBS 0.013464f
C4400 AVSS.n5425 VSUBS 0.013197f
C4401 AVSS.n5426 VSUBS 0.013197f
C4402 AVSS.n5427 VSUBS 0.012464f
C4403 AVSS.n5428 VSUBS 0.013464f
C4404 AVSS.n5430 VSUBS 0.013464f
C4405 AVSS.n5432 VSUBS 0.013464f
C4406 AVSS.n5433 VSUBS 0.013197f
C4407 AVSS.n5434 VSUBS 0.013197f
C4408 AVSS.n5435 VSUBS 0.013197f
C4409 AVSS.n5436 VSUBS 0.013464f
C4410 AVSS.n5438 VSUBS 0.013464f
C4411 AVSS.n5440 VSUBS 0.013464f
C4412 AVSS.n5441 VSUBS 0.013197f
C4413 AVSS.n5442 VSUBS 0.014713f
C4414 AVSS.n5443 VSUBS 0.017108f
C4415 AVSS.n5444 VSUBS 0.017327f
C4416 AVSS.n5445 VSUBS 0.260654f
C4417 AVSS.n5446 VSUBS 0.527322f
C4418 AVSS.n5447 VSUBS 0.021345f
C4419 AVSS.n5448 VSUBS 0.013197f
C4420 AVSS.n5449 VSUBS 0.013464f
C4421 AVSS.n5454 VSUBS 0.013464f
C4422 AVSS.n5474 VSUBS 0.015203f
C4423 AVSS.n5487 VSUBS 0.014085f
C4424 AVSS.n5488 VSUBS 0.014085f
C4425 AVSS.n5489 VSUBS 0.013536f
C4426 AVSS.n5490 VSUBS 0.013536f
C4427 AVSS.n5505 VSUBS 0.013002f
C4428 AVSS.n5506 VSUBS 0.013002f
C4429 AVSS.n5507 VSUBS 0.010886f
C4430 AVSS.n5508 VSUBS 0.010886f
C4431 AVSS.n5523 VSUBS 0.014231f
C4432 AVSS.n5524 VSUBS 0.014231f
C4433 AVSS.n5525 VSUBS 0.015203f
C4434 AVSS.n5526 VSUBS 0.015863f
C4435 AVSS.t91 VSUBS 1.58362f
C4436 AVSS.n5543 VSUBS 0.014104f
C4437 AVSS.n5544 VSUBS 0.010825f
C4438 AVSS.n5545 VSUBS 0.012104f
C4439 AVSS.n5546 VSUBS 0.09348f
C4440 AVSS.n5547 VSUBS 0.018072f
C4441 AVSS.n5550 VSUBS 0.013464f
C4442 AVSS.n5551 VSUBS 0.013464f
C4443 AVSS.n5552 VSUBS 0.013197f
C4444 AVSS.n5553 VSUBS 0.013197f
C4445 AVSS.n5554 VSUBS 0.013464f
C4446 AVSS.n5555 VSUBS 0.013464f
C4447 AVSS.n5556 VSUBS 0.013197f
C4448 AVSS.n5557 VSUBS 0.013197f
C4449 AVSS.n5558 VSUBS 0.013464f
C4450 AVSS.n5559 VSUBS 0.013464f
C4451 AVSS.n5560 VSUBS 0.013197f
C4452 AVSS.n5561 VSUBS 0.013197f
C4453 AVSS.n5562 VSUBS 0.013197f
C4454 AVSS.n5563 VSUBS 0.013464f
C4455 AVSS.n5565 VSUBS 0.135542f
C4456 AVSS.n5567 VSUBS 0.013464f
C4457 AVSS.n5568 VSUBS 0.013197f
C4458 AVSS.n5569 VSUBS 0.021004f
C4459 AVSS.n5570 VSUBS 0.01932f
C4460 AVSS.n5571 VSUBS 0.019496f
C4461 AVSS.n5572 VSUBS 0.33097f
C4462 AVSS.n5573 VSUBS 0.218223f
C4463 AVSS.n5574 VSUBS 0.218223f
C4464 AVSS.n5575 VSUBS 0.013464f
C4465 AVSS.n5576 VSUBS 0.013197f
C4466 AVSS.n5577 VSUBS 0.013197f
C4467 AVSS.n5578 VSUBS 0.013197f
C4468 AVSS.n5579 VSUBS 0.013464f
C4469 AVSS.n5580 VSUBS 0.218223f
C4470 AVSS.n5581 VSUBS 0.183064f
C4471 AVSS.t92 VSUBS 0.154434f
C4472 AVSS.n5582 VSUBS 0.144269f
C4473 AVSS.n5583 VSUBS 0.013464f
C4474 AVSS.n5584 VSUBS 0.013197f
C4475 AVSS.n5585 VSUBS 0.013197f
C4476 AVSS.n5586 VSUBS 0.013197f
C4477 AVSS.n5587 VSUBS 0.013464f
C4478 AVSS.n5588 VSUBS 0.218223f
C4479 AVSS.n5589 VSUBS 0.218223f
C4480 AVSS.n5590 VSUBS 0.218223f
C4481 AVSS.n5591 VSUBS 0.013464f
C4482 AVSS.n5592 VSUBS 0.013197f
C4483 AVSS.n5593 VSUBS 0.013197f
C4484 AVSS.n5594 VSUBS 0.013197f
C4485 AVSS.n5595 VSUBS 0.013464f
C4486 AVSS.n5596 VSUBS 0.013197f
C4487 AVSS.n5597 VSUBS 0.013197f
C4488 AVSS.n5598 VSUBS 0.013464f
C4489 AVSS.n5599 VSUBS 0.013464f
C4490 AVSS.n5600 VSUBS 0.012464f
C4491 AVSS.n5602 VSUBS 0.013464f
C4492 AVSS.n5603 VSUBS 0.013464f
C4493 AVSS.n5604 VSUBS 0.013197f
C4494 AVSS.n5605 VSUBS 0.013197f
C4495 AVSS.n5606 VSUBS 0.013464f
C4496 AVSS.n5607 VSUBS 0.013464f
C4497 AVSS.n5608 VSUBS 0.013197f
C4498 AVSS.n5609 VSUBS 0.013197f
C4499 AVSS.n5610 VSUBS 0.013464f
C4500 AVSS.n5611 VSUBS 0.013464f
C4501 AVSS.n5612 VSUBS 0.013197f
C4502 AVSS.n5613 VSUBS 0.014713f
C4503 AVSS.n5614 VSUBS 0.017108f
C4504 AVSS.n5615 VSUBS 0.017327f
C4505 AVSS.n5616 VSUBS 0.260654f
C4506 AVSS.n5617 VSUBS 0.33097f
C4507 AVSS.n5623 VSUBS 0.013464f
C4508 AVSS.n5624 VSUBS 0.019496f
C4509 AVSS.n5625 VSUBS 0.01932f
C4510 AVSS.n5626 VSUBS 0.018062f
C4511 AVSS.n5627 VSUBS 0.021194f
C4512 AVSS.n5628 VSUBS 0.019048f
C4513 AVSS.n5629 VSUBS 0.017129f
C4514 AVSS.n5630 VSUBS 0.016685f
C4515 AVSS.n5631 VSUBS 0.014676f
C4516 AVSS.n5632 VSUBS 0.027461f
C4517 AVSS.n5633 VSUBS 0.013464f
C4518 AVSS.n5634 VSUBS 0.012464f
C4519 AVSS.n5635 VSUBS 0.013464f
C4520 AVSS.n5636 VSUBS 0.013464f
C4521 AVSS.n5637 VSUBS 0.013197f
C4522 AVSS.n5638 VSUBS 0.013464f
C4523 AVSS.n5639 VSUBS 0.027461f
C4524 AVSS.n5640 VSUBS 0.013464f
C4525 AVSS.n5641 VSUBS 0.017108f
C4526 AVSS.n5642 VSUBS 0.017327f
C4527 AVSS.n5643 VSUBS 0.218223f
C4528 AVSS.n5644 VSUBS 0.013464f
C4529 AVSS.n5645 VSUBS 0.013197f
C4530 AVSS.n5646 VSUBS 0.013464f
C4531 AVSS.n5647 VSUBS 0.013464f
C4532 AVSS.n5648 VSUBS 0.013197f
C4533 AVSS.n5649 VSUBS 0.013464f
C4534 AVSS.n5650 VSUBS 0.218223f
C4535 AVSS.n5651 VSUBS 0.013464f
C4536 AVSS.n5652 VSUBS 0.013197f
C4537 AVSS.n5653 VSUBS 0.013197f
C4538 AVSS.n5654 VSUBS 0.013197f
C4539 AVSS.n5655 VSUBS 0.013464f
C4540 AVSS.n5656 VSUBS 0.218223f
C4541 AVSS.n5657 VSUBS 0.218223f
C4542 AVSS.n5658 VSUBS 0.218223f
C4543 AVSS.n5659 VSUBS 0.013464f
C4544 AVSS.n5660 VSUBS 0.013464f
C4545 AVSS.n5661 VSUBS 0.013197f
C4546 AVSS.n5662 VSUBS 0.013197f
C4547 AVSS.n5663 VSUBS 0.013197f
C4548 AVSS.n5664 VSUBS 0.013464f
C4549 AVSS.n5665 VSUBS 0.218223f
C4550 AVSS.n5666 VSUBS 0.218223f
C4551 AVSS.n5667 VSUBS 0.218223f
C4552 AVSS.n5668 VSUBS 0.013464f
C4553 AVSS.n5669 VSUBS 0.013197f
C4554 AVSS.n5670 VSUBS 0.013197f
C4555 AVSS.n5671 VSUBS 0.013197f
C4556 AVSS.n5672 VSUBS 0.013464f
C4557 AVSS.n5673 VSUBS 0.561572f
C4558 AVSS.n5674 VSUBS 0.13108f
C4559 AVSS.n5675 VSUBS 0.029139f
C4560 AVSS.n5676 VSUBS 0.014835f
C4561 AVSS.n5677 VSUBS 0.014713f
C4562 AVSS.n5678 VSUBS 0.013197f
C4563 AVSS.n5679 VSUBS 0.013197f
C4564 AVSS.n5680 VSUBS 0.013464f
C4565 AVSS.n5681 VSUBS 0.027461f
C4566 AVSS.n5682 VSUBS 0.027461f
C4567 AVSS.n5683 VSUBS 0.020291f
C4568 AVSS.n5684 VSUBS 0.027461f
C4569 AVSS.n5685 VSUBS 0.013464f
C4570 AVSS.n5686 VSUBS 0.013197f
C4571 AVSS.n5687 VSUBS 0.013197f
C4572 AVSS.n5689 VSUBS 0.013464f
C4573 AVSS.n5690 VSUBS 0.020901f
C4574 AVSS.n5691 VSUBS 0.027461f
C4575 AVSS.n5692 VSUBS 0.027461f
C4576 AVSS.n5693 VSUBS 0.013464f
C4577 AVSS.n5694 VSUBS 0.013197f
C4578 AVSS.n5695 VSUBS 0.013197f
C4579 AVSS.n5696 VSUBS 0.014549f
C4580 AVSS.n5697 VSUBS 0.013197f
C4581 AVSS.n5698 VSUBS 0.013464f
C4582 AVSS.n5699 VSUBS 0.027461f
C4583 AVSS.n5700 VSUBS 0.028377f
C4584 AVSS.n5701 VSUBS 0.030055f
C4585 AVSS.n5702 VSUBS 0.016888f
C4586 AVSS.n5703 VSUBS 0.013464f
C4587 AVSS.n5704 VSUBS 0.013197f
C4588 AVSS.n5705 VSUBS 0.013197f
C4589 AVSS.n5706 VSUBS 0.013464f
C4590 AVSS.n5707 VSUBS 0.013464f
C4591 AVSS.n5708 VSUBS 0.013197f
C4592 AVSS.n5709 VSUBS 0.013197f
C4593 AVSS.n5710 VSUBS 0.013464f
C4594 AVSS.n5711 VSUBS 0.013464f
C4595 AVSS.n5712 VSUBS 0.013197f
C4596 AVSS.n5713 VSUBS 0.013197f
C4597 AVSS.n5714 VSUBS 0.013464f
C4598 AVSS.n5715 VSUBS 0.013464f
C4599 AVSS.n5716 VSUBS 0.013197f
C4600 AVSS.n5717 VSUBS 0.013197f
C4601 AVSS.n5718 VSUBS 0.013464f
C4602 AVSS.n5719 VSUBS 0.013464f
C4603 AVSS.n5720 VSUBS 0.013197f
C4604 AVSS.n5721 VSUBS 0.013197f
C4605 AVSS.n5722 VSUBS 0.013464f
C4606 AVSS.n5723 VSUBS 0.013464f
C4607 AVSS.n5726 VSUBS 0.014516f
C4608 AVSS.n5746 VSUBS 0.015203f
C4609 AVSS.n5759 VSUBS 0.014085f
C4610 AVSS.n5760 VSUBS 0.014085f
C4611 AVSS.n5761 VSUBS 0.013536f
C4612 AVSS.n5762 VSUBS 0.013536f
C4613 AVSS.n5777 VSUBS 0.013002f
C4614 AVSS.n5778 VSUBS 0.013002f
C4615 AVSS.n5779 VSUBS 0.010886f
C4616 AVSS.n5780 VSUBS 0.010886f
C4617 AVSS.n5795 VSUBS 0.014231f
C4618 AVSS.n5796 VSUBS 0.014231f
C4619 AVSS.n5797 VSUBS 0.015203f
C4620 AVSS.n5798 VSUBS 0.015863f
C4621 AVSS.t105 VSUBS 1.58362f
C4622 AVSS.n5815 VSUBS 0.014104f
C4623 AVSS.n5816 VSUBS 0.010825f
C4624 AVSS.n5817 VSUBS 0.012104f
C4625 AVSS.n5818 VSUBS 0.025257f
C4626 AVSS.n5819 VSUBS 0.018072f
C4627 AVSS.n5822 VSUBS 0.013464f
C4628 AVSS.n5823 VSUBS 0.013464f
C4629 AVSS.n5824 VSUBS 0.013197f
C4630 AVSS.n5825 VSUBS 0.013197f
C4631 AVSS.n5826 VSUBS 0.013464f
C4632 AVSS.n5827 VSUBS 0.013464f
C4633 AVSS.n5828 VSUBS 0.013197f
C4634 AVSS.n5829 VSUBS 0.013197f
C4635 AVSS.n5830 VSUBS 0.013464f
C4636 AVSS.n5831 VSUBS 0.013464f
C4637 AVSS.n5832 VSUBS 0.013197f
C4638 AVSS.n5833 VSUBS 0.013197f
C4639 AVSS.n5834 VSUBS 0.013464f
C4640 AVSS.n5835 VSUBS 0.013464f
C4641 AVSS.n5836 VSUBS 0.013197f
C4642 AVSS.n5837 VSUBS 0.013464f
C4643 AVSS.n5838 VSUBS 0.013197f
C4644 AVSS.n5839 VSUBS 0.013197f
C4645 AVSS.n5840 VSUBS 0.021004f
C4646 AVSS.n5841 VSUBS 0.021345f
C4647 AVSS.n5843 VSUBS 0.135542f
C4648 AVSS.n5844 VSUBS 0.527322f
C4649 AVSS.n5845 VSUBS 0.135542f
C4650 AVSS.n5847 VSUBS 0.014676f
C4651 AVSS.n5848 VSUBS 0.016888f
C4652 AVSS.n5849 VSUBS 0.016685f
C4653 AVSS.n5850 VSUBS 0.013197f
C4654 AVSS.n5851 VSUBS 0.013464f
C4655 AVSS.n5852 VSUBS 0.013464f
C4656 AVSS.n5853 VSUBS 0.013197f
C4657 AVSS.n5854 VSUBS 0.013197f
C4658 AVSS.n5855 VSUBS 0.013464f
C4659 AVSS.n5856 VSUBS 0.013464f
C4660 AVSS.n5857 VSUBS 0.013197f
C4661 AVSS.n5858 VSUBS 0.013197f
C4662 AVSS.n5859 VSUBS 0.013464f
C4663 AVSS.n5860 VSUBS 0.013464f
C4664 AVSS.n5861 VSUBS 0.013197f
C4665 AVSS.n5862 VSUBS 0.013197f
C4666 AVSS.n5863 VSUBS 0.013464f
C4667 AVSS.n5864 VSUBS 0.013464f
C4668 AVSS.n5865 VSUBS 0.013197f
C4669 AVSS.n5866 VSUBS 0.013197f
C4670 AVSS.n5867 VSUBS 0.013464f
C4671 AVSS.n5868 VSUBS 0.013464f
C4672 AVSS.n5869 VSUBS 0.013197f
C4673 AVSS.n5870 VSUBS 0.013197f
C4674 AVSS.n5871 VSUBS 0.018889f
C4675 AVSS.n5872 VSUBS 0.019048f
C4676 AVSS.n5873 VSUBS 0.863324f
C4677 AVSS.n5875 VSUBS 0.013464f
C4678 AVSS.n5877 VSUBS 0.016685f
C4679 AVSS.n5878 VSUBS 0.011763f
C4680 AVSS.n5879 VSUBS 0.014676f
C4681 AVSS.n5881 VSUBS 0.013464f
C4682 AVSS.n5882 VSUBS 0.013464f
C4683 AVSS.n5883 VSUBS 0.013197f
C4684 AVSS.n5884 VSUBS 0.013197f
C4685 AVSS.n5885 VSUBS 0.012464f
C4686 AVSS.n5886 VSUBS 0.013464f
C4687 AVSS.n5888 VSUBS 0.013464f
C4688 AVSS.n5889 VSUBS 0.013464f
C4689 AVSS.n5890 VSUBS 0.013197f
C4690 AVSS.n5891 VSUBS 0.013197f
C4691 AVSS.n5892 VSUBS 0.013197f
C4692 AVSS.n5893 VSUBS 0.013464f
C4693 AVSS.n5895 VSUBS 0.013464f
C4694 AVSS.n5896 VSUBS 0.013464f
C4695 AVSS.n5897 VSUBS 0.013197f
C4696 AVSS.n5898 VSUBS 0.014713f
C4697 AVSS.n5899 VSUBS 0.017108f
C4698 AVSS.n5900 VSUBS 0.017327f
C4699 AVSS.n5901 VSUBS 0.260654f
C4700 AVSS.n5902 VSUBS 0.218223f
C4701 AVSS.n5903 VSUBS 0.218223f
C4702 AVSS.n5904 VSUBS 0.013464f
C4703 AVSS.n5905 VSUBS 0.013197f
C4704 AVSS.n5906 VSUBS 0.013197f
C4705 AVSS.n5907 VSUBS 0.013197f
C4706 AVSS.n5908 VSUBS 0.013464f
C4707 AVSS.n5909 VSUBS 0.218223f
C4708 AVSS.n5910 VSUBS 0.216542f
C4709 AVSS.n5911 VSUBS 0.437806f
C4710 AVSS.n5912 VSUBS 0.015125f
C4711 AVSS.n5913 VSUBS 0.013197f
C4712 AVSS.n5914 VSUBS 0.013197f
C4713 AVSS.n5915 VSUBS 0.013197f
C4714 AVSS.n5916 VSUBS 0.013464f
C4715 AVSS.n5917 VSUBS 0.582149f
C4716 AVSS.n5918 VSUBS 0.582149f
C4717 AVSS.n5919 VSUBS 0.582149f
C4718 AVSS.n5920 VSUBS 0.013464f
C4719 AVSS.n5921 VSUBS 0.013197f
C4720 AVSS.n5922 VSUBS 0.013197f
C4721 AVSS.n5923 VSUBS 0.01932f
C4722 AVSS.n5924 VSUBS 0.019496f
C4723 AVSS.n5925 VSUBS 2.48707f
C4724 AVSS.n5926 VSUBS 10.6675f
C4725 AVSS.n5927 VSUBS 35.083103f
C4726 AVSS.n5928 VSUBS 7.06384f
C4727 AVSS.t51 VSUBS 0.591947f
C4728 AVSS.n5929 VSUBS 0.123915f
C4729 AVSS.n5930 VSUBS 0.123915f
C4730 AVSS.n5931 VSUBS 0.123915f
C4731 AVSS.n5932 VSUBS 0.015244f
C4732 AVSS.n5933 VSUBS 0.124865f
C4733 AVSS.n5934 VSUBS 0.094775f
C4734 AVSS.n5935 VSUBS 0.180628f
C4735 AVSS.n5936 VSUBS 0.264405f
C4736 AVSS.n5937 VSUBS 0.263848f
C4737 AVSS.n5938 VSUBS 0.264962f
C4738 AVSS.n5939 VSUBS 0.263848f
C4739 AVSS.n5940 VSUBS 0.494478f
C4740 AVSS.t37 VSUBS 0.789263f
C4741 AVSS.t123 VSUBS 1.54524f
C4742 AVSS.t117 VSUBS 6.18255f
C4743 AVSS.t0 VSUBS 0.52776f
C4744 AVSS.n5941 VSUBS 1.28374f
C4745 AVSS.n5942 VSUBS 0.368481f
C4746 AVSS.n5943 VSUBS 0.04236f
C4747 AVSS.n5944 VSUBS 0.042102f
C4748 AVSS.n5945 VSUBS 0.042231f
C4749 AVSS.n5946 VSUBS 0.057377f
C4750 AVSS.n5947 VSUBS 0.042374f
C4751 AVSS.n5948 VSUBS 0.02119f
C4752 AVSS.n5950 VSUBS 0.02766f
C4753 AVSS.n5952 VSUBS 0.026467f
C4754 AVSS.n5953 VSUBS 0.058281f
C4755 AVSS.n5954 VSUBS 0.021313f
C4756 AVSS.n5955 VSUBS 0.057377f
C4757 AVSS.n5956 VSUBS 0.064447f
C4758 AVSS.n5957 VSUBS 0.042102f
C4759 AVSS.n5958 VSUBS 0.042374f
C4760 AVSS.n5959 VSUBS 0.042374f
C4761 AVSS.n5960 VSUBS 0.380368f
C4762 AVSS.t2 VSUBS 0.397009f
C4763 AVSS.n5961 VSUBS 0.869732f
C4764 AVSS.n5962 VSUBS 0.435726f
C4765 AVSS.n5963 VSUBS 0.435726f
C4766 AVSS.t46 VSUBS 2.71296f
C4767 AVSS.t9 VSUBS 14.997199f
C4768 AVSS.n5964 VSUBS 0.018977f
C4769 AVSS.n5965 VSUBS 0.70359f
C4770 AVSS.n5966 VSUBS 16.3579f
C4771 AVSS.t6 VSUBS 5.16465f
C4772 AVSS.t13 VSUBS 8.17894f
C4773 AVSS.n5967 VSUBS 0.705111f
C4774 AVSS.n5968 VSUBS 0.705111f
C4775 AVSS.n5969 VSUBS 0.89831f
C4776 AVSS.t18 VSUBS 0.017275f
C4777 AVSS.n5970 VSUBS 0.590814f
C4778 AVSS.t129 VSUBS 0.017275f
C4779 AVSS.n5971 VSUBS 0.143355f
C4780 AVSS.n5972 VSUBS 0.049193f
C4781 AVSS.t8 VSUBS 0.017259f
C4782 AVSS.t125 VSUBS 0.017259f
C4783 AVSS.n5973 VSUBS 0.590831f
C4784 AVSS.n5974 VSUBS 0.049193f
C4785 AVSS.n5975 VSUBS 0.59066f
C4786 AVSS.n5976 VSUBS 0.730673f
C4787 AVSS.t122 VSUBS 0.01648f
C4788 AVSS.n5977 VSUBS 0.399766f
C4789 AVSS.t35 VSUBS 4.25031f
C4790 AVSS.t23 VSUBS 2.14453f
C4791 AVSS.t34 VSUBS 2.14453f
C4792 AVSS.t38 VSUBS 2.14453f
C4793 AVSS.t42 VSUBS 1.66008f
C4794 AVSS.n5978 VSUBS 1.07227f
C4795 AVSS.t11 VSUBS 1.55672f
C4796 AVSS.t40 VSUBS 2.14453f
C4797 AVSS.t50 VSUBS 2.14453f
C4798 AVSS.t126 VSUBS 2.14453f
C4799 AVSS.t7 VSUBS 3.66896f
C4800 AVSS.t44 VSUBS 3.66896f
C4801 AVSS.t14 VSUBS 2.14453f
C4802 AVSS.t12 VSUBS 2.14453f
C4803 AVSS.t36 VSUBS 1.6084f
C4804 AVSS.t39 VSUBS 2.14453f
C4805 AVSS.t32 VSUBS 2.14453f
C4806 AVSS.t33 VSUBS 1.6084f
C4807 AVSS.n5979 VSUBS 1.07227f
C4808 AVSS.n5980 VSUBS 0.58644f
C4809 AVSS.n5981 VSUBS 0.58644f
C4810 AVSS.n5982 VSUBS 0.078665f
C4811 AVSS.t45 VSUBS 0.016573f
C4812 AVSS.n5983 VSUBS 0.488222f
C4813 AVSS.n5984 VSUBS 0.701796f
C4814 AVSS.n5985 VSUBS 0.689418f
C4815 AVSS.n5986 VSUBS 0.710826f
C4816 AVSS.n5987 VSUBS 0.70359f
C4817 AVSS.n5988 VSUBS 0.705111f
C4818 AVSS.n5989 VSUBS 0.703641f
C4819 AVSS.n5990 VSUBS 0.703641f
C4820 AVSS.n5991 VSUBS 9.86905f
C4821 AVSS.t10 VSUBS 29.627098f
C4822 AVSS.n5992 VSUBS 2.59669f
C4823 AVSS.n5993 VSUBS 0.434297f
C4824 AVSS.n5994 VSUBS 0.434297f
C4825 AVSS.n5995 VSUBS 0.435726f
C4826 AVSS.n5996 VSUBS 0.434297f
C4827 AVSS.n5997 VSUBS 0.434297f
C4828 AVSS.n5998 VSUBS 1.03351f
C4829 AVSS.n5999 VSUBS 2.5321f
C4830 AVSS.t5 VSUBS 4.66346f
C4831 AVSS.t47 VSUBS 4.456759f
C4832 AVSS.t120 VSUBS 0.015085f
C4833 AVSS.t119 VSUBS 0.015085f
C4834 AVSS.t118 VSUBS 0.015085f
C4835 AVSS.n6000 VSUBS 0.031937f
C4836 AVSS.t121 VSUBS 0.015085f
C4837 AVSS.n6001 VSUBS 0.102564f
C4838 AVSS.t115 VSUBS 0.015085f
C4839 AVSS.n6002 VSUBS 0.102564f
C4840 AVSS.t116 VSUBS 0.015085f
C4841 AVSS.n6003 VSUBS 0.031937f
C4842 AVSS.n6004 VSUBS 0.185706f
C4843 AVSS.n6005 VSUBS 0.103496f
C4844 AVSS.n6006 VSUBS 0.228677f
C4845 AVSS.n6007 VSUBS 0.169245f
C4846 AVSS.n6008 VSUBS 0.170485f
C4847 AVSS.n6009 VSUBS 0.114398f
C4848 AVSS.n6010 VSUBS 0.131014f
C4849 AVSS.n6011 VSUBS 0.170485f
C4850 AVSS.n6012 VSUBS 0.170485f
C4851 AVSS.n6013 VSUBS 2.17037f
C4852 AVSS.n6014 VSUBS 1.16916f
C4853 AVSS.n6015 VSUBS 0.169245f
C4854 AVSS.n6016 VSUBS 0.955997f
C4855 AVSS.t30 VSUBS 1.47921f
C4856 AVSS.t130 VSUBS 1.56318f
C4857 AVSS.t28 VSUBS 1.07227f
C4858 AVSS.t24 VSUBS 1.11748f
C4859 AVSS.n6017 VSUBS 0.124865f
C4860 AVSS.n6018 VSUBS 0.542593f
C4861 AVSS.n6019 VSUBS 0.536133f
C4862 AVSS.t127 VSUBS 1.60194f
C4863 AVSS.t22 VSUBS 1.13686f
C4864 AVSS.t27 VSUBS 1.07227f
C4865 AVSS.t48 VSUBS 1.42754f
C4866 AVSS.n6020 VSUBS 0.975375f
C4867 AVSS.n6021 VSUBS 0.955997f
C4868 AVSS.n6022 VSUBS 0.169245f
C4869 AVSS.n6023 VSUBS 0.169245f
C4870 AVSS.n6024 VSUBS 0.170485f
C4871 AVSS.n6025 VSUBS 0.192798f
C4872 AVSS.n6026 VSUBS 0.016216f
C4873 AVSS.n6027 VSUBS 0.254275f
C4874 AVSS.n6028 VSUBS 0.299832f
C4875 AVSS.n6029 VSUBS 0.310153f
C4876 AVSS.n6030 VSUBS 0.13307f
C4877 AVSS.n6031 VSUBS 0.132794f
C4878 AVSS.n6032 VSUBS 0.265586f
C4879 AVSS.n6033 VSUBS 2.54502f
C4880 AVSS.t15 VSUBS 5.12531f
C4881 AVSS.n6034 VSUBS 0.539647f
C4882 AVSS.n6035 VSUBS 0.265586f
C4883 AVSS.n6036 VSUBS 0.132794f
C4884 AVSS.n6037 VSUBS 0.13307f
C4885 AVSS.n6038 VSUBS 0.20733f
C4886 AVSS.n6039 VSUBS 0.065445f
C4887 AVSS.t52 VSUBS 0.016523f
C4888 AVSS.n6040 VSUBS 0.021923f
C4889 AVSS.t124 VSUBS 0.017242f
C4890 AVSS.n6041 VSUBS 0.194623f
C4891 AVSS.n6042 VSUBS 0.073629f
C4892 AVSS.n6043 VSUBS 0.125643f
C4893 AVSS.n6044 VSUBS 0.206531f
C4894 AVSS.t31 VSUBS 0.017226f
C4895 AVSS.n6045 VSUBS 0.165232f
C4896 AVSS.n6046 VSUBS 0.026572f
C4897 AVSS.t49 VSUBS 0.016872f
C4898 AVSS.n6047 VSUBS 0.086888f
C4899 AVSS.t21 VSUBS 0.017242f
C4900 AVSS.t26 VSUBS 0.016603f
C4901 AVSS.n6048 VSUBS 0.127674f
C4902 AVSS.n6049 VSUBS 0.194623f
C4903 AVSS.n6050 VSUBS 0.136902f
C4904 AVSS.n6051 VSUBS 0.123915f
C4905 AVSS.n6052 VSUBS 0.124865f
C4906 AVSS.n6053 VSUBS 0.124865f
C4907 AVSS.n6054 VSUBS 0.394631f
C4908 AVSS.t25 VSUBS 0.591947f
C4909 AVSS.t128 VSUBS 0.789263f
C4910 AVSS.t20 VSUBS 0.846318f
C4911 AVSS.n6055 VSUBS 0.529209f
C4912 AVSS.n6056 VSUBS 0.329246p
C4913 AVSS.n6057 VSUBS 56.4425f
C4914 AVSS.t17 VSUBS 15.429799f
C4915 AVSS.n6058 VSUBS 16.3579f
C4916 AVSS.n6059 VSUBS 0.58644f
C4917 AVSS.n6060 VSUBS 0.58644f
C4918 AVSS.n6061 VSUBS 0.055769f
C4919 AVSS.n6062 VSUBS 0.16088f
C4920 AVSS.n6063 VSUBS 1.04923f
C4921 AVSS.t55 VSUBS 17.1225f
C4922 AVSS.n6064 VSUBS 18.458f
C4923 AVSS.t71 VSUBS 17.1225f
C4924 AVSS.n6065 VSUBS 16.724901f
C4925 AVSS.t53 VSUBS 17.1225f
C4926 AVSS.n6066 VSUBS 14.814199f
C4927 AVSS.n6067 VSUBS 16.1531f
C4928 AVSS.t70 VSUBS 18.0884f
C4929 AVSS.n6068 VSUBS 5.81745f
C4930 AVSS.t73 VSUBS 17.1225f
C4931 AVSS.n6069 VSUBS 12.5678f
C4932 AVSS.t74 VSUBS 18.0884f
C4933 AVSS.n6070 VSUBS 5.38967f
C4934 AVSS.t61 VSUBS 17.1225f
C4935 AVSS.n6071 VSUBS 12.5678f
C4936 AVSS.t62 VSUBS 18.0884f
C4937 AVSS.n6072 VSUBS 5.38967f
C4938 AVSS.t63 VSUBS 17.1225f
C4939 AVSS.n6073 VSUBS 10.4677f
C4940 AVSS.n6074 VSUBS 5.28628f
C4941 AVSS.n6075 VSUBS 2.90165f
C4942 AVSS.n6076 VSUBS 1.79376f
C4943 AVSS.n6077 VSUBS 0.04959f
C4944 AVSS.n6079 VSUBS 0.07714f
C4945 AVSS.n6080 VSUBS 0.160158f
C4946 AVSS.n6081 VSUBS 0.043735f
C4947 AVSS.n6082 VSUBS 0.078223f
C4948 AVSS.n6083 VSUBS 0.110993f
C4949 AVSS.n6084 VSUBS 0.033852f
C4950 AVSS.n6085 VSUBS 0.018072f
C4951 AVSS.n6087 VSUBS 0.011633f
C4952 AVSS.n6088 VSUBS 0.014835f
C4953 AVSS.n6090 VSUBS 0.013464f
C4954 AVSS.n6092 VSUBS 0.013464f
C4955 AVSS.n6093 VSUBS 0.013197f
C4956 AVSS.n6094 VSUBS 0.013197f
C4957 AVSS.n6095 VSUBS 0.013197f
C4958 AVSS.n6096 VSUBS 0.013464f
C4959 AVSS.n6098 VSUBS 0.013464f
C4960 AVSS.n6100 VSUBS 0.013464f
C4961 AVSS.n6102 VSUBS 0.012464f
C4962 AVSS.n6103 VSUBS 0.013197f
C4963 AVSS.n6104 VSUBS 0.013464f
C4964 AVSS.n6106 VSUBS 0.013464f
C4965 AVSS.n6108 VSUBS 0.013464f
C4966 AVSS.n6109 VSUBS 0.013197f
C4967 AVSS.n6110 VSUBS 0.014549f
C4968 AVSS.n6111 VSUBS 0.016685f
C4969 AVSS.n6112 VSUBS 0.016888f
C4970 AVSS.n6113 VSUBS 0.013464f
C4971 AVSS.n6114 VSUBS 0.253149f
C4972 AVSS.n6115 VSUBS 0.253149f
C4973 AVSS.n6116 VSUBS 0.013464f
C4974 AVSS.n6117 VSUBS 0.013197f
C4975 AVSS.n6118 VSUBS 0.013197f
C4976 AVSS.n6119 VSUBS 0.013197f
C4977 AVSS.n6120 VSUBS 0.013464f
C4978 AVSS.n6121 VSUBS 0.253149f
C4979 AVSS.n6122 VSUBS 0.253149f
C4980 AVSS.n6123 VSUBS 0.167359f
C4981 AVSS.n6124 VSUBS 0.013464f
C4982 AVSS.n6125 VSUBS 0.013197f
C4983 AVSS.n6126 VSUBS 0.013197f
C4984 AVSS.n6127 VSUBS 0.013197f
C4985 AVSS.n6128 VSUBS 0.013464f
C4986 AVSS.n6129 VSUBS 0.253149f
C4987 AVSS.n6130 VSUBS 0.253149f
C4988 AVSS.n6131 VSUBS 0.253149f
C4989 AVSS.n6132 VSUBS 0.013464f
C4990 AVSS.n6133 VSUBS 0.013197f
C4991 AVSS.n6134 VSUBS 0.013197f
C4992 AVSS.n6135 VSUBS 0.018889f
C4993 AVSS.n6136 VSUBS 0.019048f
C4994 AVSS.n6137 VSUBS 0.383942f
C4995 AVSS.t84 VSUBS 2.95053f
C4996 AVSS.n6138 VSUBS 0.383942f
C4997 AVSS.n6139 VSUBS 0.019048f
C4998 AVSS.n6140 VSUBS 0.018889f
C4999 AVSS.n6141 VSUBS 0.013197f
C5000 AVSS.n6142 VSUBS 0.013197f
C5001 AVSS.n6143 VSUBS 0.013464f
C5002 AVSS.n6144 VSUBS 0.253149f
C5003 AVSS.n6145 VSUBS 0.253149f
C5004 AVSS.n6146 VSUBS 0.253149f
C5005 AVSS.n6147 VSUBS 0.013464f
C5006 AVSS.n6148 VSUBS 0.013197f
C5007 AVSS.n6149 VSUBS 0.013197f
C5008 AVSS.n6150 VSUBS 0.013197f
C5009 AVSS.n6151 VSUBS 0.013464f
C5010 AVSS.n6152 VSUBS 0.013464f
C5011 AVSS.n6153 VSUBS 0.253149f
C5012 AVSS.n6154 VSUBS 0.253149f
C5013 AVSS.n6155 VSUBS 0.013464f
C5014 AVSS.n6156 VSUBS 0.013197f
C5015 AVSS.n6157 VSUBS 0.013197f
C5016 AVSS.n6158 VSUBS 0.013197f
C5017 AVSS.n6159 VSUBS 0.013464f
C5018 AVSS.n6160 VSUBS 0.253149f
C5019 AVSS.n6161 VSUBS 0.654125f
C5020 AVSS.n6162 VSUBS 0.150221f
C5021 AVSS.n6163 VSUBS 0.016888f
C5022 AVSS.n6164 VSUBS 0.016685f
C5023 AVSS.n6165 VSUBS 0.014549f
C5024 AVSS.n6166 VSUBS 0.013197f
C5025 AVSS.n6167 VSUBS 0.013464f
C5026 AVSS.n6168 VSUBS 0.027461f
C5027 AVSS.n6169 VSUBS 0.027461f
C5028 AVSS.n6170 VSUBS 0.027461f
C5029 AVSS.n6171 VSUBS 0.013464f
C5030 AVSS.n6172 VSUBS 0.013197f
C5031 AVSS.n6173 VSUBS 0.012464f
C5032 AVSS.n6175 VSUBS 0.013464f
C5033 AVSS.n6176 VSUBS 0.020901f
C5034 AVSS.t85 VSUBS 0.200034f
C5035 AVSS.n6177 VSUBS 0.020291f
C5036 AVSS.n6178 VSUBS 0.027461f
C5037 AVSS.n6179 VSUBS 0.013464f
C5038 AVSS.n6180 VSUBS 0.013197f
C5039 AVSS.n6181 VSUBS 0.013197f
C5040 AVSS.n6182 VSUBS 0.013197f
C5041 AVSS.n6183 VSUBS 0.013464f
C5042 AVSS.n6184 VSUBS 0.027461f
C5043 AVSS.n6185 VSUBS 0.027461f
C5044 AVSS.n6186 VSUBS 0.029139f
C5045 AVSS.n6187 VSUBS 0.014835f
C5046 AVSS.n6188 VSUBS 0.014713f
C5047 AVSS.n6189 VSUBS 0.017108f
C5048 AVSS.n6190 VSUBS 0.013197f
C5049 AVSS.n6191 VSUBS 0.013464f
C5050 AVSS.n6193 VSUBS 0.013464f
C5051 AVSS.n6194 VSUBS 0.013464f
C5052 AVSS.n6195 VSUBS 0.013197f
C5053 AVSS.n6196 VSUBS 0.013197f
C5054 AVSS.n6197 VSUBS 0.013197f
C5055 AVSS.n6198 VSUBS 0.013464f
C5056 AVSS.n6200 VSUBS 0.013464f
C5057 AVSS.n6201 VSUBS 0.013464f
C5058 AVSS.n6202 VSUBS 0.013197f
C5059 AVSS.n6203 VSUBS 0.013197f
C5060 AVSS.n6204 VSUBS 0.013197f
C5061 AVSS.n6205 VSUBS 0.013464f
C5062 AVSS.n6207 VSUBS 0.013464f
C5063 AVSS.n6208 VSUBS 0.013464f
C5064 AVSS.n6211 VSUBS 0.012774f
C5065 AVSS.n6212 VSUBS 0.035594f
C5066 AVSS.n6213 VSUBS 0.157726f
C5067 AVSS.n6214 VSUBS 0.073801f
C5068 AVSS.n6215 VSUBS 0.078697f
C5069 AVSS.n6216 VSUBS 0.0733f
C5070 AVSS.n6217 VSUBS 0.149766f
C5071 AVSS.n6218 VSUBS 0.073801f
C5072 AVSS.n6219 VSUBS 0.078697f
C5073 AVSS.n6220 VSUBS 0.0733f
C5074 AVSS.n6221 VSUBS 0.149766f
C5075 AVSS.n6222 VSUBS 0.073801f
C5076 AVSS.n6223 VSUBS 0.078697f
C5077 AVSS.n6224 VSUBS 0.0733f
C5078 AVSS.n6225 VSUBS 0.129464f
C5079 AVSS.n6226 VSUBS 0.101099f
C5080 AVSS.n6227 VSUBS 0.04266f
C5081 AVSS.n6228 VSUBS 0.091973f
C5082 AVSS.n6229 VSUBS 0.166238f
C5083 AVSS.n6230 VSUBS 0.093787f
C5084 AVSS.n6231 VSUBS 0.067428f
C5085 AVSS.n6232 VSUBS 0.043157f
C5086 AVSS.n6233 VSUBS 0.033359f
C5087 AVSS.n6234 VSUBS 0.030324f
C5088 AVSS.n6235 VSUBS 0.051397f
C5089 AVSS.n6236 VSUBS 0.045828f
C5090 AVSS.t106 VSUBS 0.154434f
C5091 AVSS.n6237 VSUBS 0.205976f
C5092 AVSS.n6238 VSUBS 0.051397f
C5093 AVSS.n6239 VSUBS 0.077272f
C5094 AVSS.n6240 VSUBS 0.091803f
C5095 AVSS.n6241 VSUBS 0.160736f
C5096 AVSS.n6242 VSUBS 0.084368f
C5097 AVSS.n6243 VSUBS 0.11551f
C5098 AVSS.n6244 VSUBS 0.192018f
C5099 AVSS.n6245 VSUBS 0.210564f
C5100 AVSS.n6246 VSUBS 0.205814f
C5101 AVSS.n6247 VSUBS 0.04266f
C5102 AVSS.n6248 VSUBS 0.030324f
C5103 AVSS.n6249 VSUBS 0.090352f
C5104 AVSS.n6250 VSUBS 0.090352f
C5105 AVSS.n6251 VSUBS 0.046257f
C5106 AVSS.n6252 VSUBS 0.051397f
C5107 AVSS.n6253 VSUBS 0.077272f
C5108 AVSS.n6254 VSUBS 0.189601f
C5109 AVSS.n6255 VSUBS 0.186488f
C5110 AVSS.n6256 VSUBS 0.114153f
C5111 AVSS.n6257 VSUBS 0.192018f
C5112 AVSS.n6258 VSUBS 0.04266f
C5113 AVSS.n6259 VSUBS 0.210564f
C5114 AVSS.n6260 VSUBS 0.067428f
C5115 AVSS.n6261 VSUBS 0.090352f
C5116 AVSS.n6262 VSUBS 0.090352f
C5117 AVSS.n6263 VSUBS 0.030324f
C5118 AVSS.n6264 VSUBS 0.051397f
C5119 AVSS.n6265 VSUBS 0.045828f
C5120 AVSS.t89 VSUBS 0.154434f
C5121 AVSS.n6266 VSUBS 0.183064f
C5122 AVSS.n6267 VSUBS 0.013464f
C5123 AVSS.n6268 VSUBS 0.013197f
C5124 AVSS.n6269 VSUBS 0.013197f
C5125 AVSS.n6270 VSUBS 0.013197f
C5126 AVSS.n6271 VSUBS 0.013464f
C5127 AVSS.n6272 VSUBS 0.218223f
C5128 AVSS.n6273 VSUBS 0.218223f
C5129 AVSS.n6274 VSUBS 0.218223f
C5130 AVSS.n6275 VSUBS 0.013464f
C5131 AVSS.n6276 VSUBS 0.013197f
C5132 AVSS.n6277 VSUBS 0.01932f
C5133 AVSS.n6278 VSUBS 0.021004f
C5134 AVSS.n6279 VSUBS 0.021345f
C5135 AVSS.n6281 VSUBS 0.013464f
C5136 AVSS.n6283 VSUBS 0.013464f
C5137 AVSS.n6284 VSUBS 0.013197f
C5138 AVSS.n6285 VSUBS 0.013197f
C5139 AVSS.n6286 VSUBS 0.013197f
C5140 AVSS.n6287 VSUBS 0.013464f
C5141 AVSS.n6289 VSUBS 0.013464f
C5142 AVSS.n6291 VSUBS 0.013464f
C5143 AVSS.n6292 VSUBS 0.013197f
C5144 AVSS.n6293 VSUBS 0.013197f
C5145 AVSS.n6294 VSUBS 0.013197f
C5146 AVSS.n6295 VSUBS 0.013464f
C5147 AVSS.n6297 VSUBS 0.013464f
C5148 AVSS.n6298 VSUBS 0.013464f
C5149 AVSS.n6300 VSUBS 0.021194f
C5150 AVSS.n6301 VSUBS 0.018062f
C5151 AVSS.n6303 VSUBS 0.017854f
C5152 pmos_current_bgr_2_0.D3.n0 VSUBS 0.964488f
C5153 pmos_current_bgr_2_0.D3.n1 VSUBS 0.621049f
C5154 pmos_current_bgr_2_0.D3.t18 VSUBS 1.27469f
C5155 pmos_current_bgr_2_0.D3.t19 VSUBS 1.27469f
C5156 pmos_current_bgr_2_0.D3.t20 VSUBS 1.58062f
C5157 pmos_current_bgr_2_0.D3.t9 VSUBS 0.03203f
C5158 pmos_current_bgr_2_0.D3.t8 VSUBS 0.024637f
C5159 pmos_current_bgr_2_0.D3.n2 VSUBS 0.054715f
C5160 pmos_current_bgr_2_0.D3.t10 VSUBS 0.032456f
C5161 pmos_current_bgr_2_0.D3.t2 VSUBS 0.032456f
C5162 pmos_current_bgr_2_0.D3.t1 VSUBS 6.87815f
C5163 pmos_current_bgr_2_0.D3.n3 VSUBS 3.78633f
C5164 pmos_current_bgr_2_0.D3.t22 VSUBS 1.27469f
C5165 pmos_current_bgr_2_0.D3.n4 VSUBS 3.78633f
C5166 pmos_current_bgr_2_0.D3.n5 VSUBS 3.78633f
C5167 pmos_current_bgr_2_0.D3.t21 VSUBS 1.27469f
C5168 pmos_current_bgr_2_0.D3.t17 VSUBS 1.58062f
C5169 pmos_current_bgr_2_0.D3.n6 VSUBS 3.78633f
C5170 pmos_current_bgr_2_0.D3.t3 VSUBS 6.87787f
C5171 pmos_current_bgr_2_0.D3.t4 VSUBS 0.032456f
C5172 pmos_current_bgr_2_0.D3.t13 VSUBS 0.024637f
C5173 pmos_current_bgr_2_0.D3.t15 VSUBS 0.03203f
C5174 pmos_current_bgr_2_0.D3.n7 VSUBS 0.050407f
C5175 pmos_current_bgr_2_0.D3.t7 VSUBS 0.033815f
C5176 pmos_current_bgr_2_0.D3.t5 VSUBS 0.024912f
C5177 pmos_current_bgr_2_0.D3.n8 VSUBS 0.050953f
C5178 pmos_current_bgr_2_0.D3.n9 VSUBS 0.019008f
C5179 pmos_current_bgr_2_0.D3.n10 VSUBS 0.133232f
C5180 pmos_current_bgr_2_0.D3.t11 VSUBS 0.024912f
C5181 pmos_current_bgr_2_0.D3.n11 VSUBS 0.050953f
C5182 pmos_current_bgr_2_0.D3.t12 VSUBS 0.043057f
C5183 pmos_current_bgr_2_0.D3.n12 VSUBS 0.019008f
C5184 pmos_current_bgr_2_0.D3.n13 VSUBS 0.139741f
C5185 pmos_current_bgr_2_0.D3.n14 VSUBS 0.936257f
C5186 pmos_current_bgr_2_0.D3.t14 VSUBS 0.032456f
C5187 pmos_iptat_0.VDDE VSUBS 3.29859f
C5188 digital_0.VDDE.n0 VSUBS 2.01133f
C5189 digital_0.VDDE.n1 VSUBS 41.575302f
C5190 pmos_current_bgr_2_0.vdde VSUBS 3.88297f
C5191 digital_0.VDDE.n2 VSUBS 1.32996f
C5192 digital_0.VDDE.n3 VSUBS 0.537698f
C5193 pmos_current_bgr_2_0.VDDE VSUBS 1.89204f
C5194 pmos_current_bgr_0.vdde VSUBS 2.08863f
C5195 digital_0.VDDE.n4 VSUBS 3.08838f
C5196 pmos_startup_0.VDDE VSUBS 2.81298f
C5197 digital_0.VDDE.n5 VSUBS 4.45872f
C5198 digital_0.pmos_ena_0.VDDE VSUBS 2.36033f
C5199 digital_0.VDDE.n6 VSUBS 1.40819f
C5200 digital_0.VDDE.n7 VSUBS 2.51058f
C5201 digital_0.VDDE.t54 VSUBS 0.145776f
C5202 digital_0.VDDE.t72 VSUBS 0.145776f
C5203 digital_0.VDDE.n8 VSUBS 0.298078f
C5204 digital_0.VDDE.t53 VSUBS 0.533846f
C5205 digital_0.VDDE.n9 VSUBS 1.73189f
C5206 digital_0.VDDE.t49 VSUBS 0.145776f
C5207 digital_0.VDDE.t6 VSUBS 0.145776f
C5208 digital_0.VDDE.n10 VSUBS 0.298078f
C5209 digital_0.VDDE.t48 VSUBS 0.533846f
C5210 digital_0.VDDE.n11 VSUBS 2.21358f
C5211 digital_0.VDDE.n12 VSUBS 2.74045f
C5212 digital_0.VDDE.n13 VSUBS 2.77096f
C5213 digital_0.VDDE.n14 VSUBS 2.7836f
C5214 digital_0.VDDE.n15 VSUBS 2.7836f
C5215 digital_0.VDDE.n16 VSUBS 2.77096f
C5216 digital_0.VDDE.t73 VSUBS 0.072888f
C5217 digital_0.VDDE.t3 VSUBS 0.072888f
C5218 digital_0.VDDE.n17 VSUBS 0.149916f
C5219 digital_0.VDDE.t1 VSUBS 0.072888f
C5220 digital_0.VDDE.t24 VSUBS 0.072888f
C5221 digital_0.VDDE.n18 VSUBS 0.149916f
C5222 digital_0.VDDE.n19 VSUBS 0.63774f
C5223 digital_0.VDDE.t70 VSUBS 0.072888f
C5224 digital_0.VDDE.t9 VSUBS 0.072888f
C5225 digital_0.VDDE.n20 VSUBS 0.15509f
C5226 digital_0.VDDE.n21 VSUBS 2.0688f
C5227 digital_0.VDDE.t7 VSUBS 0.072888f
C5228 digital_0.VDDE.t10 VSUBS 0.072888f
C5229 digital_0.VDDE.n22 VSUBS 0.15509f
C5230 digital_0.VDDE.n23 VSUBS 2.06793f
C5231 digital_0.VDDE.n24 VSUBS 0.648454f
C5232 digital_0.VDDE.n25 VSUBS 2.40888f
C5233 digital_0.VDDE.n26 VSUBS 2.27903f
C5234 digital_0.VDDE.n27 VSUBS 2.284f
C5235 digital_0.VDDE.n28 VSUBS 2.27903f
C5236 digital_0.VDDE.n29 VSUBS 2.27903f
C5237 digital_0.VDDE.t0 VSUBS 0.936333f
C5238 digital_0.VDDE.n30 VSUBS 0.918738f
C5239 digital_0.VDDE.t15 VSUBS 0.072888f
C5240 digital_0.VDDE.t55 VSUBS 12.8564f
C5241 digital_0.VDDE.n31 VSUBS 2.10058f
C5242 digital_0.VDDE.t68 VSUBS 0.072888f
C5243 digital_0.VDDE.t17 VSUBS 0.072888f
C5244 digital_0.VDDE.n32 VSUBS 0.174445f
C5245 digital_0.VDDE.n33 VSUBS 2.38067f
C5246 digital_0.VDDE.n34 VSUBS 0.149916f
C5247 digital_0.VDDE.t56 VSUBS 0.145776f
C5248 digital_0.VDDE.t42 VSUBS 0.072888f
C5249 digital_0.VDDE.n35 VSUBS 0.149916f
C5250 digital_0.VDDE.t41 VSUBS 0.192014f
C5251 digital_0.VDDE.n36 VSUBS 0.214739f
C5252 digital_0.VDDE.t43 VSUBS 0.263613f
C5253 digital_0.VDDE.n37 VSUBS 0.186885f
C5254 digital_0.VDDE.n38 VSUBS 0.624756f
C5255 digital_0.VDDE.n39 VSUBS 1.66458f
C5256 digital_0.VDDE.n40 VSUBS 2.25861f
C5257 digital_0.VDDE.n41 VSUBS 2.25861f
C5258 digital_0.VDDE.n42 VSUBS 7.09551f
C5259 digital_0.VDDE.n43 VSUBS 4.56592f
C5260 digital_0.VDDE.n44 VSUBS 4.56506f
C5261 digital_0.VDDE.n45 VSUBS 2.28296f
C5262 digital_0.VDDE.n46 VSUBS 2.46694f
C5263 digital_0.VDDE.n47 VSUBS 4.58415f
C5264 digital_0.VDDE.n48 VSUBS 0.666343f
C5265 digital_0.VDDE.t67 VSUBS 0.072888f
C5266 digital_0.VDDE.t34 VSUBS 0.072888f
C5267 digital_0.VDDE.n49 VSUBS 0.15509f
C5268 digital_0.VDDE.n50 VSUBS 1.37111f
C5269 digital_0.VDDE.t66 VSUBS 0.072888f
C5270 digital_0.VDDE.t33 VSUBS 0.072888f
C5271 digital_0.VDDE.n51 VSUBS 0.15509f
C5272 digital_0.VDDE.n52 VSUBS 1.37111f
C5273 digital_0.VDDE.n53 VSUBS 0.666985f
C5274 digital_0.VDDE.t57 VSUBS 13.246201f
C5275 digital_0.VDDE.t44 VSUBS 13.246201f
C5276 digital_0.VDDE.n54 VSUBS 4.48308f
C5277 digital_0.VDDE.n55 VSUBS 0.390963f
C5278 digital_0.VDDE.t20 VSUBS 0.072888f
C5279 digital_0.VDDE.t69 VSUBS 0.072888f
C5280 digital_0.VDDE.n56 VSUBS 0.149916f
C5281 digital_0.VDDE.t46 VSUBS 0.145776f
C5282 digital_0.VDDE.n57 VSUBS 0.149916f
C5283 digital_0.VDDE.t58 VSUBS 0.145776f
C5284 digital_0.VDDE.n58 VSUBS 0.149916f
C5285 digital_0.VDDE.t71 VSUBS 0.072888f
C5286 digital_0.VDDE.t63 VSUBS 0.072888f
C5287 digital_0.VDDE.n59 VSUBS 0.149916f
C5288 digital_0.VDDE.t51 VSUBS 0.145776f
C5289 digital_0.VDDE.t39 VSUBS 13.246201f
C5290 digital_0.VDDE.t50 VSUBS 13.246201f
C5291 digital_0.VDDE.n60 VSUBS 4.48308f
C5292 digital_0.VDDE.n61 VSUBS 0.390385f
C5293 digital_0.VDDE.n62 VSUBS 0.149916f
C5294 digital_0.VDDE.t40 VSUBS 0.145776f
C5295 digital_0.VDDE.n63 VSUBS 0.149916f
C5296 digital_0.VDDE.n64 VSUBS 1.92349f
C5297 digital_0.VDDE.n65 VSUBS 2.13545f
C5298 digital_0.VDDE.t28 VSUBS 0.072888f
C5299 digital_0.VDDE.t30 VSUBS 0.072888f
C5300 digital_0.VDDE.n66 VSUBS 0.149916f
C5301 digital_0.VDDE.t27 VSUBS 0.072888f
C5302 digital_0.VDDE.t31 VSUBS 0.072888f
C5303 digital_0.VDDE.n67 VSUBS 0.149916f
C5304 digital_0.VDDE.n68 VSUBS 0.922444f
C5305 digital_0.VDDE.n69 VSUBS 0.883696f
C5306 digital_0.VDDE.n70 VSUBS 2.30552f
C5307 digital_0.VDDE.n71 VSUBS 2.30552f
C5308 digital_0.VDDE.n72 VSUBS 2.30552f
C5309 digital_0.VDDE.n73 VSUBS 2.05936f
C5310 digital_0.VDDE.n74 VSUBS 1.80964f
C5311 digital_0.VDDE.n75 VSUBS 2.3257f
C5312 digital_0.VDDE.n76 VSUBS 2.3257f
C5313 digital_0.VDDE.n77 VSUBS 2.30552f
C5314 digital_0.VDDE.t18 VSUBS 7.402339f
C5315 digital_0.VDDE.t4 VSUBS 41.1539f
C5316 digital_0.VDDE.t26 VSUBS 41.1539f
C5317 digital_0.VDDE.t19 VSUBS 39.4664f
C5318 digital_0.VDDE.n78 VSUBS 77.667f
C5319 digital_0.VDDE.t29 VSUBS 40.7321f
C5320 digital_0.VDDE.t21 VSUBS 40.7321f
C5321 digital_0.VDDE.n79 VSUBS 39.888298f
C5322 digital_0.VDDE.t8 VSUBS 6.5202f
C5323 digital_0.VDDE.n80 VSUBS 16.2609f
C5324 digital_0.VDDE.t35 VSUBS 50.959f
C5325 digital_0.VDDE.t32 VSUBS 0.120087p
C5326 digital_0.VDDE.t45 VSUBS 0.111879p
C5327 digital_0.VDDE.n81 VSUBS 39.0445f
C5328 digital_0.VDDE.n82 VSUBS 2.32484f
C5329 digital_0.VDDE.n83 VSUBS 2.32484f
C5330 digital_0.VDDE.n84 VSUBS 2.01838f
C5331 digital_0.VDDE.n85 VSUBS 2.07441f
C5332 digital_0.VDDE.n86 VSUBS 2.81367f
C5333 digital_0.VDDE.n87 VSUBS 0.65988f
C5334 digital_0.VDDE.t64 VSUBS 0.072888f
C5335 digital_0.VDDE.t22 VSUBS 0.072888f
C5336 digital_0.VDDE.n88 VSUBS 0.15509f
C5337 digital_0.VDDE.n89 VSUBS 1.37111f
C5338 digital_0.VDDE.t65 VSUBS 0.072888f
C5339 digital_0.VDDE.t23 VSUBS 0.072888f
C5340 digital_0.VDDE.n90 VSUBS 0.15509f
C5341 digital_0.VDDE.n91 VSUBS 1.37111f
C5342 digital_0.VDDE.n92 VSUBS 0.666985f
C5343 digital_0.VDDE.n93 VSUBS 3.21071f
C5344 digital_0.VDDE.n94 VSUBS 2.28467f
C5345 digital_0.VDDE.n95 VSUBS 3.213f
C5346 digital_0.VDDE.n96 VSUBS 3.82592f
C5347 digital_0.VDDE.n97 VSUBS 3.21191f
C5348 digital_0.VDDE.n98 VSUBS 2.28424f
C5349 digital_0.VDDE.n99 VSUBS 2.28253f
C5350 digital_0.VDDE.n100 VSUBS 4.58073f
C5351 digital_0.VDDE.n101 VSUBS 4.58073f
C5352 digital_0.VDDE.n102 VSUBS 11.122701f
C5353 digital_0.VDDE.n103 VSUBS 14.3061f
C5354 digital_0.VDDE.n104 VSUBS 8.36119f
C5355 digital_0.VDDE.t13 VSUBS 5.52299f
C5356 digital_0.VDDE.t12 VSUBS 41.1539f
C5357 digital_0.VDDE.t2 VSUBS 41.1539f
C5358 digital_0.VDDE.t16 VSUBS 39.4664f
C5359 digital_0.VDDE.t14 VSUBS 80.2571f
C5360 digital_0.VDDE.t25 VSUBS 39.8463f
C5361 digital_0.VDDE.t5 VSUBS 6.71071f
C5362 digital_0.VDDE.n105 VSUBS 8.91675f
C5363 digital_0.VDDE.n106 VSUBS 6.30806f
C5364 digital_0.VDDE.n107 VSUBS 2.77096f
C5365 digital_0.VDDE.n108 VSUBS 39.4664f
C5366 digital_0.VDDE.n109 VSUBS 39.4664f
C5367 digital_0.VDDE.n110 VSUBS 2.25861f
C5368 digital_0.VDDE.n111 VSUBS 2.25861f
C5369 digital_0.VDDE.n112 VSUBS 1.80865f
C5370 digital_0.VDDE.n113 VSUBS 2.17761f
C5371 digital_0.VDDE.n114 VSUBS 1.73089f
C5372 digital_0.VDDE.n115 VSUBS 2.77096f
C5373 digital_0.VDDE.n116 VSUBS 2.7836f
C5374 digital_0.VDDE.n117 VSUBS 2.41349f
C5375 digital_0.VDDE.n118 VSUBS 1.30154f
C5376 digital_0.VDDE.n119 VSUBS 46.069897f
C5377 digital_0.VDDE.t47 VSUBS 0.236377f
C5378 digital_0.VDDE.t52 VSUBS 0.236377f
C5379 digital_0.VDDE.n120 VSUBS 0.333673f
C5380 digital_0.VDDE.t61 VSUBS 0.539494f
C5381 digital_0.VDDE.t59 VSUBS 0.236377f
C5382 digital_0.VDDE.t36 VSUBS 0.236377f
C5383 digital_0.VDDE.n121 VSUBS 0.333673f
C5384 digital_0.VDDE.t38 VSUBS 0.539494f
C5385 digital_0.VDDE.n122 VSUBS 2.01117f
C5386 digital_0.VDDE.t62 VSUBS 0.145776f
C5387 digital_0.VDDE.t60 VSUBS 0.145776f
C5388 digital_0.VDDE.n123 VSUBS 0.304081f
C5389 digital_0.VDDE.t11 VSUBS 0.145776f
C5390 digital_0.VDDE.t37 VSUBS 0.145776f
C5391 digital_0.VDDE.n124 VSUBS 0.30386f
C5392 VREF.t13 VSUBS 0.01678f
C5393 VREF.n0 VSUBS 0.034697f
C5394 VREF.t14 VSUBS 0.01678f
C5395 VREF.n1 VSUBS 0.034781f
C5396 VREF.t7 VSUBS 0.078683f
C5397 VREF.t9 VSUBS 0.078683f
C5398 VREF.t8 VSUBS 0.031709f
C5399 VREF.t6 VSUBS 0.031709f
C5400 VREF.n2 VSUBS 0.068285f
C5401 VREF.n3 VSUBS 0.289158f
C5402 VREF.t1 VSUBS 0.01678f
C5403 VREF.t11 VSUBS 0.01678f
C5404 VREF.n4 VSUBS 0.034781f
C5405 VREF.t5 VSUBS 0.061653f
C5406 VREF.t2 VSUBS 0.01678f
C5407 VREF.t4 VSUBS 0.01678f
C5408 VREF.n5 VSUBS 0.034513f
C5409 VREF.t0 VSUBS 0.059536f
C5410 VREF.n6 VSUBS 1.72415f
C5411 VREF.n7 VSUBS 0.970837f
C5412 VREF.t12 VSUBS 0.061903f
C5413 VREF.t3 VSUBS 0.031709f
C5414 VREF.t10 VSUBS 0.031709f
C5415 VREF.n8 VSUBS 0.068285f
C5416 VREF.n9 VSUBS 0.176879f
C5417 VREF.n10 VSUBS 0.026169f
C5418 VREF.n11 VSUBS 1.63153f
C5419 VREF.n12 VSUBS 1.62262f
.ends

