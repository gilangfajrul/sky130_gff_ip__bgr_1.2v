magic
tech sky130A
magscale 1 2
timestamp 1762873293
<< pwell >>
rect -782 -7962 782 7962
<< psubdiff >>
rect -746 7892 -650 7926
rect 650 7892 746 7926
rect -746 7830 -712 7892
rect 712 7830 746 7892
rect -746 -7892 -712 -7830
rect 712 -7892 746 -7830
rect -746 -7926 -650 -7892
rect 650 -7926 746 -7892
<< psubdiffcont >>
rect -650 7892 650 7926
rect -746 -7830 -712 7830
rect 712 -7830 746 7830
rect -650 -7926 650 -7892
<< xpolycontact >>
rect -616 7364 -546 7796
rect -616 5284 -546 5716
rect -450 7364 -380 7796
rect -450 5284 -380 5716
rect -284 7364 -214 7796
rect -284 5284 -214 5716
rect -118 7364 -48 7796
rect -118 5284 -48 5716
rect 48 7364 118 7796
rect 48 5284 118 5716
rect 214 7364 284 7796
rect 214 5284 284 5716
rect 380 7364 450 7796
rect 380 5284 450 5716
rect 546 7364 616 7796
rect 546 5284 616 5716
rect -616 4748 -546 5180
rect -616 2668 -546 3100
rect -450 4748 -380 5180
rect -450 2668 -380 3100
rect -284 4748 -214 5180
rect -284 2668 -214 3100
rect -118 4748 -48 5180
rect -118 2668 -48 3100
rect 48 4748 118 5180
rect 48 2668 118 3100
rect 214 4748 284 5180
rect 214 2668 284 3100
rect 380 4748 450 5180
rect 380 2668 450 3100
rect 546 4748 616 5180
rect 546 2668 616 3100
rect -616 2132 -546 2564
rect -616 52 -546 484
rect -450 2132 -380 2564
rect -450 52 -380 484
rect -284 2132 -214 2564
rect -284 52 -214 484
rect -118 2132 -48 2564
rect -118 52 -48 484
rect 48 2132 118 2564
rect 48 52 118 484
rect 214 2132 284 2564
rect 214 52 284 484
rect 380 2132 450 2564
rect 380 52 450 484
rect 546 2132 616 2564
rect 546 52 616 484
rect -616 -484 -546 -52
rect -616 -2564 -546 -2132
rect -450 -484 -380 -52
rect -450 -2564 -380 -2132
rect -284 -484 -214 -52
rect -284 -2564 -214 -2132
rect -118 -484 -48 -52
rect -118 -2564 -48 -2132
rect 48 -484 118 -52
rect 48 -2564 118 -2132
rect 214 -484 284 -52
rect 214 -2564 284 -2132
rect 380 -484 450 -52
rect 380 -2564 450 -2132
rect 546 -484 616 -52
rect 546 -2564 616 -2132
rect -616 -3100 -546 -2668
rect -616 -5180 -546 -4748
rect -450 -3100 -380 -2668
rect -450 -5180 -380 -4748
rect -284 -3100 -214 -2668
rect -284 -5180 -214 -4748
rect -118 -3100 -48 -2668
rect -118 -5180 -48 -4748
rect 48 -3100 118 -2668
rect 48 -5180 118 -4748
rect 214 -3100 284 -2668
rect 214 -5180 284 -4748
rect 380 -3100 450 -2668
rect 380 -5180 450 -4748
rect 546 -3100 616 -2668
rect 546 -5180 616 -4748
rect -616 -5716 -546 -5284
rect -616 -7796 -546 -7364
rect -450 -5716 -380 -5284
rect -450 -7796 -380 -7364
rect -284 -5716 -214 -5284
rect -284 -7796 -214 -7364
rect -118 -5716 -48 -5284
rect -118 -7796 -48 -7364
rect 48 -5716 118 -5284
rect 48 -7796 118 -7364
rect 214 -5716 284 -5284
rect 214 -7796 284 -7364
rect 380 -5716 450 -5284
rect 380 -7796 450 -7364
rect 546 -5716 616 -5284
rect 546 -7796 616 -7364
<< ppolyres >>
rect -616 5716 -546 7364
rect -450 5716 -380 7364
rect -284 5716 -214 7364
rect -118 5716 -48 7364
rect 48 5716 118 7364
rect 214 5716 284 7364
rect 380 5716 450 7364
rect 546 5716 616 7364
rect -616 3100 -546 4748
rect -450 3100 -380 4748
rect -284 3100 -214 4748
rect -118 3100 -48 4748
rect 48 3100 118 4748
rect 214 3100 284 4748
rect 380 3100 450 4748
rect 546 3100 616 4748
rect -616 484 -546 2132
rect -450 484 -380 2132
rect -284 484 -214 2132
rect -118 484 -48 2132
rect 48 484 118 2132
rect 214 484 284 2132
rect 380 484 450 2132
rect 546 484 616 2132
rect -616 -2132 -546 -484
rect -450 -2132 -380 -484
rect -284 -2132 -214 -484
rect -118 -2132 -48 -484
rect 48 -2132 118 -484
rect 214 -2132 284 -484
rect 380 -2132 450 -484
rect 546 -2132 616 -484
rect -616 -4748 -546 -3100
rect -450 -4748 -380 -3100
rect -284 -4748 -214 -3100
rect -118 -4748 -48 -3100
rect 48 -4748 118 -3100
rect 214 -4748 284 -3100
rect 380 -4748 450 -3100
rect 546 -4748 616 -3100
rect -616 -7364 -546 -5716
rect -450 -7364 -380 -5716
rect -284 -7364 -214 -5716
rect -118 -7364 -48 -5716
rect 48 -7364 118 -5716
rect 214 -7364 284 -5716
rect 380 -7364 450 -5716
rect 546 -7364 616 -5716
<< locali >>
rect -666 7892 -650 7926
rect 650 7892 666 7926
rect -746 7830 -712 7846
rect 712 7830 746 7846
rect -746 -7846 -712 -7830
rect 712 -7846 746 -7830
rect -666 -7926 -650 -7892
rect 650 -7926 666 -7892
<< viali >>
rect -600 7381 -562 7778
rect -434 7381 -396 7778
rect -268 7381 -230 7778
rect -102 7381 -64 7778
rect 64 7381 102 7778
rect 230 7381 268 7778
rect 396 7381 434 7778
rect 562 7381 600 7778
rect -600 5302 -562 5699
rect -434 5302 -396 5699
rect -268 5302 -230 5699
rect -102 5302 -64 5699
rect 64 5302 102 5699
rect 230 5302 268 5699
rect 396 5302 434 5699
rect 562 5302 600 5699
rect -600 4765 -562 5162
rect -434 4765 -396 5162
rect -268 4765 -230 5162
rect -102 4765 -64 5162
rect 64 4765 102 5162
rect 230 4765 268 5162
rect 396 4765 434 5162
rect 562 4765 600 5162
rect -600 2686 -562 3083
rect -434 2686 -396 3083
rect -268 2686 -230 3083
rect -102 2686 -64 3083
rect 64 2686 102 3083
rect 230 2686 268 3083
rect 396 2686 434 3083
rect 562 2686 600 3083
rect -600 2149 -562 2546
rect -434 2149 -396 2546
rect -268 2149 -230 2546
rect -102 2149 -64 2546
rect 64 2149 102 2546
rect 230 2149 268 2546
rect 396 2149 434 2546
rect 562 2149 600 2546
rect -600 70 -562 467
rect -434 70 -396 467
rect -268 70 -230 467
rect -102 70 -64 467
rect 64 70 102 467
rect 230 70 268 467
rect 396 70 434 467
rect 562 70 600 467
rect -600 -467 -562 -70
rect -434 -467 -396 -70
rect -268 -467 -230 -70
rect -102 -467 -64 -70
rect 64 -467 102 -70
rect 230 -467 268 -70
rect 396 -467 434 -70
rect 562 -467 600 -70
rect -600 -2546 -562 -2149
rect -434 -2546 -396 -2149
rect -268 -2546 -230 -2149
rect -102 -2546 -64 -2149
rect 64 -2546 102 -2149
rect 230 -2546 268 -2149
rect 396 -2546 434 -2149
rect 562 -2546 600 -2149
rect -600 -3083 -562 -2686
rect -434 -3083 -396 -2686
rect -268 -3083 -230 -2686
rect -102 -3083 -64 -2686
rect 64 -3083 102 -2686
rect 230 -3083 268 -2686
rect 396 -3083 434 -2686
rect 562 -3083 600 -2686
rect -600 -5162 -562 -4765
rect -434 -5162 -396 -4765
rect -268 -5162 -230 -4765
rect -102 -5162 -64 -4765
rect 64 -5162 102 -4765
rect 230 -5162 268 -4765
rect 396 -5162 434 -4765
rect 562 -5162 600 -4765
rect -600 -5699 -562 -5302
rect -434 -5699 -396 -5302
rect -268 -5699 -230 -5302
rect -102 -5699 -64 -5302
rect 64 -5699 102 -5302
rect 230 -5699 268 -5302
rect 396 -5699 434 -5302
rect 562 -5699 600 -5302
rect -600 -7778 -562 -7381
rect -434 -7778 -396 -7381
rect -268 -7778 -230 -7381
rect -102 -7778 -64 -7381
rect 64 -7778 102 -7381
rect 230 -7778 268 -7381
rect 396 -7778 434 -7381
rect 562 -7778 600 -7381
<< metal1 >>
rect -606 7778 -556 7790
rect -606 7381 -600 7778
rect -562 7381 -556 7778
rect -606 7369 -556 7381
rect -440 7778 -390 7790
rect -440 7381 -434 7778
rect -396 7381 -390 7778
rect -440 7369 -390 7381
rect -274 7778 -224 7790
rect -274 7381 -268 7778
rect -230 7381 -224 7778
rect -274 7369 -224 7381
rect -108 7778 -58 7790
rect -108 7381 -102 7778
rect -64 7381 -58 7778
rect -108 7369 -58 7381
rect 58 7778 108 7790
rect 58 7381 64 7778
rect 102 7381 108 7778
rect 58 7369 108 7381
rect 224 7778 274 7790
rect 224 7381 230 7778
rect 268 7381 274 7778
rect 224 7369 274 7381
rect 390 7778 440 7790
rect 390 7381 396 7778
rect 434 7381 440 7778
rect 390 7369 440 7381
rect 556 7778 606 7790
rect 556 7381 562 7778
rect 600 7381 606 7778
rect 556 7369 606 7381
rect -606 5699 -556 5711
rect -606 5302 -600 5699
rect -562 5302 -556 5699
rect -606 5290 -556 5302
rect -440 5699 -390 5711
rect -440 5302 -434 5699
rect -396 5302 -390 5699
rect -440 5290 -390 5302
rect -274 5699 -224 5711
rect -274 5302 -268 5699
rect -230 5302 -224 5699
rect -274 5290 -224 5302
rect -108 5699 -58 5711
rect -108 5302 -102 5699
rect -64 5302 -58 5699
rect -108 5290 -58 5302
rect 58 5699 108 5711
rect 58 5302 64 5699
rect 102 5302 108 5699
rect 58 5290 108 5302
rect 224 5699 274 5711
rect 224 5302 230 5699
rect 268 5302 274 5699
rect 224 5290 274 5302
rect 390 5699 440 5711
rect 390 5302 396 5699
rect 434 5302 440 5699
rect 390 5290 440 5302
rect 556 5699 606 5711
rect 556 5302 562 5699
rect 600 5302 606 5699
rect 556 5290 606 5302
rect -606 5162 -556 5174
rect -606 4765 -600 5162
rect -562 4765 -556 5162
rect -606 4753 -556 4765
rect -440 5162 -390 5174
rect -440 4765 -434 5162
rect -396 4765 -390 5162
rect -440 4753 -390 4765
rect -274 5162 -224 5174
rect -274 4765 -268 5162
rect -230 4765 -224 5162
rect -274 4753 -224 4765
rect -108 5162 -58 5174
rect -108 4765 -102 5162
rect -64 4765 -58 5162
rect -108 4753 -58 4765
rect 58 5162 108 5174
rect 58 4765 64 5162
rect 102 4765 108 5162
rect 58 4753 108 4765
rect 224 5162 274 5174
rect 224 4765 230 5162
rect 268 4765 274 5162
rect 224 4753 274 4765
rect 390 5162 440 5174
rect 390 4765 396 5162
rect 434 4765 440 5162
rect 390 4753 440 4765
rect 556 5162 606 5174
rect 556 4765 562 5162
rect 600 4765 606 5162
rect 556 4753 606 4765
rect -606 3083 -556 3095
rect -606 2686 -600 3083
rect -562 2686 -556 3083
rect -606 2674 -556 2686
rect -440 3083 -390 3095
rect -440 2686 -434 3083
rect -396 2686 -390 3083
rect -440 2674 -390 2686
rect -274 3083 -224 3095
rect -274 2686 -268 3083
rect -230 2686 -224 3083
rect -274 2674 -224 2686
rect -108 3083 -58 3095
rect -108 2686 -102 3083
rect -64 2686 -58 3083
rect -108 2674 -58 2686
rect 58 3083 108 3095
rect 58 2686 64 3083
rect 102 2686 108 3083
rect 58 2674 108 2686
rect 224 3083 274 3095
rect 224 2686 230 3083
rect 268 2686 274 3083
rect 224 2674 274 2686
rect 390 3083 440 3095
rect 390 2686 396 3083
rect 434 2686 440 3083
rect 390 2674 440 2686
rect 556 3083 606 3095
rect 556 2686 562 3083
rect 600 2686 606 3083
rect 556 2674 606 2686
rect -606 2546 -556 2558
rect -606 2149 -600 2546
rect -562 2149 -556 2546
rect -606 2137 -556 2149
rect -440 2546 -390 2558
rect -440 2149 -434 2546
rect -396 2149 -390 2546
rect -440 2137 -390 2149
rect -274 2546 -224 2558
rect -274 2149 -268 2546
rect -230 2149 -224 2546
rect -274 2137 -224 2149
rect -108 2546 -58 2558
rect -108 2149 -102 2546
rect -64 2149 -58 2546
rect -108 2137 -58 2149
rect 58 2546 108 2558
rect 58 2149 64 2546
rect 102 2149 108 2546
rect 58 2137 108 2149
rect 224 2546 274 2558
rect 224 2149 230 2546
rect 268 2149 274 2546
rect 224 2137 274 2149
rect 390 2546 440 2558
rect 390 2149 396 2546
rect 434 2149 440 2546
rect 390 2137 440 2149
rect 556 2546 606 2558
rect 556 2149 562 2546
rect 600 2149 606 2546
rect 556 2137 606 2149
rect -606 467 -556 479
rect -606 70 -600 467
rect -562 70 -556 467
rect -606 58 -556 70
rect -440 467 -390 479
rect -440 70 -434 467
rect -396 70 -390 467
rect -440 58 -390 70
rect -274 467 -224 479
rect -274 70 -268 467
rect -230 70 -224 467
rect -274 58 -224 70
rect -108 467 -58 479
rect -108 70 -102 467
rect -64 70 -58 467
rect -108 58 -58 70
rect 58 467 108 479
rect 58 70 64 467
rect 102 70 108 467
rect 58 58 108 70
rect 224 467 274 479
rect 224 70 230 467
rect 268 70 274 467
rect 224 58 274 70
rect 390 467 440 479
rect 390 70 396 467
rect 434 70 440 467
rect 390 58 440 70
rect 556 467 606 479
rect 556 70 562 467
rect 600 70 606 467
rect 556 58 606 70
rect -606 -70 -556 -58
rect -606 -467 -600 -70
rect -562 -467 -556 -70
rect -606 -479 -556 -467
rect -440 -70 -390 -58
rect -440 -467 -434 -70
rect -396 -467 -390 -70
rect -440 -479 -390 -467
rect -274 -70 -224 -58
rect -274 -467 -268 -70
rect -230 -467 -224 -70
rect -274 -479 -224 -467
rect -108 -70 -58 -58
rect -108 -467 -102 -70
rect -64 -467 -58 -70
rect -108 -479 -58 -467
rect 58 -70 108 -58
rect 58 -467 64 -70
rect 102 -467 108 -70
rect 58 -479 108 -467
rect 224 -70 274 -58
rect 224 -467 230 -70
rect 268 -467 274 -70
rect 224 -479 274 -467
rect 390 -70 440 -58
rect 390 -467 396 -70
rect 434 -467 440 -70
rect 390 -479 440 -467
rect 556 -70 606 -58
rect 556 -467 562 -70
rect 600 -467 606 -70
rect 556 -479 606 -467
rect -606 -2149 -556 -2137
rect -606 -2546 -600 -2149
rect -562 -2546 -556 -2149
rect -606 -2558 -556 -2546
rect -440 -2149 -390 -2137
rect -440 -2546 -434 -2149
rect -396 -2546 -390 -2149
rect -440 -2558 -390 -2546
rect -274 -2149 -224 -2137
rect -274 -2546 -268 -2149
rect -230 -2546 -224 -2149
rect -274 -2558 -224 -2546
rect -108 -2149 -58 -2137
rect -108 -2546 -102 -2149
rect -64 -2546 -58 -2149
rect -108 -2558 -58 -2546
rect 58 -2149 108 -2137
rect 58 -2546 64 -2149
rect 102 -2546 108 -2149
rect 58 -2558 108 -2546
rect 224 -2149 274 -2137
rect 224 -2546 230 -2149
rect 268 -2546 274 -2149
rect 224 -2558 274 -2546
rect 390 -2149 440 -2137
rect 390 -2546 396 -2149
rect 434 -2546 440 -2149
rect 390 -2558 440 -2546
rect 556 -2149 606 -2137
rect 556 -2546 562 -2149
rect 600 -2546 606 -2149
rect 556 -2558 606 -2546
rect -606 -2686 -556 -2674
rect -606 -3083 -600 -2686
rect -562 -3083 -556 -2686
rect -606 -3095 -556 -3083
rect -440 -2686 -390 -2674
rect -440 -3083 -434 -2686
rect -396 -3083 -390 -2686
rect -440 -3095 -390 -3083
rect -274 -2686 -224 -2674
rect -274 -3083 -268 -2686
rect -230 -3083 -224 -2686
rect -274 -3095 -224 -3083
rect -108 -2686 -58 -2674
rect -108 -3083 -102 -2686
rect -64 -3083 -58 -2686
rect -108 -3095 -58 -3083
rect 58 -2686 108 -2674
rect 58 -3083 64 -2686
rect 102 -3083 108 -2686
rect 58 -3095 108 -3083
rect 224 -2686 274 -2674
rect 224 -3083 230 -2686
rect 268 -3083 274 -2686
rect 224 -3095 274 -3083
rect 390 -2686 440 -2674
rect 390 -3083 396 -2686
rect 434 -3083 440 -2686
rect 390 -3095 440 -3083
rect 556 -2686 606 -2674
rect 556 -3083 562 -2686
rect 600 -3083 606 -2686
rect 556 -3095 606 -3083
rect -606 -4765 -556 -4753
rect -606 -5162 -600 -4765
rect -562 -5162 -556 -4765
rect -606 -5174 -556 -5162
rect -440 -4765 -390 -4753
rect -440 -5162 -434 -4765
rect -396 -5162 -390 -4765
rect -440 -5174 -390 -5162
rect -274 -4765 -224 -4753
rect -274 -5162 -268 -4765
rect -230 -5162 -224 -4765
rect -274 -5174 -224 -5162
rect -108 -4765 -58 -4753
rect -108 -5162 -102 -4765
rect -64 -5162 -58 -4765
rect -108 -5174 -58 -5162
rect 58 -4765 108 -4753
rect 58 -5162 64 -4765
rect 102 -5162 108 -4765
rect 58 -5174 108 -5162
rect 224 -4765 274 -4753
rect 224 -5162 230 -4765
rect 268 -5162 274 -4765
rect 224 -5174 274 -5162
rect 390 -4765 440 -4753
rect 390 -5162 396 -4765
rect 434 -5162 440 -4765
rect 390 -5174 440 -5162
rect 556 -4765 606 -4753
rect 556 -5162 562 -4765
rect 600 -5162 606 -4765
rect 556 -5174 606 -5162
rect -606 -5302 -556 -5290
rect -606 -5699 -600 -5302
rect -562 -5699 -556 -5302
rect -606 -5711 -556 -5699
rect -440 -5302 -390 -5290
rect -440 -5699 -434 -5302
rect -396 -5699 -390 -5302
rect -440 -5711 -390 -5699
rect -274 -5302 -224 -5290
rect -274 -5699 -268 -5302
rect -230 -5699 -224 -5302
rect -274 -5711 -224 -5699
rect -108 -5302 -58 -5290
rect -108 -5699 -102 -5302
rect -64 -5699 -58 -5302
rect -108 -5711 -58 -5699
rect 58 -5302 108 -5290
rect 58 -5699 64 -5302
rect 102 -5699 108 -5302
rect 58 -5711 108 -5699
rect 224 -5302 274 -5290
rect 224 -5699 230 -5302
rect 268 -5699 274 -5302
rect 224 -5711 274 -5699
rect 390 -5302 440 -5290
rect 390 -5699 396 -5302
rect 434 -5699 440 -5302
rect 390 -5711 440 -5699
rect 556 -5302 606 -5290
rect 556 -5699 562 -5302
rect 600 -5699 606 -5302
rect 556 -5711 606 -5699
rect -606 -7381 -556 -7369
rect -606 -7778 -600 -7381
rect -562 -7778 -556 -7381
rect -606 -7790 -556 -7778
rect -440 -7381 -390 -7369
rect -440 -7778 -434 -7381
rect -396 -7778 -390 -7381
rect -440 -7790 -390 -7778
rect -274 -7381 -224 -7369
rect -274 -7778 -268 -7381
rect -230 -7778 -224 -7381
rect -274 -7790 -224 -7778
rect -108 -7381 -58 -7369
rect -108 -7778 -102 -7381
rect -64 -7778 -58 -7381
rect -108 -7790 -58 -7778
rect 58 -7381 108 -7369
rect 58 -7778 64 -7381
rect 102 -7778 108 -7381
rect 58 -7790 108 -7778
rect 224 -7381 274 -7369
rect 224 -7778 230 -7381
rect 268 -7778 274 -7381
rect 224 -7790 274 -7778
rect 390 -7381 440 -7369
rect 390 -7778 396 -7381
rect 434 -7778 440 -7381
rect 390 -7790 440 -7778
rect 556 -7381 606 -7369
rect 556 -7778 562 -7381
rect 600 -7778 606 -7381
rect 556 -7790 606 -7778
<< labels >>
rlabel psubdiffcont 0 -7909 0 -7909 0 B
port 1 nsew
rlabel xpolycontact -581 -5319 -581 -5319 0 R1_0_0
port 2 nsew
rlabel xpolycontact -581 -7761 -581 -7761 0 R2_0_0
port 3 nsew
rlabel xpolycontact -581 -2703 -581 -2703 0 R1_0_1
port 4 nsew
rlabel xpolycontact -581 -5145 -581 -5145 0 R2_0_1
port 5 nsew
rlabel xpolycontact -581 -87 -581 -87 0 R1_0_2
port 6 nsew
rlabel xpolycontact -581 -2529 -581 -2529 0 R2_0_2
port 7 nsew
rlabel xpolycontact -581 2529 -581 2529 0 R1_0_3
port 8 nsew
rlabel xpolycontact -581 87 -581 87 0 R2_0_3
port 9 nsew
rlabel xpolycontact -581 5145 -581 5145 0 R1_0_4
port 10 nsew
rlabel xpolycontact -581 2703 -581 2703 0 R2_0_4
port 11 nsew
rlabel xpolycontact -581 7761 -581 7761 0 R1_0_5
port 12 nsew
rlabel xpolycontact -581 5319 -581 5319 0 R2_0_5
port 13 nsew
rlabel xpolycontact -415 -5319 -415 -5319 0 R1_1_0
port 14 nsew
rlabel xpolycontact -415 -7761 -415 -7761 0 R2_1_0
port 15 nsew
rlabel xpolycontact -415 -2703 -415 -2703 0 R1_1_1
port 16 nsew
rlabel xpolycontact -415 -5145 -415 -5145 0 R2_1_1
port 17 nsew
rlabel xpolycontact -415 -87 -415 -87 0 R1_1_2
port 18 nsew
rlabel xpolycontact -415 -2529 -415 -2529 0 R2_1_2
port 19 nsew
rlabel xpolycontact -415 2529 -415 2529 0 R1_1_3
port 20 nsew
rlabel xpolycontact -415 87 -415 87 0 R2_1_3
port 21 nsew
rlabel xpolycontact -415 5145 -415 5145 0 R1_1_4
port 22 nsew
rlabel xpolycontact -415 2703 -415 2703 0 R2_1_4
port 23 nsew
rlabel xpolycontact -415 7761 -415 7761 0 R1_1_5
port 24 nsew
rlabel xpolycontact -415 5319 -415 5319 0 R2_1_5
port 25 nsew
rlabel xpolycontact -249 -5319 -249 -5319 0 R1_2_0
port 26 nsew
rlabel xpolycontact -249 -7761 -249 -7761 0 R2_2_0
port 27 nsew
rlabel xpolycontact -249 -2703 -249 -2703 0 R1_2_1
port 28 nsew
rlabel xpolycontact -249 -5145 -249 -5145 0 R2_2_1
port 29 nsew
rlabel xpolycontact -249 -87 -249 -87 0 R1_2_2
port 30 nsew
rlabel xpolycontact -249 -2529 -249 -2529 0 R2_2_2
port 31 nsew
rlabel xpolycontact -249 2529 -249 2529 0 R1_2_3
port 32 nsew
rlabel xpolycontact -249 87 -249 87 0 R2_2_3
port 33 nsew
rlabel xpolycontact -249 5145 -249 5145 0 R1_2_4
port 34 nsew
rlabel xpolycontact -249 2703 -249 2703 0 R2_2_4
port 35 nsew
rlabel xpolycontact -249 7761 -249 7761 0 R1_2_5
port 36 nsew
rlabel xpolycontact -249 5319 -249 5319 0 R2_2_5
port 37 nsew
rlabel xpolycontact -83 -5319 -83 -5319 0 R1_3_0
port 38 nsew
rlabel xpolycontact -83 -7761 -83 -7761 0 R2_3_0
port 39 nsew
rlabel xpolycontact -83 -2703 -83 -2703 0 R1_3_1
port 40 nsew
rlabel xpolycontact -83 -5145 -83 -5145 0 R2_3_1
port 41 nsew
rlabel xpolycontact -83 -87 -83 -87 0 R1_3_2
port 42 nsew
rlabel xpolycontact -83 -2529 -83 -2529 0 R2_3_2
port 43 nsew
rlabel xpolycontact -83 2529 -83 2529 0 R1_3_3
port 44 nsew
rlabel xpolycontact -83 87 -83 87 0 R2_3_3
port 45 nsew
rlabel xpolycontact -83 5145 -83 5145 0 R1_3_4
port 46 nsew
rlabel xpolycontact -83 2703 -83 2703 0 R2_3_4
port 47 nsew
rlabel xpolycontact -83 7761 -83 7761 0 R1_3_5
port 48 nsew
rlabel xpolycontact -83 5319 -83 5319 0 R2_3_5
port 49 nsew
rlabel xpolycontact 83 -5319 83 -5319 0 R1_4_0
port 50 nsew
rlabel xpolycontact 83 -7761 83 -7761 0 R2_4_0
port 51 nsew
rlabel xpolycontact 83 -2703 83 -2703 0 R1_4_1
port 52 nsew
rlabel xpolycontact 83 -5145 83 -5145 0 R2_4_1
port 53 nsew
rlabel xpolycontact 83 -87 83 -87 0 R1_4_2
port 54 nsew
rlabel xpolycontact 83 -2529 83 -2529 0 R2_4_2
port 55 nsew
rlabel xpolycontact 83 2529 83 2529 0 R1_4_3
port 56 nsew
rlabel xpolycontact 83 87 83 87 0 R2_4_3
port 57 nsew
rlabel xpolycontact 83 5145 83 5145 0 R1_4_4
port 58 nsew
rlabel xpolycontact 83 2703 83 2703 0 R2_4_4
port 59 nsew
rlabel xpolycontact 83 7761 83 7761 0 R1_4_5
port 60 nsew
rlabel xpolycontact 83 5319 83 5319 0 R2_4_5
port 61 nsew
rlabel xpolycontact 249 -5319 249 -5319 0 R1_5_0
port 62 nsew
rlabel xpolycontact 249 -7761 249 -7761 0 R2_5_0
port 63 nsew
rlabel xpolycontact 249 -2703 249 -2703 0 R1_5_1
port 64 nsew
rlabel xpolycontact 249 -5145 249 -5145 0 R2_5_1
port 65 nsew
rlabel xpolycontact 249 -87 249 -87 0 R1_5_2
port 66 nsew
rlabel xpolycontact 249 -2529 249 -2529 0 R2_5_2
port 67 nsew
rlabel xpolycontact 249 2529 249 2529 0 R1_5_3
port 68 nsew
rlabel xpolycontact 249 87 249 87 0 R2_5_3
port 69 nsew
rlabel xpolycontact 249 5145 249 5145 0 R1_5_4
port 70 nsew
rlabel xpolycontact 249 2703 249 2703 0 R2_5_4
port 71 nsew
rlabel xpolycontact 249 7761 249 7761 0 R1_5_5
port 72 nsew
rlabel xpolycontact 249 5319 249 5319 0 R2_5_5
port 73 nsew
rlabel xpolycontact 415 -5319 415 -5319 0 R1_6_0
port 74 nsew
rlabel xpolycontact 415 -7761 415 -7761 0 R2_6_0
port 75 nsew
rlabel xpolycontact 415 -2703 415 -2703 0 R1_6_1
port 76 nsew
rlabel xpolycontact 415 -5145 415 -5145 0 R2_6_1
port 77 nsew
rlabel xpolycontact 415 -87 415 -87 0 R1_6_2
port 78 nsew
rlabel xpolycontact 415 -2529 415 -2529 0 R2_6_2
port 79 nsew
rlabel xpolycontact 415 2529 415 2529 0 R1_6_3
port 80 nsew
rlabel xpolycontact 415 87 415 87 0 R2_6_3
port 81 nsew
rlabel xpolycontact 415 5145 415 5145 0 R1_6_4
port 82 nsew
rlabel xpolycontact 415 2703 415 2703 0 R2_6_4
port 83 nsew
rlabel xpolycontact 415 7761 415 7761 0 R1_6_5
port 84 nsew
rlabel xpolycontact 415 5319 415 5319 0 R2_6_5
port 85 nsew
rlabel xpolycontact 581 -5319 581 -5319 0 R1_7_0
port 86 nsew
rlabel xpolycontact 581 -7761 581 -7761 0 R2_7_0
port 87 nsew
rlabel xpolycontact 581 -2703 581 -2703 0 R1_7_1
port 88 nsew
rlabel xpolycontact 581 -5145 581 -5145 0 R2_7_1
port 89 nsew
rlabel xpolycontact 581 -87 581 -87 0 R1_7_2
port 90 nsew
rlabel xpolycontact 581 -2529 581 -2529 0 R2_7_2
port 91 nsew
rlabel xpolycontact 581 2529 581 2529 0 R1_7_3
port 92 nsew
rlabel xpolycontact 581 87 581 87 0 R2_7_3
port 93 nsew
rlabel xpolycontact 581 5145 581 5145 0 R1_7_4
port 94 nsew
rlabel xpolycontact 581 2703 581 2703 0 R2_7_4
port 95 nsew
rlabel xpolycontact 581 7761 581 7761 0 R1_7_5
port 96 nsew
rlabel xpolycontact 581 5319 581 5319 0 R2_7_5
port 97 nsew
<< properties >>
string FIXED_BBOX -729 -7909 729 7909
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.350 l 8.4 m 6 nx 8 wmin 0.350 lmin 0.50 class resistor rho 319.8 val 8.788k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 0 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0 doports 1
<< end >>
