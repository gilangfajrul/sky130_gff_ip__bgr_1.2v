magic
tech sky130A
magscale 1 2
timestamp 1717071607
<< nwell >>
rect -386 1770 8352 2798
rect -386 1764 8158 1770
rect 8160 1764 8352 1770
rect -386 934 8352 1764
<< nsubdiff >>
rect -350 2728 -290 2762
rect 8256 2728 8316 2762
rect -350 2702 -316 2728
rect 8282 2702 8316 2728
rect -350 1004 -316 1030
rect 8282 1004 8316 1030
rect -350 970 -290 1004
rect 8256 970 8316 1004
<< nsubdiffcont >>
rect -290 2728 8256 2762
rect -350 1030 -316 2702
rect 8282 1030 8316 2702
rect -290 970 8256 1004
<< poly >>
rect -228 2690 -162 2706
rect -228 2656 -212 2690
rect -178 2656 -162 2690
rect -228 2640 -162 2656
rect -192 2609 -162 2640
rect 8128 2690 8194 2706
rect 8128 2656 8144 2690
rect 8178 2656 8194 2690
rect 8128 2640 8194 2656
rect 8128 2609 8158 2640
rect -192 1962 -162 1993
rect -254 1946 -162 1962
rect -254 1912 -238 1946
rect -204 1912 -162 1946
rect -254 1896 -162 1912
rect 8128 1962 8158 1993
rect 8128 1946 8220 1962
rect 8128 1912 8170 1946
rect 8204 1912 8220 1946
rect 8128 1896 8220 1912
rect -254 1820 -162 1836
rect -254 1786 -238 1820
rect -204 1786 -162 1820
rect -254 1770 -162 1786
rect -192 1739 -162 1770
rect 8128 1820 8220 1836
rect 8128 1786 8170 1820
rect 8204 1786 8220 1820
rect 8128 1770 8220 1786
rect 8128 1764 8158 1770
rect -192 1092 -162 1123
rect -228 1076 -162 1092
rect -228 1042 -212 1076
rect -178 1042 -162 1076
rect -228 1026 -162 1042
rect 8128 1092 8158 1123
rect 8128 1076 8194 1092
rect 8128 1042 8144 1076
rect 8178 1042 8194 1076
rect 8128 1026 8194 1042
<< polycont >>
rect -212 2656 -178 2690
rect 8144 2656 8178 2690
rect -238 1912 -204 1946
rect 8170 1912 8204 1946
rect -238 1786 -204 1820
rect 8170 1786 8204 1820
rect -212 1042 -178 1076
rect 8144 1042 8178 1076
<< locali >>
rect -350 2728 -290 2762
rect 8256 2728 8316 2762
rect -350 2702 -316 2728
rect 8282 2702 8316 2728
rect -238 2656 -212 2690
rect -178 2656 -162 2690
rect 8128 2656 8144 2690
rect 8178 2656 8204 2690
rect -238 2609 -204 2656
rect 8170 2609 8204 2656
rect -238 1946 -204 1993
rect -238 1896 -204 1912
rect 8170 1946 8204 1993
rect 8170 1896 8204 1912
rect -238 1820 -204 1836
rect -238 1739 -204 1786
rect 8170 1820 8204 1836
rect 8170 1739 8204 1786
rect -238 1076 -204 1123
rect 8170 1076 8204 1123
rect -238 1042 -212 1076
rect -178 1042 -162 1076
rect 8128 1042 8144 1076
rect 8178 1042 8204 1076
rect -350 1004 -316 1030
rect 8282 1004 8316 1030
rect -350 970 -290 1004
rect 8256 970 8316 1004
<< viali >>
rect -212 2728 -178 2762
rect 1908 2728 1942 2762
rect 6024 2728 6058 2762
rect 8144 2728 8178 2762
rect -212 2656 -178 2690
rect 8144 2656 8178 2690
rect -350 1912 -316 1946
rect -238 1912 -204 1946
rect 8170 1912 8204 1946
rect 8282 1912 8316 1946
rect -350 1786 -316 1820
rect -238 1786 -204 1820
rect 8170 1786 8204 1820
rect 8282 1786 8316 1820
rect -212 1042 -178 1076
rect 8144 1042 8178 1076
rect -212 970 -178 1004
rect 1908 970 1942 1004
rect 6024 970 6058 1004
rect 8144 970 8178 1004
<< metal1 >>
rect -224 2762 -166 2768
rect -224 2728 -212 2762
rect -178 2728 -166 2762
rect -224 2696 -166 2728
rect -244 2690 -166 2696
rect -244 2656 -212 2690
rect -178 2656 -166 2690
rect -244 2650 -166 2656
rect 1896 2762 1954 2768
rect 1896 2728 1908 2762
rect 1942 2728 1954 2762
rect -244 2609 -198 2650
rect 1896 2597 1954 2728
rect 6012 2762 6070 2768
rect 6012 2728 6024 2762
rect 6058 2728 6070 2762
rect 6012 2597 6070 2728
rect 8132 2762 8190 2768
rect 8132 2728 8144 2762
rect 8178 2728 8190 2762
rect 8132 2696 8190 2728
rect 8132 2690 8210 2696
rect 8132 2656 8144 2690
rect 8178 2656 8210 2690
rect 8132 2650 8210 2656
rect 8164 2609 8210 2650
rect 1889 2421 1899 2597
rect 1951 2421 1961 2597
rect 3947 2421 3957 2597
rect 4009 2421 4019 2597
rect 6005 2421 6015 2597
rect 6067 2421 6077 2597
rect -156 2291 -110 2420
rect 394 2319 404 2371
rect 1388 2368 1398 2371
rect 6568 2368 6578 2371
rect 1388 2322 6578 2368
rect 1388 2319 1398 2322
rect 6568 2319 6578 2322
rect 7562 2319 7572 2371
rect 8076 2291 8122 2431
rect -169 2239 -159 2291
rect -107 2288 -97 2291
rect 8063 2288 8073 2291
rect -107 2242 8073 2288
rect -107 2239 -97 2242
rect 8063 2239 8073 2242
rect 8125 2239 8135 2291
rect -169 2005 -159 2181
rect -107 2005 -97 2181
rect 1889 2005 1899 2181
rect 1951 2005 1961 2181
rect 6005 2005 6015 2181
rect 6067 2005 6077 2181
rect 8063 2005 8073 2181
rect 8125 2005 8135 2181
rect -244 1958 -198 1993
rect -356 1946 -198 1958
rect -356 1912 -350 1946
rect -316 1912 -238 1946
rect -204 1912 -198 1946
rect -356 1900 -198 1912
rect 392 1889 1400 1906
rect 2450 1889 3458 1906
rect 3960 1889 4006 1993
rect 8164 1958 8210 1993
rect 8164 1946 8322 1958
rect 8164 1912 8170 1946
rect 8204 1912 8282 1946
rect 8316 1912 8322 1946
rect 4508 1889 5516 1906
rect 6566 1889 7574 1906
rect 8164 1900 8322 1912
rect -156 1843 8122 1889
rect -356 1820 -198 1832
rect -356 1786 -350 1820
rect -316 1786 -238 1820
rect -204 1786 -198 1820
rect -356 1774 -198 1786
rect -244 1739 -198 1774
rect -156 1739 -110 1843
rect 392 1826 1400 1843
rect 2450 1826 3458 1843
rect 4508 1826 5516 1843
rect 6566 1826 7574 1843
rect 8076 1727 8122 1843
rect 8164 1820 8322 1832
rect 8164 1786 8170 1820
rect 8204 1786 8282 1820
rect 8316 1786 8322 1820
rect 8164 1774 8322 1786
rect 8164 1735 8210 1774
rect 1889 1551 1899 1727
rect 1951 1551 1961 1727
rect 3947 1551 3957 1727
rect 4009 1551 4019 1727
rect 6005 1551 6015 1727
rect 6067 1551 6077 1727
rect -169 1438 -159 1490
rect -107 1487 -97 1490
rect 8063 1487 8073 1490
rect -107 1441 8073 1487
rect -107 1438 -97 1441
rect 8063 1438 8073 1441
rect 8125 1438 8135 1490
rect -156 1304 -110 1438
rect 394 1361 404 1413
rect 1388 1410 1398 1413
rect 6568 1410 6578 1413
rect 1388 1364 6578 1410
rect 1388 1361 1398 1364
rect 6568 1361 6578 1364
rect 7562 1361 7572 1413
rect 1889 1135 1899 1311
rect 1951 1135 1961 1311
rect 3947 1135 3957 1311
rect 4009 1135 4019 1311
rect 6005 1135 6015 1311
rect 6067 1135 6077 1311
rect 8076 1309 8122 1438
rect -244 1082 -198 1123
rect -244 1076 -166 1082
rect -244 1042 -212 1076
rect -178 1042 -166 1076
rect -244 1036 -166 1042
rect -224 1004 -166 1036
rect -224 970 -212 1004
rect -178 970 -166 1004
rect -224 964 -166 970
rect 1896 1004 1954 1135
rect 1896 970 1908 1004
rect 1942 970 1954 1004
rect 1896 964 1954 970
rect 6012 1004 6070 1135
rect 8164 1082 8210 1123
rect 6012 970 6024 1004
rect 6058 970 6070 1004
rect 6012 964 6070 970
rect 8132 1076 8210 1082
rect 8132 1042 8144 1076
rect 8178 1042 8210 1076
rect 8132 1036 8210 1042
rect 8132 1004 8190 1036
rect 8132 970 8144 1004
rect 8178 970 8190 1004
rect 8132 964 8190 970
<< via1 >>
rect 1899 2421 1951 2597
rect 3957 2421 4009 2597
rect 6015 2421 6067 2597
rect 404 2319 1388 2371
rect 6578 2319 7562 2371
rect -159 2239 -107 2291
rect 8073 2239 8125 2291
rect -159 2005 -107 2181
rect 1899 2005 1951 2181
rect 6015 2005 6067 2181
rect 8073 2005 8125 2181
rect 1899 1551 1951 1727
rect 3957 1551 4009 1727
rect 6015 1551 6067 1727
rect -159 1438 -107 1490
rect 8073 1438 8125 1490
rect 404 1361 1388 1413
rect 6578 1361 7562 1413
rect 1899 1135 1951 1311
rect 3957 1135 4009 1311
rect 6015 1135 6067 1311
<< metal2 >>
rect 1899 2597 1951 2607
rect 404 2373 1388 2383
rect 404 2307 1388 2317
rect -159 2291 -107 2301
rect -304 2239 -159 2291
rect -304 1490 -252 2239
rect -159 2229 -107 2239
rect -161 2181 -105 2191
rect -161 1995 -105 2005
rect 1899 2181 1951 2421
rect 3955 2597 4011 2607
rect 3955 2411 4011 2421
rect 6015 2597 6067 2607
rect 1899 1727 1951 2005
rect 6015 2181 6067 2421
rect 6578 2373 7562 2383
rect 6578 2307 7562 2317
rect 8073 2291 8125 2301
rect 8125 2239 8270 2291
rect 8073 2229 8125 2239
rect -159 1490 -107 1500
rect -304 1438 -159 1490
rect -159 1428 -107 1438
rect 404 1415 1388 1425
rect 404 1349 1388 1359
rect 1899 1311 1951 1551
rect 3955 1727 4011 1737
rect 3955 1541 4011 1551
rect 6015 1727 6067 2005
rect 8071 2181 8127 2191
rect 8071 1995 8127 2005
rect 1899 1125 1951 1135
rect 3955 1311 4011 1321
rect 3955 1125 4011 1135
rect 6015 1311 6067 1551
rect 8073 1490 8125 1500
rect 8218 1490 8270 2239
rect 8125 1438 8270 1490
rect 8073 1428 8125 1438
rect 6578 1415 7562 1425
rect 6578 1349 7562 1359
rect 6015 1125 6067 1135
<< via2 >>
rect 404 2371 1388 2373
rect 404 2319 1388 2371
rect 404 2317 1388 2319
rect -161 2005 -159 2181
rect -159 2005 -107 2181
rect -107 2005 -105 2181
rect 3955 2421 3957 2597
rect 3957 2421 4009 2597
rect 4009 2421 4011 2597
rect 6578 2371 7562 2373
rect 6578 2319 7562 2371
rect 6578 2317 7562 2319
rect 404 1413 1388 1415
rect 404 1361 1388 1413
rect 404 1359 1388 1361
rect 3955 1551 3957 1727
rect 3957 1551 4009 1727
rect 4009 1551 4011 1727
rect 8071 2005 8073 2181
rect 8073 2005 8125 2181
rect 8125 2005 8127 2181
rect 3955 1135 3957 1311
rect 3957 1135 4009 1311
rect 4009 1135 4011 1311
rect 6578 1413 7562 1415
rect 6578 1361 7562 1413
rect 6578 1359 7562 1361
<< metal3 >>
rect 3945 2597 4021 2602
rect 3941 2421 3951 2597
rect 4015 2421 4025 2597
rect 3945 2416 4021 2421
rect 394 2376 1398 2378
rect -312 2373 1398 2376
rect -312 2317 404 2373
rect 1388 2317 1398 2373
rect -312 2316 1398 2317
rect -312 1418 -252 2316
rect 394 2312 1398 2316
rect 6568 2375 7572 2378
rect 6568 2373 8278 2375
rect 6568 2317 6578 2373
rect 7562 2317 8278 2373
rect 6568 2315 8278 2317
rect 6568 2312 7572 2315
rect -171 2181 -95 2186
rect -171 2005 -161 2181
rect -105 2005 -95 2181
rect -171 2000 -95 2005
rect 8061 2181 8137 2186
rect 8061 2005 8071 2181
rect 8127 2005 8137 2181
rect 8061 2000 8137 2005
rect -163 1896 -103 2000
rect 8069 1896 8129 2000
rect -163 1836 8129 1896
rect 3953 1732 4013 1836
rect 3945 1727 4021 1732
rect 3945 1551 3955 1727
rect 4011 1551 4021 1727
rect 3945 1546 4021 1551
rect 394 1418 1398 1420
rect -312 1415 1398 1418
rect -312 1359 404 1415
rect 1388 1359 1398 1415
rect -312 1358 1398 1359
rect 394 1354 1398 1358
rect 6568 1417 7572 1420
rect 8218 1417 8278 2315
rect 6568 1415 8278 1417
rect 6568 1359 6578 1415
rect 7562 1359 8278 1415
rect 6568 1357 8278 1359
rect 6568 1354 7572 1357
rect 3945 1311 4021 1316
rect 3941 1135 3951 1311
rect 4015 1135 4025 1311
rect 3945 1130 4021 1135
<< via3 >>
rect 3951 2421 3955 2597
rect 3955 2421 4011 2597
rect 4011 2421 4015 2597
rect 3951 1135 3955 1311
rect 3955 1135 4011 1311
rect 4011 1135 4015 1311
<< metal4 >>
rect 3950 2597 4016 2598
rect 3950 2421 3951 2597
rect 4015 2421 4016 2597
rect 3950 2420 4016 2421
rect 3953 1312 4013 2420
rect 3950 1311 4016 1312
rect 3950 1135 3951 1311
rect 4015 1135 4016 1311
rect 3950 1134 4016 1135
use sky130_fd_pr__pfet_01v8_2XU96L  sky130_fd_pr__pfet_01v8_2XU96L_0
timestamp 1717000582
transform 1 0 -177 0 1 1223
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XU96L  sky130_fd_pr__pfet_01v8_2XU96L_1
timestamp 1717000582
transform 1 0 8143 0 1 2509
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XU96L  sky130_fd_pr__pfet_01v8_2XU96L_2
timestamp 1717000582
transform 1 0 8143 0 1 2093
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XU96L  sky130_fd_pr__pfet_01v8_2XU96L_3
timestamp 1717000582
transform 1 0 8143 0 1 1639
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XU96L  sky130_fd_pr__pfet_01v8_2XU96L_4
timestamp 1717000582
transform 1 0 8143 0 1 1223
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XU96L  sky130_fd_pr__pfet_01v8_2XU96L_5
timestamp 1717000582
transform 1 0 -177 0 1 2509
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XU96L  sky130_fd_pr__pfet_01v8_2XU96L_6
timestamp 1717000582
transform 1 0 -177 0 1 2093
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XU96L  sky130_fd_pr__pfet_01v8_2XU96L_7
timestamp 1717000582
transform 1 0 -177 0 1 1639
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_8WJJP2  sky130_fd_pr__pfet_01v8_8WJJP2_0
timestamp 1717071345
transform 1 0 3983 0 1 1675
box -4181 -198 4181 164
use sky130_fd_pr__pfet_01v8_8WJJP2  sky130_fd_pr__pfet_01v8_8WJJP2_1
timestamp 1717071345
transform 1 0 3983 0 1 1259
box -4181 -198 4181 164
use sky130_fd_pr__pfet_01v8_C2SJBD  sky130_fd_pr__pfet_01v8_C2SJBD_0
timestamp 1717071345
transform 1 0 3983 0 1 2473
box -4181 -164 4181 198
use sky130_fd_pr__pfet_01v8_C2SJBD  sky130_fd_pr__pfet_01v8_C2SJBD_1
timestamp 1717071345
transform 1 0 3983 0 1 2057
box -4181 -164 4181 198
<< labels >>
flabel metal2 8174 2266 8174 2266 0 FreeSans 160 0 0 0 D4
port 0 nsew
flabel viali 8160 2743 8160 2743 0 FreeSans 160 0 0 0 VDD
port 1 nsew
flabel metal3 8094 1928 8094 1928 0 FreeSans 160 0 0 0 D2
port 2 nsew
flabel metal1 8100 1776 8100 1776 0 FreeSans 160 0 0 0 D1
port 3 nsew
flabel metal4 3977 1420 3977 1420 0 FreeSans 160 0 0 0 D3
port 4 nsew
flabel metal3 7704 1397 7705 1397 0 FreeSans 160 0 0 0 G
port 5 nsew
<< end >>
