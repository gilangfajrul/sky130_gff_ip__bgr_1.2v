magic
tech sky130A
magscale 1 2
timestamp 1718865135
<< pwell >>
rect -782 -8202 782 8202
<< psubdiff >>
rect -746 8132 -650 8166
rect 650 8132 746 8166
rect -746 8070 -712 8132
rect 712 8070 746 8132
rect -746 -8132 -712 -8070
rect 712 -8132 746 -8070
rect -746 -8166 -650 -8132
rect 650 -8166 746 -8132
<< psubdiffcont >>
rect -650 8132 650 8166
rect -746 -8070 -712 8070
rect 712 -8070 746 8070
rect -650 -8166 650 -8132
<< xpolycontact >>
rect -616 7604 -546 8036
rect -616 5444 -546 5876
rect -450 7604 -380 8036
rect -450 5444 -380 5876
rect -284 7604 -214 8036
rect -284 5444 -214 5876
rect -118 7604 -48 8036
rect -118 5444 -48 5876
rect 48 7604 118 8036
rect 48 5444 118 5876
rect 214 7604 284 8036
rect 214 5444 284 5876
rect 380 7604 450 8036
rect 380 5444 450 5876
rect 546 7604 616 8036
rect 546 5444 616 5876
rect -616 4908 -546 5340
rect -616 2748 -546 3180
rect -450 4908 -380 5340
rect -450 2748 -380 3180
rect -284 4908 -214 5340
rect -284 2748 -214 3180
rect -118 4908 -48 5340
rect -118 2748 -48 3180
rect 48 4908 118 5340
rect 48 2748 118 3180
rect 214 4908 284 5340
rect 214 2748 284 3180
rect 380 4908 450 5340
rect 380 2748 450 3180
rect 546 4908 616 5340
rect 546 2748 616 3180
rect -616 2212 -546 2644
rect -616 52 -546 484
rect -450 2212 -380 2644
rect -450 52 -380 484
rect -284 2212 -214 2644
rect -284 52 -214 484
rect -118 2212 -48 2644
rect -118 52 -48 484
rect 48 2212 118 2644
rect 48 52 118 484
rect 214 2212 284 2644
rect 214 52 284 484
rect 380 2212 450 2644
rect 380 52 450 484
rect 546 2212 616 2644
rect 546 52 616 484
rect -616 -484 -546 -52
rect -616 -2644 -546 -2212
rect -450 -484 -380 -52
rect -450 -2644 -380 -2212
rect -284 -484 -214 -52
rect -284 -2644 -214 -2212
rect -118 -484 -48 -52
rect -118 -2644 -48 -2212
rect 48 -484 118 -52
rect 48 -2644 118 -2212
rect 214 -484 284 -52
rect 214 -2644 284 -2212
rect 380 -484 450 -52
rect 380 -2644 450 -2212
rect 546 -484 616 -52
rect 546 -2644 616 -2212
rect -616 -3180 -546 -2748
rect -616 -5340 -546 -4908
rect -450 -3180 -380 -2748
rect -450 -5340 -380 -4908
rect -284 -3180 -214 -2748
rect -284 -5340 -214 -4908
rect -118 -3180 -48 -2748
rect -118 -5340 -48 -4908
rect 48 -3180 118 -2748
rect 48 -5340 118 -4908
rect 214 -3180 284 -2748
rect 214 -5340 284 -4908
rect 380 -3180 450 -2748
rect 380 -5340 450 -4908
rect 546 -3180 616 -2748
rect 546 -5340 616 -4908
rect -616 -5876 -546 -5444
rect -616 -8036 -546 -7604
rect -450 -5876 -380 -5444
rect -450 -8036 -380 -7604
rect -284 -5876 -214 -5444
rect -284 -8036 -214 -7604
rect -118 -5876 -48 -5444
rect -118 -8036 -48 -7604
rect 48 -5876 118 -5444
rect 48 -8036 118 -7604
rect 214 -5876 284 -5444
rect 214 -8036 284 -7604
rect 380 -5876 450 -5444
rect 380 -8036 450 -7604
rect 546 -5876 616 -5444
rect 546 -8036 616 -7604
<< ppolyres >>
rect -616 5876 -546 7604
rect -450 5876 -380 7604
rect -284 5876 -214 7604
rect -118 5876 -48 7604
rect 48 5876 118 7604
rect 214 5876 284 7604
rect 380 5876 450 7604
rect 546 5876 616 7604
rect -616 3180 -546 4908
rect -450 3180 -380 4908
rect -284 3180 -214 4908
rect -118 3180 -48 4908
rect 48 3180 118 4908
rect 214 3180 284 4908
rect 380 3180 450 4908
rect 546 3180 616 4908
rect -616 484 -546 2212
rect -450 484 -380 2212
rect -284 484 -214 2212
rect -118 484 -48 2212
rect 48 484 118 2212
rect 214 484 284 2212
rect 380 484 450 2212
rect 546 484 616 2212
rect -616 -2212 -546 -484
rect -450 -2212 -380 -484
rect -284 -2212 -214 -484
rect -118 -2212 -48 -484
rect 48 -2212 118 -484
rect 214 -2212 284 -484
rect 380 -2212 450 -484
rect 546 -2212 616 -484
rect -616 -4908 -546 -3180
rect -450 -4908 -380 -3180
rect -284 -4908 -214 -3180
rect -118 -4908 -48 -3180
rect 48 -4908 118 -3180
rect 214 -4908 284 -3180
rect 380 -4908 450 -3180
rect 546 -4908 616 -3180
rect -616 -7604 -546 -5876
rect -450 -7604 -380 -5876
rect -284 -7604 -214 -5876
rect -118 -7604 -48 -5876
rect 48 -7604 118 -5876
rect 214 -7604 284 -5876
rect 380 -7604 450 -5876
rect 546 -7604 616 -5876
<< locali >>
rect -666 8132 -650 8166
rect 650 8132 666 8166
rect -746 8070 -712 8086
rect 712 8070 746 8086
rect -746 -8086 -712 -8070
rect 712 -8086 746 -8070
rect -666 -8166 -650 -8132
rect 650 -8166 666 -8132
<< viali >>
rect -600 7621 -562 8018
rect -434 7621 -396 8018
rect -268 7621 -230 8018
rect -102 7621 -64 8018
rect 64 7621 102 8018
rect 230 7621 268 8018
rect 396 7621 434 8018
rect 562 7621 600 8018
rect -600 5462 -562 5859
rect -434 5462 -396 5859
rect -268 5462 -230 5859
rect -102 5462 -64 5859
rect 64 5462 102 5859
rect 230 5462 268 5859
rect 396 5462 434 5859
rect 562 5462 600 5859
rect -600 4925 -562 5322
rect -434 4925 -396 5322
rect -268 4925 -230 5322
rect -102 4925 -64 5322
rect 64 4925 102 5322
rect 230 4925 268 5322
rect 396 4925 434 5322
rect 562 4925 600 5322
rect -600 2766 -562 3163
rect -434 2766 -396 3163
rect -268 2766 -230 3163
rect -102 2766 -64 3163
rect 64 2766 102 3163
rect 230 2766 268 3163
rect 396 2766 434 3163
rect 562 2766 600 3163
rect -600 2229 -562 2626
rect -434 2229 -396 2626
rect -268 2229 -230 2626
rect -102 2229 -64 2626
rect 64 2229 102 2626
rect 230 2229 268 2626
rect 396 2229 434 2626
rect 562 2229 600 2626
rect -600 70 -562 467
rect -434 70 -396 467
rect -268 70 -230 467
rect -102 70 -64 467
rect 64 70 102 467
rect 230 70 268 467
rect 396 70 434 467
rect 562 70 600 467
rect -600 -467 -562 -70
rect -434 -467 -396 -70
rect -268 -467 -230 -70
rect -102 -467 -64 -70
rect 64 -467 102 -70
rect 230 -467 268 -70
rect 396 -467 434 -70
rect 562 -467 600 -70
rect -600 -2626 -562 -2229
rect -434 -2626 -396 -2229
rect -268 -2626 -230 -2229
rect -102 -2626 -64 -2229
rect 64 -2626 102 -2229
rect 230 -2626 268 -2229
rect 396 -2626 434 -2229
rect 562 -2626 600 -2229
rect -600 -3163 -562 -2766
rect -434 -3163 -396 -2766
rect -268 -3163 -230 -2766
rect -102 -3163 -64 -2766
rect 64 -3163 102 -2766
rect 230 -3163 268 -2766
rect 396 -3163 434 -2766
rect 562 -3163 600 -2766
rect -600 -5322 -562 -4925
rect -434 -5322 -396 -4925
rect -268 -5322 -230 -4925
rect -102 -5322 -64 -4925
rect 64 -5322 102 -4925
rect 230 -5322 268 -4925
rect 396 -5322 434 -4925
rect 562 -5322 600 -4925
rect -600 -5859 -562 -5462
rect -434 -5859 -396 -5462
rect -268 -5859 -230 -5462
rect -102 -5859 -64 -5462
rect 64 -5859 102 -5462
rect 230 -5859 268 -5462
rect 396 -5859 434 -5462
rect 562 -5859 600 -5462
rect -600 -8018 -562 -7621
rect -434 -8018 -396 -7621
rect -268 -8018 -230 -7621
rect -102 -8018 -64 -7621
rect 64 -8018 102 -7621
rect 230 -8018 268 -7621
rect 396 -8018 434 -7621
rect 562 -8018 600 -7621
<< metal1 >>
rect -606 8018 -556 8030
rect -606 7621 -600 8018
rect -562 7621 -556 8018
rect -606 7609 -556 7621
rect -440 8018 -390 8030
rect -440 7621 -434 8018
rect -396 7621 -390 8018
rect -440 7609 -390 7621
rect -274 8018 -224 8030
rect -274 7621 -268 8018
rect -230 7621 -224 8018
rect -274 7609 -224 7621
rect -108 8018 -58 8030
rect -108 7621 -102 8018
rect -64 7621 -58 8018
rect -108 7609 -58 7621
rect 58 8018 108 8030
rect 58 7621 64 8018
rect 102 7621 108 8018
rect 58 7609 108 7621
rect 224 8018 274 8030
rect 224 7621 230 8018
rect 268 7621 274 8018
rect 224 7609 274 7621
rect 390 8018 440 8030
rect 390 7621 396 8018
rect 434 7621 440 8018
rect 390 7609 440 7621
rect 556 8018 606 8030
rect 556 7621 562 8018
rect 600 7621 606 8018
rect 556 7609 606 7621
rect -606 5859 -556 5871
rect -606 5462 -600 5859
rect -562 5462 -556 5859
rect -606 5450 -556 5462
rect -440 5859 -390 5871
rect -440 5462 -434 5859
rect -396 5462 -390 5859
rect -440 5450 -390 5462
rect -274 5859 -224 5871
rect -274 5462 -268 5859
rect -230 5462 -224 5859
rect -274 5450 -224 5462
rect -108 5859 -58 5871
rect -108 5462 -102 5859
rect -64 5462 -58 5859
rect -108 5450 -58 5462
rect 58 5859 108 5871
rect 58 5462 64 5859
rect 102 5462 108 5859
rect 58 5450 108 5462
rect 224 5859 274 5871
rect 224 5462 230 5859
rect 268 5462 274 5859
rect 224 5450 274 5462
rect 390 5859 440 5871
rect 390 5462 396 5859
rect 434 5462 440 5859
rect 390 5450 440 5462
rect 556 5859 606 5871
rect 556 5462 562 5859
rect 600 5462 606 5859
rect 556 5450 606 5462
rect -606 5322 -556 5334
rect -606 4925 -600 5322
rect -562 4925 -556 5322
rect -606 4913 -556 4925
rect -440 5322 -390 5334
rect -440 4925 -434 5322
rect -396 4925 -390 5322
rect -440 4913 -390 4925
rect -274 5322 -224 5334
rect -274 4925 -268 5322
rect -230 4925 -224 5322
rect -274 4913 -224 4925
rect -108 5322 -58 5334
rect -108 4925 -102 5322
rect -64 4925 -58 5322
rect -108 4913 -58 4925
rect 58 5322 108 5334
rect 58 4925 64 5322
rect 102 4925 108 5322
rect 58 4913 108 4925
rect 224 5322 274 5334
rect 224 4925 230 5322
rect 268 4925 274 5322
rect 224 4913 274 4925
rect 390 5322 440 5334
rect 390 4925 396 5322
rect 434 4925 440 5322
rect 390 4913 440 4925
rect 556 5322 606 5334
rect 556 4925 562 5322
rect 600 4925 606 5322
rect 556 4913 606 4925
rect -606 3163 -556 3175
rect -606 2766 -600 3163
rect -562 2766 -556 3163
rect -606 2754 -556 2766
rect -440 3163 -390 3175
rect -440 2766 -434 3163
rect -396 2766 -390 3163
rect -440 2754 -390 2766
rect -274 3163 -224 3175
rect -274 2766 -268 3163
rect -230 2766 -224 3163
rect -274 2754 -224 2766
rect -108 3163 -58 3175
rect -108 2766 -102 3163
rect -64 2766 -58 3163
rect -108 2754 -58 2766
rect 58 3163 108 3175
rect 58 2766 64 3163
rect 102 2766 108 3163
rect 58 2754 108 2766
rect 224 3163 274 3175
rect 224 2766 230 3163
rect 268 2766 274 3163
rect 224 2754 274 2766
rect 390 3163 440 3175
rect 390 2766 396 3163
rect 434 2766 440 3163
rect 390 2754 440 2766
rect 556 3163 606 3175
rect 556 2766 562 3163
rect 600 2766 606 3163
rect 556 2754 606 2766
rect -606 2626 -556 2638
rect -606 2229 -600 2626
rect -562 2229 -556 2626
rect -606 2217 -556 2229
rect -440 2626 -390 2638
rect -440 2229 -434 2626
rect -396 2229 -390 2626
rect -440 2217 -390 2229
rect -274 2626 -224 2638
rect -274 2229 -268 2626
rect -230 2229 -224 2626
rect -274 2217 -224 2229
rect -108 2626 -58 2638
rect -108 2229 -102 2626
rect -64 2229 -58 2626
rect -108 2217 -58 2229
rect 58 2626 108 2638
rect 58 2229 64 2626
rect 102 2229 108 2626
rect 58 2217 108 2229
rect 224 2626 274 2638
rect 224 2229 230 2626
rect 268 2229 274 2626
rect 224 2217 274 2229
rect 390 2626 440 2638
rect 390 2229 396 2626
rect 434 2229 440 2626
rect 390 2217 440 2229
rect 556 2626 606 2638
rect 556 2229 562 2626
rect 600 2229 606 2626
rect 556 2217 606 2229
rect -606 467 -556 479
rect -606 70 -600 467
rect -562 70 -556 467
rect -606 58 -556 70
rect -440 467 -390 479
rect -440 70 -434 467
rect -396 70 -390 467
rect -440 58 -390 70
rect -274 467 -224 479
rect -274 70 -268 467
rect -230 70 -224 467
rect -274 58 -224 70
rect -108 467 -58 479
rect -108 70 -102 467
rect -64 70 -58 467
rect -108 58 -58 70
rect 58 467 108 479
rect 58 70 64 467
rect 102 70 108 467
rect 58 58 108 70
rect 224 467 274 479
rect 224 70 230 467
rect 268 70 274 467
rect 224 58 274 70
rect 390 467 440 479
rect 390 70 396 467
rect 434 70 440 467
rect 390 58 440 70
rect 556 467 606 479
rect 556 70 562 467
rect 600 70 606 467
rect 556 58 606 70
rect -606 -70 -556 -58
rect -606 -467 -600 -70
rect -562 -467 -556 -70
rect -606 -479 -556 -467
rect -440 -70 -390 -58
rect -440 -467 -434 -70
rect -396 -467 -390 -70
rect -440 -479 -390 -467
rect -274 -70 -224 -58
rect -274 -467 -268 -70
rect -230 -467 -224 -70
rect -274 -479 -224 -467
rect -108 -70 -58 -58
rect -108 -467 -102 -70
rect -64 -467 -58 -70
rect -108 -479 -58 -467
rect 58 -70 108 -58
rect 58 -467 64 -70
rect 102 -467 108 -70
rect 58 -479 108 -467
rect 224 -70 274 -58
rect 224 -467 230 -70
rect 268 -467 274 -70
rect 224 -479 274 -467
rect 390 -70 440 -58
rect 390 -467 396 -70
rect 434 -467 440 -70
rect 390 -479 440 -467
rect 556 -70 606 -58
rect 556 -467 562 -70
rect 600 -467 606 -70
rect 556 -479 606 -467
rect -606 -2229 -556 -2217
rect -606 -2626 -600 -2229
rect -562 -2626 -556 -2229
rect -606 -2638 -556 -2626
rect -440 -2229 -390 -2217
rect -440 -2626 -434 -2229
rect -396 -2626 -390 -2229
rect -440 -2638 -390 -2626
rect -274 -2229 -224 -2217
rect -274 -2626 -268 -2229
rect -230 -2626 -224 -2229
rect -274 -2638 -224 -2626
rect -108 -2229 -58 -2217
rect -108 -2626 -102 -2229
rect -64 -2626 -58 -2229
rect -108 -2638 -58 -2626
rect 58 -2229 108 -2217
rect 58 -2626 64 -2229
rect 102 -2626 108 -2229
rect 58 -2638 108 -2626
rect 224 -2229 274 -2217
rect 224 -2626 230 -2229
rect 268 -2626 274 -2229
rect 224 -2638 274 -2626
rect 390 -2229 440 -2217
rect 390 -2626 396 -2229
rect 434 -2626 440 -2229
rect 390 -2638 440 -2626
rect 556 -2229 606 -2217
rect 556 -2626 562 -2229
rect 600 -2626 606 -2229
rect 556 -2638 606 -2626
rect -606 -2766 -556 -2754
rect -606 -3163 -600 -2766
rect -562 -3163 -556 -2766
rect -606 -3175 -556 -3163
rect -440 -2766 -390 -2754
rect -440 -3163 -434 -2766
rect -396 -3163 -390 -2766
rect -440 -3175 -390 -3163
rect -274 -2766 -224 -2754
rect -274 -3163 -268 -2766
rect -230 -3163 -224 -2766
rect -274 -3175 -224 -3163
rect -108 -2766 -58 -2754
rect -108 -3163 -102 -2766
rect -64 -3163 -58 -2766
rect -108 -3175 -58 -3163
rect 58 -2766 108 -2754
rect 58 -3163 64 -2766
rect 102 -3163 108 -2766
rect 58 -3175 108 -3163
rect 224 -2766 274 -2754
rect 224 -3163 230 -2766
rect 268 -3163 274 -2766
rect 224 -3175 274 -3163
rect 390 -2766 440 -2754
rect 390 -3163 396 -2766
rect 434 -3163 440 -2766
rect 390 -3175 440 -3163
rect 556 -2766 606 -2754
rect 556 -3163 562 -2766
rect 600 -3163 606 -2766
rect 556 -3175 606 -3163
rect -606 -4925 -556 -4913
rect -606 -5322 -600 -4925
rect -562 -5322 -556 -4925
rect -606 -5334 -556 -5322
rect -440 -4925 -390 -4913
rect -440 -5322 -434 -4925
rect -396 -5322 -390 -4925
rect -440 -5334 -390 -5322
rect -274 -4925 -224 -4913
rect -274 -5322 -268 -4925
rect -230 -5322 -224 -4925
rect -274 -5334 -224 -5322
rect -108 -4925 -58 -4913
rect -108 -5322 -102 -4925
rect -64 -5322 -58 -4925
rect -108 -5334 -58 -5322
rect 58 -4925 108 -4913
rect 58 -5322 64 -4925
rect 102 -5322 108 -4925
rect 58 -5334 108 -5322
rect 224 -4925 274 -4913
rect 224 -5322 230 -4925
rect 268 -5322 274 -4925
rect 224 -5334 274 -5322
rect 390 -4925 440 -4913
rect 390 -5322 396 -4925
rect 434 -5322 440 -4925
rect 390 -5334 440 -5322
rect 556 -4925 606 -4913
rect 556 -5322 562 -4925
rect 600 -5322 606 -4925
rect 556 -5334 606 -5322
rect -606 -5462 -556 -5450
rect -606 -5859 -600 -5462
rect -562 -5859 -556 -5462
rect -606 -5871 -556 -5859
rect -440 -5462 -390 -5450
rect -440 -5859 -434 -5462
rect -396 -5859 -390 -5462
rect -440 -5871 -390 -5859
rect -274 -5462 -224 -5450
rect -274 -5859 -268 -5462
rect -230 -5859 -224 -5462
rect -274 -5871 -224 -5859
rect -108 -5462 -58 -5450
rect -108 -5859 -102 -5462
rect -64 -5859 -58 -5462
rect -108 -5871 -58 -5859
rect 58 -5462 108 -5450
rect 58 -5859 64 -5462
rect 102 -5859 108 -5462
rect 58 -5871 108 -5859
rect 224 -5462 274 -5450
rect 224 -5859 230 -5462
rect 268 -5859 274 -5462
rect 224 -5871 274 -5859
rect 390 -5462 440 -5450
rect 390 -5859 396 -5462
rect 434 -5859 440 -5462
rect 390 -5871 440 -5859
rect 556 -5462 606 -5450
rect 556 -5859 562 -5462
rect 600 -5859 606 -5462
rect 556 -5871 606 -5859
rect -606 -7621 -556 -7609
rect -606 -8018 -600 -7621
rect -562 -8018 -556 -7621
rect -606 -8030 -556 -8018
rect -440 -7621 -390 -7609
rect -440 -8018 -434 -7621
rect -396 -8018 -390 -7621
rect -440 -8030 -390 -8018
rect -274 -7621 -224 -7609
rect -274 -8018 -268 -7621
rect -230 -8018 -224 -7621
rect -274 -8030 -224 -8018
rect -108 -7621 -58 -7609
rect -108 -8018 -102 -7621
rect -64 -8018 -58 -7621
rect -108 -8030 -58 -8018
rect 58 -7621 108 -7609
rect 58 -8018 64 -7621
rect 102 -8018 108 -7621
rect 58 -8030 108 -8018
rect 224 -7621 274 -7609
rect 224 -8018 230 -7621
rect 268 -8018 274 -7621
rect 224 -8030 274 -8018
rect 390 -7621 440 -7609
rect 390 -8018 396 -7621
rect 434 -8018 440 -7621
rect 390 -8030 440 -8018
rect 556 -7621 606 -7609
rect 556 -8018 562 -7621
rect 600 -8018 606 -7621
rect 556 -8030 606 -8018
<< properties >>
string FIXED_BBOX -729 -8149 729 8149
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.350 l 8.8 m 6 nx 8 wmin 0.350 lmin 0.50 rho 319.8 val 9.153k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 0 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
