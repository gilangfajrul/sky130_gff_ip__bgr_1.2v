magic
tech sky130A
magscale 1 2
timestamp 1717768441
<< error_p >>
rect -29 245 29 251
rect -29 211 -17 245
rect -29 205 29 211
<< nwell >>
rect -109 -298 109 264
<< pmos >>
rect -15 -236 15 164
<< pdiff >>
rect -73 152 -15 164
rect -73 -224 -61 152
rect -27 -224 -15 152
rect -73 -236 -15 -224
rect 15 152 73 164
rect 15 -224 27 152
rect 61 -224 73 152
rect 15 -236 73 -224
<< pdiffc >>
rect -61 -224 -27 152
rect 27 -224 61 152
<< poly >>
rect -33 245 33 261
rect -33 211 -17 245
rect 17 211 33 245
rect -33 195 33 211
rect -15 164 15 195
rect -15 -262 15 -236
<< polycont >>
rect -17 211 17 245
<< locali >>
rect -33 211 -17 245
rect 17 211 33 245
rect -61 152 -27 168
rect -61 -240 -27 -224
rect 27 152 61 168
rect 27 -240 61 -224
<< viali >>
rect -17 211 17 245
rect -61 -224 -27 152
rect 27 -224 61 152
<< metal1 >>
rect -29 245 29 251
rect -29 211 -17 245
rect 17 211 29 245
rect -29 205 29 211
rect -67 152 -21 164
rect -67 -224 -61 152
rect -27 -224 -21 152
rect -67 -236 -21 -224
rect 21 152 67 164
rect 21 -224 27 152
rect 61 -224 67 152
rect 21 -236 67 -224
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
