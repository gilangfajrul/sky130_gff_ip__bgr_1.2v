magic
tech sky130A
magscale 1 2
timestamp 1717421032
<< nwell >>
rect -2123 -198 2123 164
<< pmos >>
rect -2029 -136 -29 64
rect 29 -136 2029 64
<< pdiff >>
rect -2087 52 -2029 64
rect -2087 -124 -2075 52
rect -2041 -124 -2029 52
rect -2087 -136 -2029 -124
rect -29 52 29 64
rect -29 -124 -17 52
rect 17 -124 29 52
rect -29 -136 29 -124
rect 2029 52 2087 64
rect 2029 -124 2041 52
rect 2075 -124 2087 52
rect 2029 -136 2087 -124
<< pdiffc >>
rect -2075 -124 -2041 52
rect -17 -124 17 52
rect 2041 -124 2075 52
<< poly >>
rect -1537 145 -521 161
rect -1537 128 -1521 145
rect -2029 111 -1521 128
rect -537 128 -521 145
rect 521 145 1537 161
rect 521 128 537 145
rect -537 111 -29 128
rect -2029 64 -29 111
rect 29 111 537 128
rect 1521 128 1537 145
rect 1521 111 2029 128
rect 29 64 2029 111
rect -2029 -162 -29 -136
rect 29 -162 2029 -136
<< polycont >>
rect -1521 111 -537 145
rect 537 111 1521 145
<< locali >>
rect -1537 111 -1521 145
rect -537 111 -521 145
rect 521 111 537 145
rect 1521 111 1537 145
rect -2075 52 -2041 68
rect -2075 -140 -2041 -124
rect -17 52 17 68
rect -17 -140 17 -124
rect 2041 52 2075 68
rect 2041 -140 2075 -124
<< viali >>
rect -1521 111 -537 145
rect 537 111 1521 145
rect -2075 -124 -2041 52
rect -17 -124 17 52
rect 2041 -124 2075 52
<< metal1 >>
rect -1533 145 -525 151
rect -1533 111 -1521 145
rect -537 111 -525 145
rect -1533 105 -525 111
rect 525 145 1533 151
rect 525 111 537 145
rect 1521 111 1533 145
rect 525 105 1533 111
rect -2081 52 -2035 64
rect -2081 -124 -2075 52
rect -2041 -124 -2035 52
rect -2081 -136 -2035 -124
rect -23 52 23 64
rect -23 -124 -17 52
rect 17 -124 23 52
rect -23 -136 23 -124
rect 2035 52 2081 64
rect 2035 -124 2041 52
rect 2075 -124 2081 52
rect 2035 -136 2081 -124
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 10 m 1 nf 2 diffcov 100 polycov 50 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
