magic
tech sky130A
magscale 1 2
timestamp 1716993797
<< dnwell >>
rect -244 -407 8430 1175
<< nwell >>
rect -357 -510 8543 1278
<< pmos >>
rect 589 875 1425 879
<< nsubdiff >>
rect -321 1208 -261 1242
rect 8447 1208 8507 1242
rect -321 1182 -287 1208
rect 8473 1182 8507 1208
rect -321 -440 -287 -414
rect 8473 -440 8507 -414
rect -321 -474 -261 -440
rect 8447 -474 8507 -440
<< nsubdiffcont >>
rect -261 1208 8447 1242
rect -321 -414 -287 1182
rect 8473 -414 8507 1182
rect -261 -474 8447 -440
<< poly >>
rect -170 1095 -52 1148
rect -82 1075 -52 1095
rect 8238 1095 8356 1148
rect 8238 1075 8268 1095
rect 589 879 1425 887
rect 589 795 1425 875
rect 2651 795 3477 875
rect 4709 795 5535 875
rect 6771 795 7597 875
rect -82 461 -52 481
rect -170 408 -52 461
rect 593 414 1419 481
rect 2651 414 3477 481
rect 4709 414 5535 481
rect 6767 414 7593 481
rect 8238 461 8268 481
rect 8238 408 8356 461
rect -170 307 -52 360
rect -82 287 -52 307
rect 593 287 1419 354
rect 2651 307 3477 354
rect 4709 306 5535 354
rect 6767 287 7593 354
rect 8238 312 8356 360
rect 8260 307 8356 312
rect 589 -81 1425 -27
rect 2651 -81 3477 -27
rect 4709 -81 5535 -27
rect 6771 -81 7597 -27
rect 589 -107 2006 -81
rect 2064 -107 4064 -81
rect 4124 -107 6122 -81
rect 6180 -107 7597 -81
rect 8238 -107 8268 -81
rect -82 -327 -52 -307
rect -170 -380 -52 -327
rect 8238 -327 8268 -307
rect 8238 -380 8356 -327
<< locali >>
rect -321 1208 -261 1242
rect 8447 1208 8507 1242
rect -321 1182 -287 1208
rect 8473 1182 8507 1208
rect -128 1075 -94 1102
rect 8280 1075 8314 1102
rect -128 454 -94 481
rect 8280 454 8314 481
rect -128 287 -94 314
rect 8280 278 8314 314
rect 2018 -107 2052 -103
rect 6134 -107 6168 -103
rect 8192 -107 8226 -103
rect 8280 -107 8314 -103
rect -128 -334 -94 -307
rect 8280 -334 8314 -307
rect -321 -440 -287 -414
rect 8473 -440 8507 -414
rect -321 -474 -261 -440
rect 8447 -474 8507 -440
<< viali >>
rect 2012 1208 2058 1242
rect 6128 1208 6174 1242
rect -158 1102 -86 1138
rect 4067 1113 4119 1165
rect 8272 1102 8344 1138
rect 606 815 1406 849
rect 2664 815 3464 849
rect 4722 815 5522 849
rect 6784 815 7584 849
rect -158 418 -86 454
rect 594 415 1418 455
rect 2652 415 3476 455
rect 4710 415 5534 455
rect 6768 415 7592 455
rect 8272 418 8344 454
rect -158 314 -86 350
rect 594 313 1418 353
rect 2652 313 3476 353
rect 4710 313 5534 353
rect 6768 313 7592 353
rect 8272 314 8344 350
rect 606 -81 1406 -47
rect 2664 -81 3464 -47
rect 4722 -81 5522 -47
rect 6784 -81 7584 -47
rect -158 -370 -86 -334
rect 4067 -397 4119 -345
rect 8272 -370 8344 -334
rect 2012 -474 2058 -440
rect 6128 -474 6174 -440
<< metal1 >>
rect 2000 1242 2070 1248
rect 2000 1208 2012 1242
rect 2058 1208 2070 1242
rect 2000 1202 2070 1208
rect 6116 1242 6186 1248
rect 6116 1208 6128 1242
rect 6174 1208 6186 1242
rect 6116 1202 6186 1208
rect -170 1138 -74 1144
rect -170 1102 -158 1138
rect -86 1102 -74 1138
rect -170 1095 -74 1102
rect -134 1075 -88 1095
rect -46 1063 0 1075
rect 2012 1063 2058 1202
rect 4055 1165 4131 1171
rect 4055 1113 4067 1165
rect 4119 1113 4131 1165
rect 4055 1107 4131 1113
rect -46 887 -40 1063
rect -6 887 0 1063
rect 1999 887 2009 1063
rect 2061 887 2071 1063
rect 4070 1057 4116 1107
rect 6128 1063 6174 1202
rect 8260 1138 8356 1144
rect 8260 1102 8272 1138
rect 8344 1102 8356 1138
rect 8260 1095 8356 1102
rect 8274 1075 8320 1095
rect 6115 887 6125 1063
rect 6177 887 6187 1063
rect -134 824 -88 878
rect -46 824 0 887
rect -244 778 0 824
rect 594 806 606 858
rect 1406 806 1418 858
rect 2652 806 2664 858
rect 3464 806 3476 858
rect 4710 806 4722 858
rect 5522 806 5534 858
rect 6772 806 6784 858
rect 7584 806 7596 858
rect 8186 824 8232 875
rect 8274 824 8320 877
rect 8186 778 8430 824
rect -244 732 8430 778
rect -244 36 -198 732
rect -59 493 -49 669
rect 3 493 13 669
rect 1999 493 2009 669
rect 2061 493 2071 669
rect 6115 493 6125 669
rect 6177 493 6187 669
rect 8173 493 8183 669
rect 8235 493 8245 669
rect -134 463 -88 481
rect -46 463 0 486
rect -134 461 0 463
rect -170 454 0 461
rect -170 418 -158 454
rect -86 435 0 454
rect 582 455 1430 461
rect -86 418 -74 435
rect -170 412 -74 418
rect 582 415 594 455
rect 1418 415 1430 455
rect 582 407 1430 415
rect 2640 455 3488 461
rect 2640 415 2652 455
rect 3476 415 3488 455
rect 2640 407 3488 415
rect 4070 407 4116 481
rect 8186 463 8232 493
rect 8274 463 8320 481
rect 8186 461 8320 463
rect 4698 455 5546 461
rect 4698 415 4710 455
rect 5534 415 5546 455
rect 4698 407 5546 415
rect 6756 455 7604 461
rect 6756 415 6768 455
rect 7592 415 7604 455
rect 8186 454 8356 461
rect 8186 435 8272 454
rect 6756 407 7604 415
rect 8260 418 8272 435
rect 8344 418 8356 454
rect 8260 412 8356 418
rect -46 361 8232 407
rect -46 356 0 361
rect -170 350 0 356
rect -170 314 -158 350
rect -86 314 0 350
rect -170 307 0 314
rect 582 353 1430 361
rect 582 313 594 353
rect 1418 313 1430 353
rect 582 307 1430 313
rect 2640 353 3488 361
rect 2640 313 2652 353
rect 3476 313 3488 353
rect 2640 307 3488 313
rect 4698 353 5546 361
rect 4698 313 4710 353
rect 5534 313 5546 353
rect 4698 307 5546 313
rect 6756 353 7604 361
rect 6756 313 6768 353
rect 7592 313 7604 353
rect 6756 307 7604 313
rect 8186 356 8232 361
rect 8186 350 8356 356
rect 8186 314 8272 350
rect 8344 314 8356 350
rect 8186 307 8356 314
rect -134 287 -88 307
rect -46 285 0 307
rect 8186 280 8232 307
rect 8274 279 8320 307
rect 8280 278 8314 279
rect 1999 99 2009 275
rect 2061 99 2071 275
rect 4057 99 4067 275
rect 4119 99 4129 275
rect 6115 99 6125 275
rect 6177 99 6187 275
rect 8384 36 8430 732
rect -244 -10 8430 36
rect -244 -56 0 -10
rect -134 -107 -88 -56
rect -46 -119 0 -56
rect 594 -90 606 -38
rect 1406 -90 1418 -38
rect 2652 -90 2664 -38
rect 3464 -90 3476 -38
rect 4710 -90 4722 -38
rect 5522 -90 5534 -38
rect 6772 -90 6784 -38
rect 7584 -90 7596 -38
rect 8186 -56 8430 -10
rect 8186 -107 8232 -56
rect 8274 -109 8320 -56
rect -46 -295 -40 -119
rect -6 -295 0 -119
rect 1999 -295 2009 -119
rect 2061 -295 2071 -119
rect 6115 -295 6125 -119
rect 6177 -295 6187 -119
rect -46 -307 0 -295
rect -134 -327 -88 -307
rect -170 -334 -74 -327
rect -170 -370 -158 -334
rect -86 -370 -74 -334
rect -170 -376 -74 -370
rect 2012 -434 2058 -307
rect 4070 -339 4116 -307
rect 4055 -345 4131 -339
rect 4055 -397 4067 -345
rect 4119 -397 4131 -345
rect 4055 -403 4131 -397
rect 6128 -434 6174 -307
rect 8274 -327 8320 -307
rect 8260 -334 8356 -327
rect 8260 -370 8272 -334
rect 8344 -370 8356 -334
rect 8260 -376 8356 -370
rect 2000 -440 2070 -434
rect 2000 -474 2012 -440
rect 2058 -474 2070 -440
rect 2000 -480 2070 -474
rect 6116 -440 6186 -434
rect 6116 -474 6128 -440
rect 6174 -474 6186 -440
rect 6116 -480 6186 -474
<< via1 >>
rect 4067 1113 4119 1165
rect 2009 887 2061 1063
rect 6125 887 6177 1063
rect 606 849 1406 858
rect 606 815 1406 849
rect 606 806 1406 815
rect 2664 849 3464 858
rect 2664 815 3464 849
rect 2664 806 3464 815
rect 4722 849 5522 858
rect 4722 815 5522 849
rect 4722 806 5522 815
rect 6784 849 7584 858
rect 6784 815 7584 849
rect 6784 806 7584 815
rect -49 493 3 669
rect 2009 493 2061 669
rect 6125 493 6177 669
rect 8183 493 8235 669
rect 2009 99 2061 275
rect 4067 99 4119 275
rect 6125 99 6177 275
rect 606 -47 1406 -38
rect 606 -81 1406 -47
rect 606 -90 1406 -81
rect 2664 -47 3464 -38
rect 2664 -81 3464 -47
rect 2664 -90 3464 -81
rect 4722 -47 5522 -38
rect 4722 -81 5522 -47
rect 4722 -90 5522 -81
rect 6784 -47 7584 -38
rect 6784 -81 7584 -47
rect 6784 -90 7584 -81
rect 2009 -295 2061 -119
rect 6125 -295 6177 -119
rect 4067 -397 4119 -345
<< metal2 >>
rect 4067 1165 4119 1175
rect -244 1113 4067 1165
rect 4119 1113 8430 1165
rect -244 -345 -198 1113
rect 4067 1103 4119 1113
rect 2007 1063 2063 1073
rect 2007 877 2063 887
rect 6123 1063 6179 1073
rect 6123 877 6179 887
rect 606 860 1406 870
rect 2664 858 3464 868
rect 1406 806 2664 849
rect 4722 858 5522 868
rect 3464 806 4722 849
rect 6784 860 7584 870
rect 5522 806 6784 849
rect 1406 804 6784 806
rect 606 796 7584 804
rect 606 794 1406 796
rect 6784 794 7584 796
rect -49 669 3 679
rect -49 410 3 493
rect 2007 669 2063 679
rect 2007 483 2063 493
rect 6123 669 6179 679
rect 6123 483 6179 493
rect 8183 669 8235 679
rect 8183 410 8235 493
rect -49 358 8235 410
rect 2007 275 2063 285
rect 2007 89 2063 99
rect 4067 275 4119 358
rect 4067 89 4119 99
rect 6123 275 6179 285
rect 6123 89 6179 99
rect 606 -28 1406 -26
rect 6784 -28 7584 -26
rect 606 -36 7584 -28
rect 1406 -38 6784 -36
rect 1406 -81 2664 -38
rect 606 -102 1406 -92
rect 3464 -81 4722 -38
rect 2664 -100 3464 -90
rect 5522 -81 6784 -38
rect 4722 -100 5522 -90
rect 6784 -102 7584 -92
rect 2007 -119 2063 -109
rect 2007 -305 2063 -295
rect 6123 -119 6179 -109
rect 6123 -305 6179 -295
rect 4067 -345 4119 -335
rect 8384 -345 8430 1113
rect -244 -397 4067 -345
rect 4119 -397 8430 -345
rect 4067 -407 4119 -397
<< via2 >>
rect 2007 887 2009 1063
rect 2009 887 2061 1063
rect 2061 887 2063 1063
rect 6123 887 6125 1063
rect 6125 887 6177 1063
rect 6177 887 6179 1063
rect 606 858 1406 860
rect 606 806 1406 858
rect 6784 858 7584 860
rect 6784 806 7584 858
rect 606 804 1406 806
rect 6784 804 7584 806
rect 2007 493 2009 669
rect 2009 493 2061 669
rect 2061 493 2063 669
rect 6123 493 6125 669
rect 6125 493 6177 669
rect 6177 493 6179 669
rect 2007 99 2009 275
rect 2009 99 2061 275
rect 2061 99 2063 275
rect 6123 99 6125 275
rect 6125 99 6177 275
rect 6177 99 6179 275
rect 606 -38 1406 -36
rect 6784 -38 7584 -36
rect 606 -90 1406 -38
rect 606 -92 1406 -90
rect 6784 -90 7584 -38
rect 6784 -92 7584 -90
rect 2007 -295 2009 -119
rect 2009 -295 2061 -119
rect 2061 -295 2063 -119
rect 6123 -295 6125 -119
rect 6125 -295 6177 -119
rect 6177 -295 6179 -119
<< metal3 >>
rect 1997 1063 2073 1068
rect 1997 887 2007 1063
rect 2063 887 2073 1063
rect 1997 882 2073 887
rect 6113 1063 6189 1068
rect 6113 887 6123 1063
rect 6179 887 6189 1063
rect 6113 882 6189 887
rect -244 860 1416 865
rect -244 804 606 860
rect 1406 804 1416 860
rect -244 799 1416 804
rect -244 -31 -178 799
rect 2005 674 2065 882
rect 6121 674 6181 882
rect 6774 860 8430 865
rect 6774 804 6784 860
rect 7584 804 8430 860
rect 6774 799 8430 804
rect 1997 669 2073 674
rect 1997 493 2007 669
rect 2063 493 2073 669
rect 1997 488 2073 493
rect 6113 669 6189 674
rect 6113 493 6123 669
rect 6179 493 6189 669
rect 6113 488 6189 493
rect 2005 280 2065 488
rect 6121 280 6181 488
rect 1997 275 2073 280
rect 1997 99 2007 275
rect 2063 99 2073 275
rect 1997 94 2073 99
rect 6113 275 6189 280
rect 6113 99 6123 275
rect 6179 99 6189 275
rect 6113 94 6189 99
rect -244 -36 1416 -31
rect -244 -92 606 -36
rect 1406 -92 1416 -36
rect -244 -97 1416 -92
rect 2005 -114 2065 94
rect 6121 -114 6181 94
rect 8364 -31 8430 799
rect 6774 -36 8430 -31
rect 6774 -92 6784 -36
rect 7584 -92 8430 -36
rect 6774 -97 8430 -92
rect 1997 -119 2073 -114
rect 1997 -295 2007 -119
rect 2063 -295 2073 -119
rect 1997 -300 2073 -295
rect 6113 -119 6189 -114
rect 6113 -295 6123 -119
rect 6179 -295 6189 -119
rect 6113 -300 6189 -295
use sky130_fd_pr__pfet_01v8_2XU96L  sky130_fd_pr__pfet_01v8_2XU96L_0
timestamp 1716189928
transform 1 0 -67 0 1 -207
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XU96L  sky130_fd_pr__pfet_01v8_2XU96L_1
timestamp 1716189928
transform 1 0 8253 0 1 975
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XU96L  sky130_fd_pr__pfet_01v8_2XU96L_2
timestamp 1716189928
transform 1 0 8253 0 1 581
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XU96L  sky130_fd_pr__pfet_01v8_2XU96L_3
timestamp 1716189928
transform 1 0 8253 0 1 187
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XU96L  sky130_fd_pr__pfet_01v8_2XU96L_4
timestamp 1716189928
transform 1 0 8253 0 1 -207
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XU96L  sky130_fd_pr__pfet_01v8_2XU96L_5
timestamp 1716189928
transform 1 0 -67 0 1 975
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XU96L  sky130_fd_pr__pfet_01v8_2XU96L_6
timestamp 1716189928
transform 1 0 -67 0 1 581
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XU96L  sky130_fd_pr__pfet_01v8_2XU96L_7
timestamp 1716189928
transform 1 0 -67 0 1 187
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_UKGYDC  sky130_fd_pr__pfet_01v8_UKGYDC_0
timestamp 1716128209
transform 1 0 4093 0 1 -207
box -4181 -162 4181 162
use sky130_fd_pr__pfet_01v8_UKGYDC  sky130_fd_pr__pfet_01v8_UKGYDC_1
timestamp 1716128209
transform 1 0 4093 0 1 975
box -4181 -162 4181 162
use sky130_fd_pr__pfet_01v8_UKGYDC  sky130_fd_pr__pfet_01v8_UKGYDC_2
timestamp 1716128209
transform 1 0 4093 0 1 581
box -4181 -162 4181 162
use sky130_fd_pr__pfet_01v8_UKGYDC  sky130_fd_pr__pfet_01v8_UKGYDC_3
timestamp 1716128209
transform 1 0 4093 0 1 187
box -4181 -162 4181 162
<< labels >>
flabel metal1 6136 1182 6160 1196 0 FreeSans 320 0 0 0 VDD
port 6 nsew
flabel metal2 8192 412 8228 434 0 FreeSans 320 0 0 0 net5
port 5 nsew
flabel metal1 8192 322 8228 342 0 FreeSans 320 0 0 0 net4
port 4 nsew
flabel metal1 8240 784 8268 798 0 FreeSans 320 0 0 0 net3
port 2 nsew
flabel metal2 4240 1128 4288 1152 0 FreeSans 320 0 0 0 net2
port 1 nsew
flabel metal3 7786 810 7840 844 0 FreeSans 320 0 0 0 net1
port 0 nsew
<< end >>
