magic
tech sky130A
magscale 1 2
timestamp 1717262354
<< nwell >>
rect -181 -67 8543 861
<< nsubdiff >>
rect -145 791 -85 825
rect 8447 791 8507 825
rect -145 765 -111 791
rect 8473 765 8507 791
rect -145 3 -111 29
rect 8473 3 8507 29
rect -145 -31 -85 3
rect 8447 -31 8507 3
<< nsubdiffcont >>
rect -85 791 8447 825
rect -145 29 -111 765
rect 8473 29 8507 765
rect -85 -31 8447 3
<< poly >>
rect 6 501 36 532
rect -56 485 36 501
rect -56 451 -40 485
rect -6 451 36 485
rect -56 435 36 451
rect 8326 501 8356 532
rect 8326 485 8418 501
rect 8326 451 8368 485
rect 8402 451 8418 485
rect 8326 435 8418 451
rect -56 343 36 359
rect -56 309 -40 343
rect -6 309 36 343
rect -56 293 36 309
rect 6 288 36 293
rect 8326 343 8418 359
rect 8326 309 8368 343
rect 8402 309 8418 343
rect 8326 293 8418 309
rect 8326 262 8356 293
<< polycont >>
rect -40 451 -6 485
rect 8368 451 8402 485
rect -40 309 -6 343
rect 8368 309 8402 343
<< locali >>
rect -145 791 -85 825
rect 8447 791 8507 825
rect -145 765 -111 791
rect 8473 765 8507 791
rect -40 485 -6 532
rect -40 435 -6 451
rect 8368 485 8402 532
rect 8368 435 8402 451
rect -40 343 -6 359
rect -40 257 -6 309
rect 8368 343 8402 359
rect 8368 262 8402 309
rect -145 3 -111 29
rect 8473 3 8507 29
rect -145 -31 -85 3
rect 8447 -31 8507 3
<< viali >>
rect 2106 791 2140 825
rect 6222 791 6256 825
rect -145 451 -111 485
rect -40 451 -6 485
rect 8368 451 8402 485
rect 8473 451 8507 485
rect -145 309 -111 343
rect -40 309 -6 343
rect 8368 309 8402 343
rect 8473 309 8507 343
rect 2106 -31 2140 3
rect 6222 -31 6256 3
<< metal1 >>
rect 2094 825 2152 831
rect 2094 791 2106 825
rect 2140 791 2152 825
rect 2094 720 2152 791
rect 6210 825 6268 831
rect 6210 791 6222 825
rect 6256 791 6268 825
rect 6210 720 6268 791
rect 29 544 39 720
rect 91 544 101 720
rect 2087 544 2097 720
rect 2149 544 2159 720
rect -46 497 0 532
rect -151 485 0 497
rect -151 451 -145 485
rect -111 451 -40 485
rect -6 451 0 485
rect -151 439 0 451
rect 590 420 1598 453
rect 2648 420 3656 451
rect 4158 420 4204 570
rect 6203 544 6213 720
rect 6265 544 6275 720
rect 8261 544 8271 720
rect 8323 544 8333 720
rect 8362 497 8408 532
rect 8362 485 8513 497
rect 4706 420 5714 453
rect 6764 420 7772 455
rect 8362 451 8368 485
rect 8402 451 8473 485
rect 8507 451 8513 485
rect 8362 439 8513 451
rect 42 374 8320 420
rect -151 343 0 355
rect -151 309 -145 343
rect -111 309 -40 343
rect -6 309 0 343
rect -151 297 0 309
rect -46 256 0 297
rect 42 252 88 374
rect 590 342 1598 374
rect 2648 340 3656 374
rect 4706 342 5714 374
rect 6764 344 7772 374
rect 2087 74 2097 250
rect 2149 74 2159 250
rect 4145 74 4155 250
rect 4207 74 4217 250
rect 6203 74 6213 250
rect 6265 74 6275 250
rect 8274 238 8320 374
rect 8362 343 8513 355
rect 8362 309 8368 343
rect 8402 309 8473 343
rect 8507 309 8513 343
rect 8362 297 8513 309
rect 8362 262 8408 297
rect 2094 3 2152 74
rect 2094 -31 2106 3
rect 2140 -31 2152 3
rect 2094 -37 2152 -31
rect 6210 3 6268 74
rect 6210 -31 6222 3
rect 6256 -31 6268 3
rect 6210 -37 6268 -31
<< via1 >>
rect 39 544 91 720
rect 2097 544 2149 720
rect 6213 544 6265 720
rect 8271 544 8323 720
rect 2097 74 2149 250
rect 4155 74 4207 250
rect 6213 74 6265 250
<< metal2 >>
rect 39 720 91 730
rect 39 423 91 544
rect 2095 720 2151 730
rect 2095 534 2151 544
rect 6211 720 6267 730
rect 6211 534 6267 544
rect 8271 720 8323 730
rect 8271 423 8323 544
rect 39 371 8323 423
rect 2095 250 2151 260
rect 2095 64 2151 74
rect 4155 250 4207 371
rect 4155 64 4207 74
rect 6211 250 6267 260
rect 6211 64 6267 74
<< via2 >>
rect 2095 544 2097 720
rect 2097 544 2149 720
rect 2149 544 2151 720
rect 6211 544 6213 720
rect 6213 544 6265 720
rect 6265 544 6267 720
rect 2095 74 2097 250
rect 2097 74 2149 250
rect 2149 74 2151 250
rect 6211 74 6213 250
rect 6213 74 6265 250
rect 6265 74 6267 250
<< metal3 >>
rect 2085 720 2161 725
rect 2085 544 2095 720
rect 2151 544 2161 720
rect 2085 539 2161 544
rect 6201 720 6277 725
rect 6201 544 6211 720
rect 6267 544 6277 720
rect 6201 539 6277 544
rect 2093 255 2153 539
rect 6209 255 6269 539
rect 2085 250 2161 255
rect 2085 74 2095 250
rect 2151 74 2161 250
rect 2085 69 2161 74
rect 6201 250 6277 255
rect 6201 74 6211 250
rect 6267 74 6277 250
rect 6201 69 6277 74
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_0
timestamp 1717262354
transform 1 0 8341 0 1 632
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_2
timestamp 1717262354
transform 1 0 8341 0 1 162
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_3
timestamp 1717262354
transform 1 0 21 0 1 632
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_4
timestamp 1717262354
transform 1 0 21 0 1 162
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_8WJSP2  sky130_fd_pr__pfet_01v8_8WJSP2_1
timestamp 1717262354
transform 1 0 4181 0 1 198
box -4181 -198 4181 164
use sky130_fd_pr__pfet_01v8_C2SSBD  sky130_fd_pr__pfet_01v8_C2SSBD_0
timestamp 1717262354
transform 1 0 4181 0 1 596
box -4181 -164 4181 198
<< labels >>
flabel metal2 8293 436 8293 436 0 FreeSans 160 0 0 0 D8
port 0 nsew
flabel metal1 8301 321 8301 321 0 FreeSans 160 0 0 0 D9
port 1 nsew
flabel metal1 6239 21 6239 21 0 FreeSans 160 0 0 0 VDD
port 2 nsew
<< end >>
