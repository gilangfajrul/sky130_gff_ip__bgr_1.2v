magic
tech sky130A
magscale 1 2
timestamp 1717511437
<< checkpaint >>
rect -883 -1766 1638 755
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
use sky130_fd_pr__res_high_po_0p35_KLM4B5  XR1
timestamp 0
transform 1 0 148 0 1 1776
box -201 -2282 201 2282
use sky130_fd_pr__res_high_po_0p35_YVVSCA  XR2
timestamp 0
transform 1 0 349 0 1 -506
box 0 0 1 1
use sky130_fd_pr__res_high_po_0p35_YVVSCA  XR3
timestamp 0
transform 1 0 350 0 1 -506
box 0 0 1 1
use sky130_fd_pr__res_high_po_0p35_YVVSCA  XR4
timestamp 0
transform 1 0 351 0 1 -506
box 0 0 1 1
use sky130_fd_pr__res_high_po_0p35_YVVSCA  XR5
timestamp 0
transform 1 0 352 0 1 -506
box 0 0 1 1
use sky130_fd_pr__res_high_po_0p35_YVVSCA  XR6
timestamp 0
transform 1 0 353 0 1 -506
box 0 0 1 1
use sky130_fd_pr__res_high_po_0p35_YVVSCA  XR7
timestamp 0
transform 1 0 354 0 1 -506
box 0 0 1 1
use sky130_fd_pr__res_high_po_0p35_YVVSCA  XR8
timestamp 0
transform 1 0 355 0 1 -506
box 0 0 1 1
use sky130_fd_pr__res_high_po_0p35_YVVSCA  XR9
timestamp 0
transform 1 0 356 0 1 -506
box 0 0 1 1
use sky130_fd_pr__res_high_po_0p35_YVVSCA  XR10
timestamp 0
transform 1 0 357 0 1 -506
box 0 0 1 1
use sky130_fd_pr__res_high_po_0p35_YVVSCA  XR11
timestamp 0
transform 1 0 358 0 1 -506
box 0 0 1 1
use sky130_fd_pr__res_high_po_0p35_YVVSCA  XR12
timestamp 0
transform 1 0 359 0 1 -506
box 0 0 1 1
use sky130_fd_pr__res_high_po_0p35_YVVSCA  XR13
timestamp 0
transform 1 0 360 0 1 -506
box 0 0 1 1
use sky130_fd_pr__res_high_po_0p35_YVVSCA  XR14
timestamp 0
transform 1 0 361 0 1 -506
box 0 0 1 1
use sky130_fd_pr__res_high_po_0p35_YVVSCA  XR15
timestamp 0
transform 1 0 362 0 1 -506
box 0 0 1 1
use sky130_fd_pr__res_high_po_0p35_YVVSCA  XR16
timestamp 0
transform 1 0 363 0 1 -506
box 0 0 1 1
use sky130_fd_pr__res_high_po_0p35_YVVSCA  XR17
timestamp 0
transform 1 0 364 0 1 -506
box 0 0 1 1
use sky130_fd_pr__res_high_po_0p35_YVVSCA  XR18
timestamp 0
transform 1 0 365 0 1 -506
box 0 0 1 1
use sky130_fd_pr__res_high_po_0p35_YVVSCA  XR19
timestamp 0
transform 1 0 366 0 1 -506
box 0 0 1 1
use sky130_fd_pr__res_high_po_0p35_YVVSCA  XR20
timestamp 0
transform 1 0 367 0 1 -506
box 0 0 1 1
use sky130_fd_pr__res_high_po_0p35_YVVSCA  XR21
timestamp 0
transform 1 0 368 0 1 -506
box 0 0 1 1
use sky130_fd_pr__res_high_po_0p35_YVVSCA  XR22
timestamp 0
transform 1 0 369 0 1 -506
box 0 0 1 1
use sky130_fd_pr__res_high_po_0p35_YVVSCA  XR23
timestamp 0
transform 1 0 370 0 1 -506
box 0 0 1 1
use sky130_fd_pr__res_high_po_0p35_YVVSCA  XR24
timestamp 0
transform 1 0 371 0 1 -506
box 0 0 1 1
use sky130_fd_pr__res_high_po_0p35_YVVSCA  XR25
timestamp 0
transform 1 0 372 0 1 -506
box 0 0 1 1
use sky130_fd_pr__res_high_po_0p35_YVVSCA  XR26
timestamp 0
transform 1 0 373 0 1 -506
box 0 0 1 1
use sky130_fd_pr__res_high_po_0p35_YVVSCA  XR27
timestamp 0
transform 1 0 374 0 1 -506
box 0 0 1 1
use sky130_fd_pr__res_high_po_0p35_YVVSCA  XR28
timestamp 0
transform 1 0 375 0 1 -506
box 0 0 1 1
use sky130_fd_pr__res_high_po_0p35_YVVSCA  XR29
timestamp 0
transform 1 0 376 0 1 -506
box 0 0 1 1
use sky130_fd_pr__res_high_po_0p35_YVVSCA  XR30
timestamp 0
transform 1 0 377 0 1 -506
box 0 0 1 1
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 B
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 A
port 1 nsew
<< end >>
