magic
tech sky130A
magscale 1 2
timestamp 1716351939
<< xpolycontact >>
rect -450 590 -380 1022
rect -450 52 -380 484
rect -284 590 -214 1022
rect -284 52 -214 484
rect -118 590 -48 1022
rect -118 52 -48 484
rect 48 590 118 1022
rect 48 52 118 484
rect 214 590 284 1022
rect 214 52 284 484
rect 380 590 450 1022
rect 380 52 450 484
rect -450 -484 -380 -52
rect -450 -1022 -380 -590
rect -284 -484 -214 -52
rect -284 -1022 -214 -590
rect -118 -484 -48 -52
rect -118 -1022 -48 -590
rect 48 -484 118 -52
rect 48 -1022 118 -590
rect 214 -484 284 -52
rect 214 -1022 284 -590
rect 380 -484 450 -52
rect 380 -1022 450 -590
<< ppolyres >>
rect -450 484 -380 590
rect -284 484 -214 590
rect -118 484 -48 590
rect 48 484 118 590
rect 214 484 284 590
rect 380 484 450 590
rect -450 -590 -380 -484
rect -284 -590 -214 -484
rect -118 -590 -48 -484
rect 48 -590 118 -484
rect 214 -590 284 -484
rect 380 -590 450 -484
<< viali >>
rect -434 607 -396 1004
rect -268 607 -230 1004
rect -102 607 -64 1004
rect 64 607 102 1004
rect 230 607 268 1004
rect 396 607 434 1004
rect -434 70 -396 467
rect -268 70 -230 467
rect -102 70 -64 467
rect 64 70 102 467
rect 230 70 268 467
rect 396 70 434 467
rect -434 -467 -396 -70
rect -268 -467 -230 -70
rect -102 -467 -64 -70
rect 64 -467 102 -70
rect 230 -467 268 -70
rect 396 -467 434 -70
rect -434 -1004 -396 -607
rect -268 -1004 -230 -607
rect -102 -1004 -64 -607
rect 64 -1004 102 -607
rect 230 -1004 268 -607
rect 396 -1004 434 -607
<< metal1 >>
rect -440 1004 -390 1016
rect -440 607 -434 1004
rect -396 607 -390 1004
rect -440 595 -390 607
rect -274 1004 -224 1016
rect -274 607 -268 1004
rect -230 607 -224 1004
rect -274 595 -224 607
rect -108 1004 -58 1016
rect -108 607 -102 1004
rect -64 607 -58 1004
rect -108 595 -58 607
rect 58 1004 108 1016
rect 58 607 64 1004
rect 102 607 108 1004
rect 58 595 108 607
rect 224 1004 274 1016
rect 224 607 230 1004
rect 268 607 274 1004
rect 224 595 274 607
rect 390 1004 440 1016
rect 390 607 396 1004
rect 434 607 440 1004
rect 390 595 440 607
rect -440 467 -390 479
rect -440 70 -434 467
rect -396 70 -390 467
rect -440 58 -390 70
rect -274 467 -224 479
rect -274 70 -268 467
rect -230 70 -224 467
rect -274 58 -224 70
rect -108 467 -58 479
rect -108 70 -102 467
rect -64 70 -58 467
rect -108 58 -58 70
rect 58 467 108 479
rect 58 70 64 467
rect 102 70 108 467
rect 58 58 108 70
rect 224 467 274 479
rect 224 70 230 467
rect 268 70 274 467
rect 224 58 274 70
rect 390 467 440 479
rect 390 70 396 467
rect 434 70 440 467
rect 390 58 440 70
rect -440 -70 -390 -58
rect -440 -467 -434 -70
rect -396 -467 -390 -70
rect -440 -479 -390 -467
rect -274 -70 -224 -58
rect -274 -467 -268 -70
rect -230 -467 -224 -70
rect -274 -479 -224 -467
rect -108 -70 -58 -58
rect -108 -467 -102 -70
rect -64 -467 -58 -70
rect -108 -479 -58 -467
rect 58 -70 108 -58
rect 58 -467 64 -70
rect 102 -467 108 -70
rect 58 -479 108 -467
rect 224 -70 274 -58
rect 224 -467 230 -70
rect 268 -467 274 -70
rect 224 -479 274 -467
rect 390 -70 440 -58
rect 390 -467 396 -70
rect 434 -467 440 -70
rect 390 -479 440 -467
rect -440 -607 -390 -595
rect -440 -1004 -434 -607
rect -396 -1004 -390 -607
rect -440 -1016 -390 -1004
rect -274 -607 -224 -595
rect -274 -1004 -268 -607
rect -230 -1004 -224 -607
rect -274 -1016 -224 -1004
rect -108 -607 -58 -595
rect -108 -1004 -102 -607
rect -64 -1004 -58 -607
rect -108 -1016 -58 -1004
rect 58 -607 108 -595
rect 58 -1004 64 -607
rect 102 -1004 108 -607
rect 58 -1016 108 -1004
rect 224 -607 274 -595
rect 224 -1004 230 -607
rect 268 -1004 274 -607
rect 224 -1016 274 -1004
rect 390 -607 440 -595
rect 390 -1004 396 -607
rect 434 -1004 440 -607
rect 390 -1016 440 -1004
<< properties >>
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.350 l 0.69 m 2 nx 6 wmin 0.350 lmin 0.50 rho 319.8 val 1.743k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
