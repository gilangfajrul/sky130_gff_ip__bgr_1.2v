magic
tech sky130A
magscale 1 2
timestamp 1720269525
<< psubdiff >>
rect 2269 -2147 2329 -2113
rect 28411 -2147 28471 -2113
rect 2269 -2173 2303 -2147
rect 2269 -3918 2303 -3892
rect 28437 -2173 28471 -2147
rect 28437 -3918 28471 -3892
rect 2269 -3952 2329 -3918
rect 28411 -3952 28471 -3918
<< psubdiffcont >>
rect 2329 -2147 28411 -2113
rect 2269 -3892 2303 -2173
rect 28437 -3892 28471 -2173
rect 2329 -3952 28411 -3918
<< viali >>
rect 2269 -2147 2329 -2113
rect 2329 -2147 28411 -2113
rect 28411 -2147 28471 -2113
rect 2269 -2173 2303 -2147
rect 2269 -3892 2303 -2173
rect 2269 -3918 2303 -3892
rect 28437 -2173 28471 -2147
rect 28437 -3892 28471 -2173
rect 28437 -3918 28471 -3892
rect 2269 -3952 2329 -3918
rect 2329 -3952 28411 -3918
rect 28411 -3952 28471 -3918
<< metal1 >>
rect 2263 -2107 2309 -2103
rect 28431 -2107 28477 -2103
rect 2257 -2113 28483 -2107
rect 2257 -2153 2269 -2113
rect 2263 -3912 2269 -2153
rect 2257 -3952 2269 -3912
rect 2303 -2153 28437 -2147
rect 2303 -2253 2309 -2153
rect 28431 -2253 28437 -2153
rect 2303 -2303 2452 -2253
rect 6628 -2303 6768 -2253
rect 10964 -2303 11104 -2253
rect 15300 -2303 15440 -2253
rect 19636 -2303 19776 -2253
rect 23972 -2303 24112 -2253
rect 28270 -2303 28437 -2253
rect 2303 -3747 2309 -2303
rect 6768 -2418 6820 -2408
rect 2432 -2469 2471 -2419
rect 6628 -2469 6723 -2419
rect 6576 -2584 6628 -2574
rect 2432 -2635 2461 -2585
rect 6673 -2585 6723 -2469
rect 6768 -2480 6820 -2470
rect 10912 -2418 10964 -2408
rect 15440 -2418 15492 -2408
rect 10912 -2480 10964 -2470
rect 11009 -2469 11104 -2419
rect 15300 -2469 15395 -2419
rect 11009 -2585 11059 -2469
rect 6673 -2635 6768 -2585
rect 10964 -2635 11059 -2585
rect 11104 -2584 11156 -2574
rect 6576 -2646 6628 -2636
rect 11104 -2646 11156 -2636
rect 15248 -2584 15300 -2574
rect 15345 -2585 15395 -2469
rect 15440 -2480 15492 -2470
rect 19584 -2418 19636 -2408
rect 24112 -2418 24164 -2408
rect 19584 -2480 19636 -2470
rect 19681 -2469 19776 -2419
rect 23972 -2469 24067 -2419
rect 19681 -2585 19731 -2469
rect 15345 -2635 15440 -2585
rect 19636 -2635 19731 -2585
rect 19776 -2584 19828 -2574
rect 15248 -2646 15300 -2636
rect 19776 -2646 19828 -2636
rect 23920 -2584 23972 -2574
rect 24017 -2585 24067 -2469
rect 24112 -2480 24164 -2470
rect 28256 -2418 28308 -2408
rect 28256 -2480 28308 -2470
rect 24017 -2635 24112 -2585
rect 28308 -2635 28403 -2585
rect 23920 -2646 23972 -2636
rect 6768 -2750 6820 -2740
rect 2337 -2801 2432 -2751
rect 6628 -2801 6723 -2751
rect 2337 -3249 2387 -2801
rect 6576 -2916 6628 -2906
rect 2420 -3133 2470 -2917
rect 6673 -2917 6723 -2801
rect 6768 -2812 6820 -2802
rect 10912 -2750 10964 -2740
rect 15440 -2750 15492 -2740
rect 10912 -2812 10964 -2802
rect 11009 -2801 11104 -2751
rect 15300 -2801 15395 -2751
rect 11009 -2917 11059 -2801
rect 15345 -2840 15395 -2801
rect 15440 -2812 15492 -2802
rect 19584 -2750 19636 -2740
rect 24112 -2750 24164 -2740
rect 19584 -2812 19636 -2802
rect 19681 -2801 19776 -2751
rect 23972 -2801 24067 -2751
rect 19681 -2840 19731 -2801
rect 15345 -2878 19731 -2840
rect 6673 -2967 6768 -2917
rect 10964 -2967 11059 -2917
rect 11104 -2916 11156 -2906
rect 6576 -2978 6628 -2968
rect 11104 -2978 11156 -2968
rect 15248 -2916 15300 -2906
rect 19776 -2916 19828 -2906
rect 15248 -2978 15300 -2968
rect 15428 -3006 15475 -2917
rect 19616 -2966 19638 -2918
rect 19776 -2978 19828 -2968
rect 23920 -2916 23972 -2906
rect 24017 -2917 24067 -2801
rect 24112 -2812 24164 -2802
rect 28256 -2750 28308 -2740
rect 28256 -2812 28308 -2802
rect 28353 -2917 28403 -2635
rect 24017 -2967 24112 -2917
rect 28308 -2967 28403 -2917
rect 23920 -2978 23972 -2968
rect 15265 -3053 15475 -3006
rect 6576 -3082 6628 -3072
rect 11104 -3082 11156 -3072
rect 6576 -3144 6628 -3134
rect 6673 -3133 6768 -3083
rect 10964 -3133 11059 -3083
rect 6673 -3249 6723 -3133
rect 2337 -3299 2432 -3249
rect 6628 -3299 6723 -3249
rect 6768 -3248 6820 -3238
rect 6768 -3310 6820 -3300
rect 10912 -3248 10964 -3238
rect 11009 -3249 11059 -3133
rect 15265 -3133 15312 -3053
rect 19776 -3082 19828 -3072
rect 15345 -3133 15440 -3083
rect 19636 -3133 19731 -3083
rect 11104 -3144 11156 -3134
rect 15345 -3161 15395 -3133
rect 19681 -3161 19731 -3133
rect 19776 -3144 19828 -3134
rect 23920 -3082 23972 -3072
rect 23920 -3144 23972 -3134
rect 24017 -3133 24112 -3083
rect 28308 -3133 28403 -3083
rect 15345 -3210 19731 -3161
rect 15345 -3249 15395 -3210
rect 11009 -3299 11104 -3249
rect 15300 -3299 15395 -3249
rect 15440 -3248 15492 -3238
rect 10912 -3310 10964 -3300
rect 15440 -3310 15492 -3300
rect 19584 -3248 19636 -3238
rect 19681 -3249 19731 -3210
rect 24017 -3249 24067 -3133
rect 19681 -3299 19776 -3249
rect 23972 -3299 24067 -3249
rect 24112 -3248 24164 -3238
rect 19584 -3310 19636 -3300
rect 24112 -3310 24164 -3300
rect 28256 -3248 28308 -3238
rect 28256 -3310 28308 -3300
rect 6576 -3414 6628 -3404
rect 2432 -3465 2463 -3415
rect 11104 -3414 11156 -3404
rect 6576 -3476 6628 -3466
rect 6673 -3465 6768 -3415
rect 10964 -3465 11059 -3415
rect 6673 -3581 6723 -3465
rect 2432 -3631 2457 -3581
rect 6628 -3631 6723 -3581
rect 6768 -3580 6820 -3570
rect 6768 -3642 6820 -3632
rect 10912 -3580 10964 -3570
rect 11009 -3581 11059 -3465
rect 11104 -3476 11156 -3466
rect 15248 -3414 15300 -3404
rect 19776 -3414 19828 -3404
rect 15248 -3476 15300 -3466
rect 15345 -3465 15440 -3415
rect 19636 -3465 19731 -3415
rect 15345 -3581 15395 -3465
rect 11009 -3631 11104 -3581
rect 15300 -3631 15395 -3581
rect 15440 -3580 15492 -3570
rect 10912 -3642 10964 -3632
rect 15440 -3642 15492 -3632
rect 19584 -3580 19636 -3570
rect 19681 -3581 19731 -3465
rect 19776 -3476 19828 -3466
rect 23920 -3414 23972 -3404
rect 28353 -3415 28403 -3133
rect 23920 -3476 23972 -3466
rect 24017 -3465 24112 -3415
rect 28308 -3465 28403 -3415
rect 24017 -3581 24067 -3465
rect 19681 -3631 19776 -3581
rect 23972 -3631 24067 -3581
rect 24112 -3580 24164 -3570
rect 19584 -3642 19636 -3632
rect 24112 -3642 24164 -3632
rect 28256 -3580 28308 -3570
rect 28256 -3642 28308 -3632
rect 28431 -3747 28437 -2303
rect 2303 -3797 2467 -3747
rect 6628 -3797 6768 -3747
rect 10964 -3797 11104 -3747
rect 15300 -3797 15440 -3747
rect 19636 -3797 19776 -3747
rect 23972 -3797 24112 -3747
rect 28279 -3797 28437 -3747
rect 2303 -3912 2309 -3797
rect 28431 -3912 28437 -3797
rect 2303 -3918 28437 -3912
rect 28471 -2153 28483 -2113
rect 28471 -3912 28477 -2153
rect 28471 -3952 28483 -3912
rect 2257 -3958 28483 -3952
rect 2263 -3964 2309 -3958
rect 28431 -3964 28477 -3958
<< via1 >>
rect 6576 -2636 6628 -2584
rect 6768 -2470 6820 -2418
rect 10912 -2470 10964 -2418
rect 11104 -2636 11156 -2584
rect 15248 -2636 15300 -2584
rect 15440 -2470 15492 -2418
rect 19584 -2470 19636 -2418
rect 19776 -2636 19828 -2584
rect 23920 -2636 23972 -2584
rect 24112 -2470 24164 -2418
rect 28256 -2470 28308 -2418
rect 6576 -2968 6628 -2916
rect 6768 -2802 6820 -2750
rect 10912 -2802 10964 -2750
rect 15440 -2802 15492 -2750
rect 19584 -2802 19636 -2750
rect 11104 -2968 11156 -2916
rect 15248 -2968 15300 -2916
rect 19776 -2968 19828 -2916
rect 23920 -2968 23972 -2916
rect 24112 -2802 24164 -2750
rect 28256 -2802 28308 -2750
rect 6576 -3134 6628 -3082
rect 6768 -3300 6820 -3248
rect 10912 -3300 10964 -3248
rect 11104 -3134 11156 -3082
rect 19776 -3134 19828 -3082
rect 23920 -3134 23972 -3082
rect 15440 -3300 15492 -3248
rect 19584 -3300 19636 -3248
rect 24112 -3300 24164 -3248
rect 28256 -3300 28308 -3248
rect 6576 -3466 6628 -3414
rect 6768 -3632 6820 -3580
rect 10912 -3632 10964 -3580
rect 11104 -3466 11156 -3414
rect 15248 -3466 15300 -3414
rect 15440 -3632 15492 -3580
rect 19584 -3632 19636 -3580
rect 19776 -3466 19828 -3414
rect 23920 -3466 23972 -3414
rect 24112 -3632 24164 -3580
rect 28256 -3632 28308 -3580
<< metal2 >>
rect 6672 -2470 6768 -2418
rect 6820 -2470 6830 -2418
rect 10902 -2470 10912 -2418
rect 10964 -2470 11060 -2418
rect 6672 -2584 6724 -2470
rect 6566 -2636 6576 -2584
rect 6628 -2636 6724 -2584
rect 11008 -2584 11060 -2470
rect 15344 -2470 15440 -2418
rect 15492 -2470 15502 -2418
rect 19574 -2470 19584 -2418
rect 19636 -2470 19732 -2418
rect 15344 -2584 15396 -2470
rect 11008 -2636 11104 -2584
rect 11156 -2636 11166 -2584
rect 15238 -2636 15248 -2584
rect 15300 -2636 15396 -2584
rect 19680 -2584 19732 -2470
rect 24016 -2470 24112 -2418
rect 24164 -2470 24174 -2418
rect 28246 -2470 28256 -2418
rect 28308 -2470 28404 -2418
rect 24016 -2584 24068 -2470
rect 19680 -2636 19776 -2584
rect 19828 -2636 19838 -2584
rect 23910 -2636 23920 -2584
rect 23972 -2636 24068 -2584
rect 28352 -2750 28404 -2470
rect 6672 -2802 6768 -2750
rect 6820 -2802 6830 -2750
rect 10902 -2802 10912 -2750
rect 10964 -2802 11060 -2750
rect 6672 -2916 6724 -2802
rect 6566 -2968 6576 -2916
rect 6628 -2968 6724 -2916
rect 11008 -2833 11060 -2802
rect 15344 -2802 15440 -2750
rect 15492 -2802 15502 -2750
rect 19574 -2802 19584 -2750
rect 19636 -2802 19732 -2750
rect 15344 -2833 15396 -2802
rect 11008 -2885 15396 -2833
rect 11008 -2916 11060 -2885
rect 15344 -2916 15396 -2885
rect 11008 -2968 11104 -2916
rect 11156 -2968 11166 -2916
rect 15238 -2968 15248 -2916
rect 15300 -2968 15396 -2916
rect 19680 -2916 19732 -2802
rect 24016 -2802 24112 -2750
rect 24164 -2802 24174 -2750
rect 28246 -2802 28256 -2750
rect 28308 -2802 28404 -2750
rect 24016 -2916 24068 -2802
rect 19680 -2968 19776 -2916
rect 19828 -2968 19838 -2916
rect 23910 -2968 23920 -2916
rect 23972 -2968 24068 -2916
rect 6566 -3134 6576 -3082
rect 6628 -3134 6724 -3082
rect 11094 -3134 11104 -3082
rect 11156 -3134 11166 -3082
rect 19680 -3134 19776 -3082
rect 19828 -3134 19838 -3082
rect 23910 -3134 23920 -3082
rect 23972 -3134 24068 -3082
rect 6672 -3248 6724 -3134
rect 11008 -3217 15396 -3165
rect 11008 -3248 11060 -3217
rect 6672 -3300 6768 -3248
rect 6820 -3300 6830 -3248
rect 10902 -3300 10912 -3248
rect 10964 -3300 11060 -3248
rect 15344 -3248 15396 -3217
rect 19680 -3248 19732 -3134
rect 15344 -3300 15440 -3248
rect 15492 -3300 15502 -3248
rect 19574 -3300 19584 -3248
rect 19636 -3300 19732 -3248
rect 24016 -3248 24068 -3134
rect 24016 -3300 24112 -3248
rect 24164 -3300 24174 -3248
rect 28246 -3300 28256 -3248
rect 28308 -3300 28404 -3248
rect 6566 -3466 6576 -3414
rect 6628 -3466 6724 -3414
rect 6672 -3580 6724 -3466
rect 11008 -3466 11104 -3414
rect 11156 -3466 11166 -3414
rect 15238 -3466 15248 -3414
rect 15300 -3466 15396 -3414
rect 11008 -3580 11060 -3466
rect 6672 -3632 6768 -3580
rect 6820 -3632 6830 -3580
rect 10902 -3632 10912 -3580
rect 10964 -3632 11060 -3580
rect 15344 -3580 15396 -3466
rect 19680 -3466 19776 -3414
rect 19828 -3466 19838 -3414
rect 23910 -3466 23920 -3414
rect 23972 -3466 24068 -3414
rect 19680 -3580 19732 -3466
rect 15344 -3632 15440 -3580
rect 15492 -3632 15502 -3580
rect 19574 -3632 19584 -3580
rect 19636 -3632 19732 -3580
rect 24016 -3580 24068 -3466
rect 28352 -3580 28404 -3300
rect 24016 -3632 24112 -3580
rect 24164 -3632 24174 -3580
rect 28246 -3632 28256 -3580
rect 28308 -3632 28404 -3580
use sky130_fd_pr__res_high_po_0p35_SU58NF  sky130_fd_pr__res_high_po_0p35_SU58NF_0
timestamp 1718867607
transform 0 -1 15370 1 0 -3025
box -782 -12956 782 12956
<< labels >>
flabel metal1 2435 -3628 2435 -3628 0 FreeSans 800 0 0 0 B
port 12 nsew
flabel metal1 2441 -3462 2441 -3462 0 FreeSans 800 0 0 0 D
port 11 nsew
flabel metal1 18977 -2863 18977 -2863 0 FreeSans 800 0 0 0 VBGSC
port 10 nsew
flabel metal1 24081 -2940 24081 -2940 0 FreeSans 800 0 0 0 VBGTC
port 8 nsew
flabel metal1 2442 -2632 2442 -2632 0 FreeSans 800 0 0 0 C
port 3 nsew
flabel metal1 2451 -2466 2451 -2466 0 FreeSans 800 0 0 0 A
port 2 nsew
flabel metal1 2281 -3956 2281 -3956 0 FreeSans 800 0 0 0 AVSS
port 15 nsew
flabel metal1 11111 -3080 11111 -3080 0 FreeSans 800 0 0 0 E
port 7 nsew
flabel metal1 19626 -2932 19626 -2932 0 FreeSans 1600 0 0 0 F
port 16 nsew
<< end >>
