magic
tech sky130A
magscale 1 2
timestamp 1716353109
<< psubdiff >>
rect -239 616 -179 650
rect 8343 616 8403 650
rect -239 590 -205 616
rect 8369 590 8403 616
rect -239 -141 -205 -115
rect 8369 -141 8403 -115
rect -239 -175 -179 -141
rect 8343 -175 8403 -141
<< psubdiffcont >>
rect -179 616 8343 650
rect -239 -115 -205 590
rect 8369 -115 8403 590
rect -179 -175 8343 -141
<< poly >>
rect -93 335 -63 354
rect -170 287 -63 335
rect 1282 328 1995 354
rect 2053 328 2766 354
rect 8227 335 8257 354
rect 1282 284 1908 328
rect 2140 284 2766 328
rect 3314 287 3966 328
rect 4198 287 4824 328
rect 5398 284 6024 328
rect 6256 284 6882 328
rect 8227 287 8334 335
rect -170 146 -63 194
rect 1282 167 1908 211
rect 2140 167 2766 211
rect 1282 145 1995 167
rect 2053 145 2766 167
rect 3314 147 3966 188
rect 4198 147 4824 188
rect 5398 147 6024 191
rect 6256 147 6882 191
rect 1282 141 1959 145
rect 2093 141 2766 145
rect 8227 140 8334 188
rect 8227 121 8257 140
<< locali >>
rect -239 616 -179 650
rect 8343 616 8403 650
rect -239 590 -205 616
rect 8369 590 8403 616
rect -139 328 -105 354
rect 2007 350 2041 354
rect 8269 328 8303 354
rect -139 119 -105 153
rect 8269 121 8303 147
rect -239 -141 -205 -115
rect 8369 -141 8403 -115
rect -239 -175 -179 -141
rect 8343 -175 8403 -141
<< viali >>
rect 1998 616 2050 650
rect 6114 616 6166 650
rect -239 294 -205 328
rect -157 294 -93 328
rect 1295 294 1895 328
rect 2153 294 2753 328
rect 3327 294 3953 328
rect 4211 294 4811 328
rect 5411 294 6011 328
rect 6269 294 6869 328
rect 8257 294 8321 328
rect 8369 294 8403 328
rect -239 153 -205 187
rect -157 153 -93 187
rect 1295 167 1895 201
rect 2153 167 2753 201
rect 3327 147 3953 181
rect 4211 147 4811 181
rect 5411 147 6011 181
rect 6269 147 6869 181
rect 8257 147 8321 181
rect 8369 147 8403 181
rect 1998 -175 2050 -141
rect 6114 -175 6166 -141
<< metal1 >>
rect 1988 656 1998 659
rect 1986 610 1998 656
rect 2050 656 2060 659
rect 6104 656 6114 659
rect 1988 607 1998 610
rect 2050 610 2062 656
rect 6102 610 6114 656
rect 6166 656 6176 659
rect 2050 607 2060 610
rect 6104 607 6114 610
rect 6166 610 6178 656
rect 6166 607 6176 610
rect -57 531 8221 579
rect -57 476 -11 531
rect 1988 366 1998 502
rect 2050 366 2060 502
rect 4059 461 4105 531
rect 6104 366 6114 502
rect 6166 366 6176 502
rect 8175 465 8221 531
rect -145 334 -99 354
rect -251 328 -81 334
rect -251 294 -239 328
rect -205 294 -157 328
rect -93 294 -81 328
rect -251 288 -81 294
rect 1283 285 1295 337
rect 1895 285 1907 337
rect -251 187 -81 193
rect -251 153 -239 187
rect -205 153 -157 187
rect -93 153 -81 187
rect 1283 158 1295 210
rect 1895 158 1907 210
rect -251 147 -81 153
rect -145 121 -99 147
rect 2001 111 2047 354
rect 2141 285 2153 337
rect 2753 285 2765 337
rect 3315 328 3965 334
rect 3315 294 3327 328
rect 3953 326 3965 328
rect 4199 328 4823 334
rect 4199 326 4211 328
rect 3953 294 4211 326
rect 4811 294 4823 328
rect 3315 286 4823 294
rect 5399 285 5411 337
rect 6011 285 6023 337
rect 2141 158 2153 210
rect 2753 158 2765 210
rect 3315 181 4823 189
rect 3315 147 3327 181
rect 3953 149 4211 181
rect 3953 147 3965 149
rect 3315 141 3965 147
rect 4199 147 4211 149
rect 4811 147 4823 181
rect 4199 141 4823 147
rect 5399 138 5411 190
rect 6011 138 6023 190
rect 6117 115 6163 366
rect 6257 285 6269 337
rect 6869 285 6881 337
rect 8263 334 8309 354
rect 8245 328 8415 334
rect 8245 294 8257 328
rect 8321 294 8369 328
rect 8403 294 8415 328
rect 8245 288 8415 294
rect 6257 138 6269 190
rect 6869 138 6881 190
rect 8245 181 8415 187
rect 8245 147 8257 181
rect 8321 147 8369 181
rect 8403 147 8415 181
rect 8245 141 8415 147
rect 8263 121 8309 141
rect -57 -56 -11 29
rect 4059 -56 4105 66
rect 6104 -7 6114 109
rect 6166 -7 6176 109
rect 8175 -56 8221 18
rect -57 -104 8221 -56
rect 1988 -135 1998 -132
rect 1986 -181 1998 -135
rect 2050 -135 2060 -132
rect 6104 -135 6114 -132
rect 1988 -184 1998 -181
rect 2050 -181 2062 -135
rect 6102 -181 6114 -135
rect 6166 -135 6176 -132
rect 2050 -184 2060 -181
rect 6104 -184 6114 -181
rect 6166 -181 6178 -135
rect 6166 -184 6176 -181
<< via1 >>
rect 1998 650 2050 659
rect 1998 616 2050 650
rect 1998 607 2050 616
rect 6114 650 6166 659
rect 6114 616 6166 650
rect 6114 607 6166 616
rect 1998 366 2050 502
rect 6114 366 6166 502
rect 1295 328 1895 337
rect 1295 294 1895 328
rect 1295 285 1895 294
rect 1295 201 1895 210
rect 1295 167 1895 201
rect 1295 158 1895 167
rect 2153 328 2753 337
rect 2153 294 2753 328
rect 2153 285 2753 294
rect 5411 328 6011 337
rect 5411 294 6011 328
rect 5411 285 6011 294
rect 2153 201 2753 210
rect 2153 167 2753 201
rect 2153 158 2753 167
rect 5411 181 6011 190
rect 5411 147 6011 181
rect 5411 138 6011 147
rect 6269 328 6869 337
rect 6269 294 6869 328
rect 6269 285 6869 294
rect 6269 181 6869 190
rect 6269 147 6869 181
rect 6269 138 6869 147
rect 6114 -7 6166 109
rect 1998 -141 2050 -132
rect 1998 -175 2050 -141
rect 1998 -184 2050 -175
rect 6114 -141 6166 -132
rect 6114 -175 6166 -141
rect 6114 -184 6166 -175
<< metal2 >>
rect 1998 659 2050 669
rect 1998 502 2050 607
rect 1998 356 2050 366
rect 6114 659 6166 669
rect 6114 502 6166 607
rect 6114 356 6166 366
rect 1295 339 1895 349
rect 2153 337 2753 347
rect 1295 273 1895 283
rect 2007 294 2153 328
rect 1295 210 1895 220
rect 2007 201 2041 294
rect 2153 275 2753 285
rect 5411 337 6011 347
rect 6269 339 6869 349
rect 6011 294 6157 328
rect 5411 275 6011 285
rect 1895 167 2041 201
rect 2153 212 2753 222
rect 1295 148 1895 158
rect 2153 146 2753 156
rect 5411 192 6011 202
rect 6123 181 6157 294
rect 6269 273 6869 283
rect 6269 190 6869 200
rect 6123 147 6269 181
rect 5411 126 6011 136
rect 6269 128 6869 138
rect 6114 109 6166 119
rect 1998 -132 2050 -54
rect 1998 -194 2050 -184
rect 6114 -132 6166 -7
rect 6114 -194 6166 -184
<< via2 >>
rect 1295 337 1895 339
rect 1295 285 1895 337
rect 1295 283 1895 285
rect 6269 337 6869 339
rect 2153 210 2753 212
rect 2153 158 2753 210
rect 2153 156 2753 158
rect 5411 190 6011 192
rect 5411 138 6011 190
rect 6269 285 6869 337
rect 6269 283 6869 285
rect 5411 136 6011 138
<< metal3 >>
rect 1285 342 1905 344
rect 6259 342 6879 344
rect 1285 339 2055 342
rect 1285 283 1295 339
rect 1895 283 2055 339
rect 1285 280 2055 283
rect 1285 278 1905 280
rect 1993 215 2055 280
rect 6109 339 6879 342
rect 6109 283 6269 339
rect 6869 283 6879 339
rect 6109 280 6879 283
rect 2143 215 2763 217
rect 1993 212 2763 215
rect 1993 156 2153 212
rect 2753 156 2763 212
rect 1993 153 2763 156
rect 2143 151 2763 153
rect 5401 195 6021 197
rect 6109 195 6171 280
rect 6259 278 6879 280
rect 5401 192 6171 195
rect 5401 136 5411 192
rect 6011 136 6171 192
rect 5401 133 6171 136
rect 5401 131 6021 133
use sky130_fd_pr__nfet_01v8_EDB9KC  sky130_fd_pr__nfet_01v8_EDB9KC_0
timestamp 1716303658
transform 1 0 148 0 1 207
box 0 0 1 1
use sky130_fd_pr__nfet_01v8_S9SDYN  sky130_fd_pr__nfet_01v8_S9SDYN_0
timestamp 1716353109
transform 1 0 -78 0 1 51
box -73 -96 73 96
use sky130_fd_pr__nfet_01v8_S9SDYN  sky130_fd_pr__nfet_01v8_S9SDYN_1
timestamp 1716353109
transform 1 0 -78 0 1 424
box -73 -96 73 96
use sky130_fd_pr__nfet_01v8_S9SDYN  sky130_fd_pr__nfet_01v8_S9SDYN_2
timestamp 1716353109
transform 1 0 8242 0 1 424
box -73 -96 73 96
use sky130_fd_pr__nfet_01v8_S9SDYN  sky130_fd_pr__nfet_01v8_S9SDYN_3
timestamp 1716353109
transform 1 0 8242 0 1 51
box -73 -96 73 96
use sky130_fd_pr__nfet_01v8_X6WGLW  sky130_fd_pr__nfet_01v8_X6WGLW_0
timestamp 1716353109
transform -1 0 4082 0 1 51
box -4145 -96 4145 96
use sky130_fd_pr__nfet_01v8_X6WGLW  sky130_fd_pr__nfet_01v8_X6WGLW_1
timestamp 1716353109
transform -1 0 4082 0 1 424
box -4145 -96 4145 96
<< end >>
