magic
tech sky130A
magscale 1 2
timestamp 1717267244
<< nwell >>
rect -677 -3195 677 3195
<< nsubdiff >>
rect -641 3125 -545 3159
rect 545 3125 641 3159
rect -641 3063 -607 3125
rect 607 3063 641 3125
rect -641 -3125 -607 -3063
rect 607 -3125 641 -3063
rect -641 -3159 -545 -3125
rect 545 -3159 641 -3125
<< nsubdiffcont >>
rect -545 3125 545 3159
rect -641 -3063 -607 3063
rect 607 -3063 641 3063
rect -545 -3159 545 -3125
<< xpolycontact >>
rect -450 2588 -380 3020
rect -450 1588 -380 2020
rect -284 2588 -214 3020
rect -284 1588 -214 2020
rect -118 2588 -48 3020
rect -118 1588 -48 2020
rect 48 2588 118 3020
rect 48 1588 118 2020
rect 214 2588 284 3020
rect 214 1588 284 2020
rect 380 2588 450 3020
rect 380 1588 450 2020
rect -450 1052 -380 1484
rect -450 52 -380 484
rect -284 1052 -214 1484
rect -284 52 -214 484
rect -118 1052 -48 1484
rect -118 52 -48 484
rect 48 1052 118 1484
rect 48 52 118 484
rect 214 1052 284 1484
rect 214 52 284 484
rect 380 1052 450 1484
rect 380 52 450 484
rect -450 -484 -380 -52
rect -450 -1484 -380 -1052
rect -284 -484 -214 -52
rect -284 -1484 -214 -1052
rect -118 -484 -48 -52
rect -118 -1484 -48 -1052
rect 48 -484 118 -52
rect 48 -1484 118 -1052
rect 214 -484 284 -52
rect 214 -1484 284 -1052
rect 380 -484 450 -52
rect 380 -1484 450 -1052
rect -450 -2020 -380 -1588
rect -450 -3020 -380 -2588
rect -284 -2020 -214 -1588
rect -284 -3020 -214 -2588
rect -118 -2020 -48 -1588
rect -118 -3020 -48 -2588
rect 48 -2020 118 -1588
rect 48 -3020 118 -2588
rect 214 -2020 284 -1588
rect 214 -3020 284 -2588
rect 380 -2020 450 -1588
rect 380 -3020 450 -2588
<< ppolyres >>
rect -450 2020 -380 2588
rect -284 2020 -214 2588
rect -118 2020 -48 2588
rect 48 2020 118 2588
rect 214 2020 284 2588
rect 380 2020 450 2588
rect -450 484 -380 1052
rect -284 484 -214 1052
rect -118 484 -48 1052
rect 48 484 118 1052
rect 214 484 284 1052
rect 380 484 450 1052
rect -450 -1052 -380 -484
rect -284 -1052 -214 -484
rect -118 -1052 -48 -484
rect 48 -1052 118 -484
rect 214 -1052 284 -484
rect 380 -1052 450 -484
rect -450 -2588 -380 -2020
rect -284 -2588 -214 -2020
rect -118 -2588 -48 -2020
rect 48 -2588 118 -2020
rect 214 -2588 284 -2020
rect 380 -2588 450 -2020
<< locali >>
rect -641 3125 -545 3159
rect 545 3125 641 3159
rect -641 3063 -607 3125
rect 607 3063 641 3125
rect -641 -3125 -607 -3063
rect 607 -3125 641 -3063
rect -641 -3159 -545 -3125
rect 545 -3159 641 -3125
<< viali >>
rect -434 2605 -396 3002
rect -268 2605 -230 3002
rect -102 2605 -64 3002
rect 64 2605 102 3002
rect 230 2605 268 3002
rect 396 2605 434 3002
rect -434 1606 -396 2003
rect -268 1606 -230 2003
rect -102 1606 -64 2003
rect 64 1606 102 2003
rect 230 1606 268 2003
rect 396 1606 434 2003
rect -434 1069 -396 1466
rect -268 1069 -230 1466
rect -102 1069 -64 1466
rect 64 1069 102 1466
rect 230 1069 268 1466
rect 396 1069 434 1466
rect -434 70 -396 467
rect -268 70 -230 467
rect -102 70 -64 467
rect 64 70 102 467
rect 230 70 268 467
rect 396 70 434 467
rect -434 -467 -396 -70
rect -268 -467 -230 -70
rect -102 -467 -64 -70
rect 64 -467 102 -70
rect 230 -467 268 -70
rect 396 -467 434 -70
rect -434 -1466 -396 -1069
rect -268 -1466 -230 -1069
rect -102 -1466 -64 -1069
rect 64 -1466 102 -1069
rect 230 -1466 268 -1069
rect 396 -1466 434 -1069
rect -434 -2003 -396 -1606
rect -268 -2003 -230 -1606
rect -102 -2003 -64 -1606
rect 64 -2003 102 -1606
rect 230 -2003 268 -1606
rect 396 -2003 434 -1606
rect -434 -3002 -396 -2605
rect -268 -3002 -230 -2605
rect -102 -3002 -64 -2605
rect 64 -3002 102 -2605
rect 230 -3002 268 -2605
rect 396 -3002 434 -2605
<< metal1 >>
rect -440 3002 -390 3014
rect -440 2605 -434 3002
rect -396 2605 -390 3002
rect -440 2593 -390 2605
rect -274 3002 -224 3014
rect -274 2605 -268 3002
rect -230 2605 -224 3002
rect -274 2593 -224 2605
rect -108 3002 -58 3014
rect -108 2605 -102 3002
rect -64 2605 -58 3002
rect -108 2593 -58 2605
rect 58 3002 108 3014
rect 58 2605 64 3002
rect 102 2605 108 3002
rect 58 2593 108 2605
rect 224 3002 274 3014
rect 224 2605 230 3002
rect 268 2605 274 3002
rect 224 2593 274 2605
rect 390 3002 440 3014
rect 390 2605 396 3002
rect 434 2605 440 3002
rect 390 2593 440 2605
rect -440 2003 -390 2015
rect -440 1606 -434 2003
rect -396 1606 -390 2003
rect -440 1594 -390 1606
rect -274 2003 -224 2015
rect -274 1606 -268 2003
rect -230 1606 -224 2003
rect -274 1594 -224 1606
rect -108 2003 -58 2015
rect -108 1606 -102 2003
rect -64 1606 -58 2003
rect -108 1594 -58 1606
rect 58 2003 108 2015
rect 58 1606 64 2003
rect 102 1606 108 2003
rect 58 1594 108 1606
rect 224 2003 274 2015
rect 224 1606 230 2003
rect 268 1606 274 2003
rect 224 1594 274 1606
rect 390 2003 440 2015
rect 390 1606 396 2003
rect 434 1606 440 2003
rect 390 1594 440 1606
rect -440 1466 -390 1478
rect -440 1069 -434 1466
rect -396 1069 -390 1466
rect -440 1057 -390 1069
rect -274 1466 -224 1478
rect -274 1069 -268 1466
rect -230 1069 -224 1466
rect -274 1057 -224 1069
rect -108 1466 -58 1478
rect -108 1069 -102 1466
rect -64 1069 -58 1466
rect -108 1057 -58 1069
rect 58 1466 108 1478
rect 58 1069 64 1466
rect 102 1069 108 1466
rect 58 1057 108 1069
rect 224 1466 274 1478
rect 224 1069 230 1466
rect 268 1069 274 1466
rect 224 1057 274 1069
rect 390 1466 440 1478
rect 390 1069 396 1466
rect 434 1069 440 1466
rect 390 1057 440 1069
rect -440 467 -390 479
rect -440 70 -434 467
rect -396 70 -390 467
rect -440 58 -390 70
rect -274 467 -224 479
rect -274 70 -268 467
rect -230 70 -224 467
rect -274 58 -224 70
rect -108 467 -58 479
rect -108 70 -102 467
rect -64 70 -58 467
rect -108 58 -58 70
rect 58 467 108 479
rect 58 70 64 467
rect 102 70 108 467
rect 58 58 108 70
rect 224 467 274 479
rect 224 70 230 467
rect 268 70 274 467
rect 224 58 274 70
rect 390 467 440 479
rect 390 70 396 467
rect 434 70 440 467
rect 390 58 440 70
rect -440 -70 -390 -58
rect -440 -467 -434 -70
rect -396 -467 -390 -70
rect -440 -479 -390 -467
rect -274 -70 -224 -58
rect -274 -467 -268 -70
rect -230 -467 -224 -70
rect -274 -479 -224 -467
rect -108 -70 -58 -58
rect -108 -467 -102 -70
rect -64 -467 -58 -70
rect -108 -479 -58 -467
rect 58 -70 108 -58
rect 58 -467 64 -70
rect 102 -467 108 -70
rect 58 -479 108 -467
rect 224 -70 274 -58
rect 224 -467 230 -70
rect 268 -467 274 -70
rect 224 -479 274 -467
rect 390 -70 440 -58
rect 390 -467 396 -70
rect 434 -467 440 -70
rect 390 -479 440 -467
rect -440 -1069 -390 -1057
rect -440 -1466 -434 -1069
rect -396 -1466 -390 -1069
rect -440 -1478 -390 -1466
rect -274 -1069 -224 -1057
rect -274 -1466 -268 -1069
rect -230 -1466 -224 -1069
rect -274 -1478 -224 -1466
rect -108 -1069 -58 -1057
rect -108 -1466 -102 -1069
rect -64 -1466 -58 -1069
rect -108 -1478 -58 -1466
rect 58 -1069 108 -1057
rect 58 -1466 64 -1069
rect 102 -1466 108 -1069
rect 58 -1478 108 -1466
rect 224 -1069 274 -1057
rect 224 -1466 230 -1069
rect 268 -1466 274 -1069
rect 224 -1478 274 -1466
rect 390 -1069 440 -1057
rect 390 -1466 396 -1069
rect 434 -1466 440 -1069
rect 390 -1478 440 -1466
rect -440 -1606 -390 -1594
rect -440 -2003 -434 -1606
rect -396 -2003 -390 -1606
rect -440 -2015 -390 -2003
rect -274 -1606 -224 -1594
rect -274 -2003 -268 -1606
rect -230 -2003 -224 -1606
rect -274 -2015 -224 -2003
rect -108 -1606 -58 -1594
rect -108 -2003 -102 -1606
rect -64 -2003 -58 -1606
rect -108 -2015 -58 -2003
rect 58 -1606 108 -1594
rect 58 -2003 64 -1606
rect 102 -2003 108 -1606
rect 58 -2015 108 -2003
rect 224 -1606 274 -1594
rect 224 -2003 230 -1606
rect 268 -2003 274 -1606
rect 224 -2015 274 -2003
rect 390 -1606 440 -1594
rect 390 -2003 396 -1606
rect 434 -2003 440 -1606
rect 390 -2015 440 -2003
rect -440 -2605 -390 -2593
rect -440 -3002 -434 -2605
rect -396 -3002 -390 -2605
rect -440 -3014 -390 -3002
rect -274 -2605 -224 -2593
rect -274 -3002 -268 -2605
rect -230 -3002 -224 -2605
rect -274 -3014 -224 -3002
rect -108 -2605 -58 -2593
rect -108 -3002 -102 -2605
rect -64 -3002 -58 -2605
rect -108 -3014 -58 -3002
rect 58 -2605 108 -2593
rect 58 -3002 64 -2605
rect 102 -3002 108 -2605
rect 58 -3014 108 -3002
rect 224 -2605 274 -2593
rect 224 -3002 230 -2605
rect 268 -3002 274 -2605
rect 224 -3014 274 -3002
rect 390 -2605 440 -2593
rect 390 -3002 396 -2605
rect 434 -3002 440 -2605
rect 390 -3014 440 -3002
<< properties >>
string FIXED_BBOX -624 -3142 624 3142
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.350 l 3 m 4 nx 6 wmin 0.350 lmin 0.50 rho 319.8 val 3.854k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.350 vias 1 n_guard 1 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
