magic
tech sky130A
magscale 1 2
timestamp 1720109855
<< nwell >>
rect -176 -521 1222 851
<< nsubdiff >>
rect -140 781 -80 815
rect 1126 781 1186 815
rect -140 755 -106 781
rect 1152 755 1186 781
rect -140 -451 -106 -425
rect 1152 -451 1186 -425
rect -140 -485 -80 -451
rect 1126 -485 1186 -451
<< nsubdiffcont >>
rect -80 781 1126 815
rect -140 -425 -106 755
rect 1152 -425 1186 755
rect -80 -485 1126 -451
<< poly >>
rect 6 198 36 236
rect -50 182 36 198
rect -50 148 -40 182
rect -6 148 36 182
rect -50 132 36 148
rect 6 94 36 132
rect 94 94 952 236
rect 1010 198 1040 236
rect 1010 182 1096 198
rect 1010 148 1052 182
rect 1086 148 1096 182
rect 1010 132 1096 148
rect 1010 94 1040 132
<< polycont >>
rect -40 148 -6 182
rect 1052 148 1086 182
<< locali >>
rect -140 781 -80 815
rect 1126 781 1186 815
rect -140 755 -106 781
rect 1152 755 1186 781
rect -40 182 -6 198
rect -40 132 -6 148
rect 1052 182 1086 198
rect 1052 132 1086 148
rect -140 -451 -106 -425
rect 1152 -451 1186 -425
rect -140 -485 -80 -451
rect 1126 -485 1186 -451
<< viali >>
rect -40 148 -6 182
rect 1052 148 1086 182
<< metal1 >>
rect 389 703 660 748
rect 824 703 856 748
rect 487 274 497 650
rect 549 274 559 650
rect -46 188 0 263
rect 42 188 88 269
rect 958 188 1004 267
rect 1046 188 1092 265
rect -46 182 1092 188
rect -46 148 -40 182
rect -6 148 1052 182
rect 1086 148 1092 182
rect -46 142 1092 148
rect -46 67 0 142
rect 42 63 88 142
rect 958 61 1004 142
rect 1046 65 1092 142
rect 487 -320 497 56
rect 549 -320 559 56
rect 390 -419 661 -373
<< via1 >>
rect 497 274 549 650
rect 497 -320 549 56
<< metal2 >>
rect 497 650 549 660
rect 497 56 549 274
rect 497 -330 549 -320
use sky130_fd_pr__pfet_01v8_2ZH9EN  sky130_fd_pr__pfet_01v8_2ZH9EN_0
timestamp 1720109454
transform 1 0 21 0 1 -132
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9EN  sky130_fd_pr__pfet_01v8_2ZH9EN_1
timestamp 1720109454
transform 1 0 1025 0 1 -132
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9EN  sky130_fd_pr__pfet_01v8_2ZH9EN_2
timestamp 1720109454
transform 1 0 1025 0 1 462
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9EN  sky130_fd_pr__pfet_01v8_2ZH9EN_3
timestamp 1720109454
transform 1 0 21 0 1 462
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_9XC4R9  sky130_fd_pr__pfet_01v8_9XC4R9_0
timestamp 1720109454
transform 1 0 523 0 1 498
box -523 -298 523 264
use sky130_fd_pr__pfet_01v8_CVH45E  sky130_fd_pr__pfet_01v8_CVH45E_0
timestamp 1720109454
transform 1 0 523 0 1 -168
box -523 -264 523 298
<< labels >>
flabel metal1 982 156 982 156 0 FreeSans 160 0 0 0 VDDE
port 2 nsew
flabel metal2 528 257 528 257 0 FreeSans 160 0 0 0 AVDD
port 3 nsew
flabel metal1 848 730 848 730 0 FreeSans 160 0 0 0 G
port 0 nsew
flabel nsubdiffcont 1158 687 1158 687 0 FreeSans 160 0 0 0 DVDD
port 4 nsew
<< end >>
