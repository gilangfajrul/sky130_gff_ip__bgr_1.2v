magic
tech sky130A
magscale 1 2
timestamp 1717312722
<< metal3 >>
rect -4288 -2028 -3898 -1932
rect -6354 -4018 -6258 -3628
rect -2321 -4065 -2225 -3675
rect -4369 -5748 -3902 -5652
<< metal4 >>
rect -8858 1692 3764 1788
rect -6 1690 3764 1692
rect -10344 -7792 -10248 1395
rect -8365 -8015 -8267 618
rect -6354 -3792 -6258 -3603
rect -2321 -3792 -2225 -3535
rect -6354 -3888 -2225 -3792
rect -6354 -4132 -6258 -3888
rect -2321 -4064 -2225 -3888
rect 1691 -7826 1787 1361
rect 3670 -7828 3768 805
rect -8739 -9372 448 -9371
rect -8739 -9467 3764 -9372
rect -348 -9470 3764 -9467
use sky130_fd_pr__cap_mim_m3_1_SXWHWZ  sky130_fd_pr__cap_mim_m3_1_SXWHWZ_0
timestamp 1716453347
transform 1 0 -4133 0 1 -3840
box -7904 -7320 7904 7320
<< labels >>
flabel metal4 -3508 -3840 -3508 -3840 0 FreeSans 1600 0 0 0 A
port 0 nsew
flabel metal3 -4163 -1986 -4163 -1986 0 FreeSans 1600 0 0 0 B
port 1 nsew
flabel metal4 1735 -7571 1735 -7571 0 FreeSans 1600 0 0 0 GND
port 5 nsew
<< end >>
