magic
tech sky130A
magscale 1 2
timestamp 1762707440
<< nwell >>
rect -4181 -364 4181 364
<< pmos >>
rect -4087 64 -2087 264
rect -2029 64 -29 264
rect 29 64 2029 264
rect 2087 64 4087 264
rect -4087 -264 -2087 -64
rect -2029 -264 -29 -64
rect 29 -264 2029 -64
rect 2087 -264 4087 -64
<< pdiff >>
rect -4145 252 -4087 264
rect -4145 76 -4133 252
rect -4099 76 -4087 252
rect -4145 64 -4087 76
rect -2087 252 -2029 264
rect -2087 76 -2075 252
rect -2041 76 -2029 252
rect -2087 64 -2029 76
rect -29 252 29 264
rect -29 76 -17 252
rect 17 76 29 252
rect -29 64 29 76
rect 2029 252 2087 264
rect 2029 76 2041 252
rect 2075 76 2087 252
rect 2029 64 2087 76
rect 4087 252 4145 264
rect 4087 76 4099 252
rect 4133 76 4145 252
rect 4087 64 4145 76
rect -4145 -76 -4087 -64
rect -4145 -252 -4133 -76
rect -4099 -252 -4087 -76
rect -4145 -264 -4087 -252
rect -2087 -76 -2029 -64
rect -2087 -252 -2075 -76
rect -2041 -252 -2029 -76
rect -2087 -264 -2029 -252
rect -29 -76 29 -64
rect -29 -252 -17 -76
rect 17 -252 29 -76
rect -29 -264 29 -252
rect 2029 -76 2087 -64
rect 2029 -252 2041 -76
rect 2075 -252 2087 -76
rect 2029 -264 2087 -252
rect 4087 -76 4145 -64
rect 4087 -252 4099 -76
rect 4133 -252 4145 -76
rect 4087 -264 4145 -252
<< pdiffc >>
rect -4133 76 -4099 252
rect -2075 76 -2041 252
rect -17 76 17 252
rect 2041 76 2075 252
rect 4099 76 4133 252
rect -4133 -252 -4099 -76
rect -2075 -252 -2041 -76
rect -17 -252 17 -76
rect 2041 -252 2075 -76
rect 4099 -252 4133 -76
<< poly >>
rect -4087 345 -2087 361
rect -4087 311 -4071 345
rect -2103 311 -2087 345
rect -4087 264 -2087 311
rect -2029 345 -29 361
rect -2029 311 -2013 345
rect -45 311 -29 345
rect -2029 264 -29 311
rect 29 345 2029 361
rect 29 311 45 345
rect 2013 311 2029 345
rect 29 264 2029 311
rect 2087 345 4087 361
rect 2087 311 2103 345
rect 4071 311 4087 345
rect 2087 264 4087 311
rect -4087 17 -2087 64
rect -4087 -17 -4071 17
rect -2103 -17 -2087 17
rect -4087 -64 -2087 -17
rect -2029 17 -29 64
rect -2029 -17 -2013 17
rect -45 -17 -29 17
rect -2029 -64 -29 -17
rect 29 17 2029 64
rect 29 -17 45 17
rect 2013 -17 2029 17
rect 29 -64 2029 -17
rect 2087 17 4087 64
rect 2087 -17 2103 17
rect 4071 -17 4087 17
rect 2087 -64 4087 -17
rect -4087 -311 -2087 -264
rect -4087 -345 -4071 -311
rect -2103 -345 -2087 -311
rect -4087 -361 -2087 -345
rect -2029 -311 -29 -264
rect -2029 -345 -2013 -311
rect -45 -345 -29 -311
rect -2029 -361 -29 -345
rect 29 -311 2029 -264
rect 29 -345 45 -311
rect 2013 -345 2029 -311
rect 29 -361 2029 -345
rect 2087 -311 4087 -264
rect 2087 -345 2103 -311
rect 4071 -345 4087 -311
rect 2087 -361 4087 -345
<< polycont >>
rect -4071 311 -2103 345
rect -2013 311 -45 345
rect 45 311 2013 345
rect 2103 311 4071 345
rect -4071 -17 -2103 17
rect -2013 -17 -45 17
rect 45 -17 2013 17
rect 2103 -17 4071 17
rect -4071 -345 -2103 -311
rect -2013 -345 -45 -311
rect 45 -345 2013 -311
rect 2103 -345 4071 -311
<< locali >>
rect -4087 311 -4071 345
rect -2103 311 -2087 345
rect -2029 311 -2013 345
rect -45 311 -29 345
rect 29 311 45 345
rect 2013 311 2029 345
rect 2087 311 2103 345
rect 4071 311 4087 345
rect -4133 252 -4099 268
rect -4133 60 -4099 76
rect -2075 252 -2041 268
rect -2075 60 -2041 76
rect -17 252 17 268
rect -17 60 17 76
rect 2041 252 2075 268
rect 2041 60 2075 76
rect 4099 252 4133 268
rect 4099 60 4133 76
rect -4087 -17 -4071 17
rect -2103 -17 -2087 17
rect -2029 -17 -2013 17
rect -45 -17 -29 17
rect 29 -17 45 17
rect 2013 -17 2029 17
rect 2087 -17 2103 17
rect 4071 -17 4087 17
rect -4133 -76 -4099 -60
rect -4133 -268 -4099 -252
rect -2075 -76 -2041 -60
rect -2075 -268 -2041 -252
rect -17 -76 17 -60
rect -17 -268 17 -252
rect 2041 -76 2075 -60
rect 2041 -268 2075 -252
rect 4099 -76 4133 -60
rect 4099 -268 4133 -252
rect -4087 -345 -4071 -311
rect -2103 -345 -2087 -311
rect -2029 -345 -2013 -311
rect -45 -345 -29 -311
rect 29 -345 45 -311
rect 2013 -345 2029 -311
rect 2087 -345 2103 -311
rect 4071 -345 4087 -311
<< viali >>
rect -4071 311 -2103 345
rect -2013 311 -45 345
rect 45 311 2013 345
rect 2103 311 4071 345
rect -4133 76 -4099 252
rect -2075 76 -2041 252
rect -17 76 17 252
rect 2041 76 2075 252
rect 4099 76 4133 252
rect -4071 -17 -2103 17
rect -2013 -17 -45 17
rect 45 -17 2013 17
rect 2103 -17 4071 17
rect -4133 -252 -4099 -76
rect -2075 -252 -2041 -76
rect -17 -252 17 -76
rect 2041 -252 2075 -76
rect 4099 -252 4133 -76
rect -4071 -345 -2103 -311
rect -2013 -345 -45 -311
rect 45 -345 2013 -311
rect 2103 -345 4071 -311
<< metal1 >>
rect -4083 345 -2091 351
rect -4083 311 -4071 345
rect -2103 311 -2091 345
rect -4083 305 -2091 311
rect -2025 345 -33 351
rect -2025 311 -2013 345
rect -45 311 -33 345
rect -2025 305 -33 311
rect 33 345 2025 351
rect 33 311 45 345
rect 2013 311 2025 345
rect 33 305 2025 311
rect 2091 345 4083 351
rect 2091 311 2103 345
rect 4071 311 4083 345
rect 2091 305 4083 311
rect -4139 252 -4093 264
rect -4139 76 -4133 252
rect -4099 76 -4093 252
rect -4139 64 -4093 76
rect -2081 252 -2035 264
rect -2081 76 -2075 252
rect -2041 76 -2035 252
rect -2081 64 -2035 76
rect -23 252 23 264
rect -23 76 -17 252
rect 17 76 23 252
rect -23 64 23 76
rect 2035 252 2081 264
rect 2035 76 2041 252
rect 2075 76 2081 252
rect 2035 64 2081 76
rect 4093 252 4139 264
rect 4093 76 4099 252
rect 4133 76 4139 252
rect 4093 64 4139 76
rect -4083 17 -2091 23
rect -4083 -17 -4071 17
rect -2103 -17 -2091 17
rect -4083 -23 -2091 -17
rect -2025 17 -33 23
rect -2025 -17 -2013 17
rect -45 -17 -33 17
rect -2025 -23 -33 -17
rect 33 17 2025 23
rect 33 -17 45 17
rect 2013 -17 2025 17
rect 33 -23 2025 -17
rect 2091 17 4083 23
rect 2091 -17 2103 17
rect 4071 -17 4083 17
rect 2091 -23 4083 -17
rect -4139 -76 -4093 -64
rect -4139 -252 -4133 -76
rect -4099 -252 -4093 -76
rect -4139 -264 -4093 -252
rect -2081 -76 -2035 -64
rect -2081 -252 -2075 -76
rect -2041 -252 -2035 -76
rect -2081 -264 -2035 -252
rect -23 -76 23 -64
rect -23 -252 -17 -76
rect 17 -252 23 -76
rect -23 -264 23 -252
rect 2035 -76 2081 -64
rect 2035 -252 2041 -76
rect 2075 -252 2081 -76
rect 2035 -264 2081 -252
rect 4093 -76 4139 -64
rect 4093 -252 4099 -76
rect 4133 -252 4139 -76
rect 4093 -264 4139 -252
rect -4083 -311 -2091 -305
rect -4083 -345 -4071 -311
rect -2103 -345 -2091 -311
rect -4083 -351 -2091 -345
rect -2025 -311 -33 -305
rect -2025 -345 -2013 -311
rect -45 -345 -33 -311
rect -2025 -351 -33 -345
rect 33 -311 2025 -305
rect 33 -345 45 -311
rect 2013 -345 2025 -311
rect 33 -351 2025 -345
rect 2091 -311 4083 -305
rect 2091 -345 2103 -311
rect 4071 -345 4083 -311
rect 2091 -351 4083 -345
<< labels >>
rlabel pdiffc -4116 -164 -4116 -164 0 D0_0
port 1 nsew
rlabel polycont -3087 0 -3087 0 0 G0
port 2 nsew
rlabel pdiffc -4116 164 -4116 164 0 D0_1
port 3 nsew
rlabel pdiffc -2058 -164 -2058 -164 0 S1_0
port 4 nsew
rlabel polycont -1029 0 -1029 0 0 G1
port 5 nsew
rlabel pdiffc -2058 164 -2058 164 0 S1_1
port 6 nsew
rlabel pdiffc 0 -164 0 -164 0 D2_0
port 7 nsew
rlabel polycont 1029 0 1029 0 0 G2
port 8 nsew
rlabel pdiffc 0 164 0 164 0 D2_1
port 9 nsew
rlabel pdiffc 2058 -164 2058 -164 0 S3_0
port 10 nsew
rlabel polycont 3087 0 3087 0 0 G3
port 11 nsew
rlabel pdiffc 2058 164 2058 164 0 S3_1
port 12 nsew
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 10 m 2 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 conn_gates 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 doports 1
<< end >>
