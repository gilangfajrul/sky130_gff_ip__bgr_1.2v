magic
tech sky130A
magscale 1 2
timestamp 1717917475
<< pwell >>
rect -31 2717 1533 15873
rect -31 2712 618 2717
rect 706 2712 1533 2717
rect -31 -51 1533 2712
<< metal1 >>
rect 311 15734 1440 15784
rect 311 15689 361 15734
rect 643 15689 693 15734
rect 1390 15701 1440 15734
rect 134 15637 144 15689
rect 196 15637 206 15689
rect 466 15637 476 15689
rect 528 15637 538 15689
rect 798 15637 808 15689
rect 860 15637 870 15689
rect 1141 15651 1440 15701
rect 964 15464 974 15516
rect 1026 15464 1036 15516
rect 964 13385 974 13437
rect 1026 13385 1036 13437
rect 134 13213 144 13265
rect 196 13213 206 13265
rect 466 13213 476 13265
rect 528 13213 538 13265
rect 798 13213 808 13265
rect 860 13213 870 13265
rect 1390 13251 1440 15651
rect 311 13168 361 13213
rect 643 13168 693 13213
rect 1143 13201 1440 13251
rect 62 13118 1191 13168
rect 62 13085 112 13118
rect 62 13035 360 13085
rect 477 13073 527 13118
rect 809 13073 859 13118
rect 1141 13073 1191 13118
rect 1390 13085 1440 13201
rect 62 10635 112 13035
rect 632 13021 642 13073
rect 694 13021 704 13073
rect 964 13021 974 13073
rect 1026 13021 1036 13073
rect 1307 13035 1440 13085
rect 62 10585 361 10635
rect 632 10597 642 10649
rect 694 10597 704 10649
rect 964 10597 974 10649
rect 1026 10597 1036 10649
rect 1390 10635 1440 13035
rect 62 10469 112 10585
rect 477 10552 527 10597
rect 809 10552 859 10597
rect 1141 10552 1191 10597
rect 1307 10585 1440 10635
rect 1390 10552 1440 10585
rect 311 10502 1440 10552
rect 62 10419 195 10469
rect 311 10457 361 10502
rect 643 10457 693 10502
rect 975 10457 1025 10502
rect 1390 10469 1440 10502
rect 62 8019 112 10419
rect 466 10405 476 10457
rect 528 10405 538 10457
rect 798 10405 808 10457
rect 860 10405 870 10457
rect 1141 10419 1440 10469
rect 1390 10023 1440 10419
rect 1379 8415 1389 10023
rect 1441 8415 1451 10023
rect 62 7969 195 8019
rect 466 7981 476 8033
rect 528 7981 538 8033
rect 798 7981 808 8033
rect 860 7981 870 8033
rect 1390 8019 1440 8415
rect 62 7936 112 7969
rect 311 7936 361 7981
rect 643 7936 693 7981
rect 975 7936 1025 7981
rect 1141 7969 1440 8019
rect 62 7886 1191 7936
rect 62 7853 112 7886
rect 62 7803 361 7853
rect 477 7841 527 7886
rect 809 7841 859 7886
rect 1141 7841 1191 7886
rect 1390 7853 1440 7969
rect 62 5403 112 7803
rect 632 7789 642 7841
rect 694 7789 704 7841
rect 964 7789 974 7841
rect 1026 7789 1036 7841
rect 1307 7803 1440 7853
rect 1390 7407 1440 7803
rect 1379 5799 1389 7407
rect 1441 5799 1451 7407
rect 62 5353 360 5403
rect 632 5365 642 5417
rect 694 5365 704 5417
rect 964 5365 974 5417
rect 1026 5365 1036 5417
rect 1390 5403 1440 5799
rect 62 5237 112 5353
rect 477 5320 527 5365
rect 809 5320 859 5365
rect 1141 5320 1191 5365
rect 1307 5353 1440 5403
rect 1390 5320 1440 5353
rect 311 5270 1440 5320
rect 62 5187 195 5237
rect 311 5225 361 5270
rect 643 5225 693 5270
rect 975 5225 1025 5270
rect 1390 5237 1440 5270
rect 62 2787 112 5187
rect 466 5173 476 5225
rect 528 5173 538 5225
rect 798 5173 808 5225
rect 860 5173 870 5225
rect 1141 5187 1440 5237
rect 62 2737 188 2787
rect 466 2749 476 2801
rect 528 2749 538 2801
rect 798 2749 808 2801
rect 860 2749 870 2801
rect 1390 2787 1440 5187
rect 62 2704 112 2737
rect 311 2704 361 2749
rect 643 2704 693 2749
rect 975 2704 1025 2749
rect 1141 2737 1440 2787
rect 62 2654 1191 2704
rect 145 2611 195 2654
rect 228 171 278 2654
rect 311 2613 361 2654
rect 809 2609 859 2654
rect 1141 2609 1191 2654
rect 1390 2621 1440 2737
rect 632 2557 642 2609
rect 694 2557 704 2609
rect 964 2557 974 2609
rect 1026 2557 1036 2609
rect 1307 2571 1440 2621
rect 466 2384 476 2436
rect 528 2384 538 2436
rect 466 305 476 357
rect 528 305 538 357
rect 145 121 346 171
rect 632 133 642 185
rect 694 133 704 185
rect 964 133 974 185
rect 1026 133 1036 185
rect 1390 171 1440 2571
rect 809 88 859 133
rect 1141 88 1191 133
rect 1307 121 1440 171
rect 1390 88 1440 121
rect 809 38 1440 88
<< via1 >>
rect 144 15637 196 15689
rect 476 15637 528 15689
rect 808 15637 860 15689
rect 974 15464 1026 15516
rect 974 13385 1026 13437
rect 144 13213 196 13265
rect 476 13213 528 13265
rect 808 13213 860 13265
rect 642 13021 694 13073
rect 974 13021 1026 13073
rect 642 10597 694 10649
rect 974 10597 1026 10649
rect 476 10405 528 10457
rect 808 10405 860 10457
rect 1389 8415 1441 10023
rect 476 7981 528 8033
rect 808 7981 860 8033
rect 642 7789 694 7841
rect 974 7789 1026 7841
rect 1389 5799 1441 7407
rect 642 5365 694 5417
rect 974 5365 1026 5417
rect 476 5173 528 5225
rect 808 5173 860 5225
rect 476 2749 528 2801
rect 808 2749 860 2801
rect 642 2557 694 2609
rect 974 2557 1026 2609
rect 476 2384 528 2436
rect 476 305 528 357
rect 642 133 694 185
rect 974 133 1026 185
<< metal2 >>
rect 61 15729 528 15781
rect 61 15699 113 15729
rect 61 15689 196 15699
rect 61 15637 144 15689
rect 61 15627 196 15637
rect 476 15689 528 15729
rect 476 15627 528 15637
rect 806 15691 862 15701
rect 61 13275 113 15627
rect 806 15625 862 15635
rect 972 15518 1028 15528
rect 972 15452 1028 15462
rect 972 13439 1028 13449
rect 972 13373 1028 13383
rect 61 13265 196 13275
rect 61 13213 144 13265
rect 61 13203 196 13213
rect 476 13265 528 13275
rect 61 10553 113 13203
rect 476 13169 528 13213
rect 806 13267 862 13277
rect 806 13201 862 13211
rect 476 13117 1441 13169
rect 642 13073 694 13117
rect 642 13011 694 13021
rect 972 13075 1028 13085
rect 972 13009 1028 13019
rect 642 10649 694 10659
rect 642 10553 694 10597
rect 972 10651 1028 10661
rect 972 10585 1028 10595
rect 61 10501 860 10553
rect 61 10033 113 10501
rect 476 10457 528 10501
rect 476 10395 528 10405
rect 808 10457 860 10501
rect 808 10395 860 10405
rect 54 10023 120 10033
rect 54 8405 120 8415
rect 1389 10023 1441 13117
rect 61 7417 113 8405
rect 476 8033 528 8043
rect 476 7937 528 7981
rect 808 8033 860 8043
rect 808 7937 860 7981
rect 1389 7937 1441 8415
rect 476 7885 1441 7937
rect 642 7841 694 7885
rect 642 7779 694 7789
rect 974 7841 1026 7885
rect 974 7779 1026 7789
rect 54 7407 120 7417
rect 54 5789 120 5799
rect 1389 7407 1441 7885
rect 61 5321 113 5789
rect 642 5417 694 5427
rect 642 5321 694 5365
rect 974 5417 1026 5427
rect 974 5321 1026 5365
rect 61 5269 1026 5321
rect 61 89 113 5269
rect 474 5227 530 5237
rect 474 5161 530 5171
rect 808 5225 860 5269
rect 808 5163 860 5173
rect 474 2803 530 2813
rect 474 2737 530 2747
rect 808 2801 860 2811
rect 808 2705 860 2749
rect 1389 2705 1441 5799
rect 808 2653 1441 2705
rect 640 2611 696 2621
rect 640 2545 696 2555
rect 974 2609 1026 2653
rect 974 2547 1026 2557
rect 474 2438 530 2448
rect 474 2372 530 2382
rect 474 359 530 369
rect 474 293 530 303
rect 640 187 696 197
rect 640 121 696 131
rect 974 185 1026 195
rect 974 89 1026 133
rect 61 37 1026 89
<< via2 >>
rect 806 15689 862 15691
rect 806 15637 808 15689
rect 808 15637 860 15689
rect 860 15637 862 15689
rect 806 15635 862 15637
rect 972 15516 1028 15518
rect 972 15464 974 15516
rect 974 15464 1026 15516
rect 1026 15464 1028 15516
rect 972 15462 1028 15464
rect 972 13437 1028 13439
rect 972 13385 974 13437
rect 974 13385 1026 13437
rect 1026 13385 1028 13437
rect 972 13383 1028 13385
rect 806 13265 862 13267
rect 806 13213 808 13265
rect 808 13213 860 13265
rect 860 13213 862 13265
rect 806 13211 862 13213
rect 972 13073 1028 13075
rect 972 13021 974 13073
rect 974 13021 1026 13073
rect 1026 13021 1028 13073
rect 972 13019 1028 13021
rect 972 10649 1028 10651
rect 972 10597 974 10649
rect 974 10597 1026 10649
rect 1026 10597 1028 10649
rect 972 10595 1028 10597
rect 54 8415 120 10023
rect 54 5799 120 7407
rect 474 5225 530 5227
rect 474 5173 476 5225
rect 476 5173 528 5225
rect 528 5173 530 5225
rect 474 5171 530 5173
rect 474 2801 530 2803
rect 474 2749 476 2801
rect 476 2749 528 2801
rect 528 2749 530 2801
rect 474 2747 530 2749
rect 640 2609 696 2611
rect 640 2557 642 2609
rect 642 2557 694 2609
rect 694 2557 696 2609
rect 640 2555 696 2557
rect 474 2436 530 2438
rect 474 2384 476 2436
rect 476 2384 528 2436
rect 528 2384 530 2436
rect 474 2382 530 2384
rect 474 357 530 359
rect 474 305 476 357
rect 476 305 528 357
rect 528 305 530 357
rect 474 303 530 305
rect 640 185 696 187
rect 640 133 642 185
rect 642 133 694 185
rect 694 133 696 185
rect 640 131 696 133
<< metal3 >>
rect 796 15717 1448 15793
rect 796 15691 872 15717
rect 796 15635 806 15691
rect 862 15635 872 15691
rect 796 15630 872 15635
rect 962 15522 1038 15567
rect 958 15458 968 15522
rect 1032 15458 1042 15522
rect 962 15413 1038 15458
rect 962 13443 1038 13488
rect 958 13379 968 13443
rect 1032 13379 1042 13443
rect 962 13334 1038 13379
rect 796 13267 950 13272
rect 796 13211 806 13267
rect 862 13211 950 13267
rect 796 13176 950 13211
rect 54 13110 1038 13176
rect 54 10028 120 13110
rect 884 13075 1038 13110
rect 884 13019 972 13075
rect 1028 13019 1038 13075
rect 884 13014 1038 13019
rect 962 10651 1038 10656
rect 962 10595 972 10651
rect 1028 10595 1038 10651
rect 962 10565 1038 10595
rect 1382 10565 1448 15717
rect 962 10489 1448 10565
rect 44 10023 130 10028
rect 1382 10023 1448 10489
rect 44 8415 54 10023
rect 120 8415 130 10023
rect 1372 8415 1382 10023
rect 1448 8415 1458 10023
rect 44 8410 130 8415
rect 54 7412 120 8410
rect 44 7407 130 7412
rect 1382 7407 1448 8415
rect 44 5799 54 7407
rect 120 5799 130 7407
rect 1372 5799 1382 7407
rect 1448 5799 1458 7407
rect 44 5794 130 5799
rect 54 2712 120 5794
rect 1382 5333 1448 5799
rect 464 5257 1448 5333
rect 464 5227 540 5257
rect 464 5171 474 5227
rect 530 5171 540 5227
rect 464 5166 540 5171
rect 464 2803 618 2808
rect 464 2747 474 2803
rect 530 2747 618 2803
rect 464 2712 618 2747
rect 54 2646 706 2712
rect 552 2611 706 2646
rect 552 2555 640 2611
rect 696 2555 706 2611
rect 552 2550 706 2555
rect 464 2442 540 2487
rect 460 2378 470 2442
rect 534 2378 544 2442
rect 464 2333 540 2378
rect 464 363 540 407
rect 460 299 470 363
rect 534 299 544 363
rect 464 254 540 299
rect 630 187 706 192
rect 630 131 640 187
rect 696 131 706 187
rect 630 105 706 131
rect 1382 105 1448 5257
rect 630 29 1448 105
<< via3 >>
rect 968 15518 1032 15522
rect 968 15462 972 15518
rect 972 15462 1028 15518
rect 1028 15462 1032 15518
rect 968 15458 1032 15462
rect 968 13439 1032 13443
rect 968 13383 972 13439
rect 972 13383 1028 13439
rect 1028 13383 1032 13439
rect 968 13379 1032 13383
rect 1382 8415 1448 10023
rect 1382 5799 1448 7407
rect 470 2438 534 2442
rect 470 2382 474 2438
rect 474 2382 530 2438
rect 530 2382 534 2438
rect 470 2378 534 2382
rect 470 359 534 363
rect 470 303 474 359
rect 474 303 530 359
rect 530 303 534 359
rect 470 299 534 303
<< metal4 >>
rect 54 15522 1033 15523
rect 54 15458 968 15522
rect 1032 15458 1033 15522
rect 54 15457 1033 15458
rect 54 364 120 15457
rect 967 13443 1448 13444
rect 967 13379 968 13443
rect 1032 13379 1448 13443
rect 967 13378 1448 13379
rect 1382 10024 1448 13378
rect 1381 10023 1449 10024
rect 1381 8415 1382 10023
rect 1448 8415 1449 10023
rect 1381 8414 1449 8415
rect 1382 7408 1448 8414
rect 1381 7407 1449 7408
rect 1381 5799 1382 7407
rect 1448 5799 1449 7407
rect 1381 5798 1449 5799
rect 1382 2443 1448 5798
rect 469 2442 1448 2443
rect 469 2378 470 2442
rect 534 2378 1448 2442
rect 469 2377 1448 2378
rect 54 363 535 364
rect 54 299 470 363
rect 534 299 535 363
rect 54 298 535 299
use sky130_fd_pr__res_high_po_0p35_KQ9YC9  sky130_fd_pr__res_high_po_0p35_KQ9YC9_0
timestamp 1717669726
transform 1 0 751 0 1 7911
box -782 -7962 782 7962
<< labels >>
flabel metal1 224 7908 224 7908 0 FreeSans 1600 0 0 0 B
port 0 nsew
flabel metal4 80 7474 80 7474 0 FreeSans 1600 0 0 0 A
port 1 nsew
flabel pwell 12 -35 12 -35 0 FreeSans 1600 0 0 0 AVSS
port 4 nsew
flabel metal4 1420 7946 1420 7946 0 FreeSans 1600 0 0 0 1
port 5 nsew
flabel metal3 118 8070 118 8070 0 FreeSans 1600 0 0 0 2
port 6 nsew
flabel metal2 1418 8274 1418 8274 0 FreeSans 1600 0 0 0 3
port 7 nsew
<< end >>
