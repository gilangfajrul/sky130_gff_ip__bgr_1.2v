magic
tech sky130A
magscale 1 2
timestamp 1718868641
<< viali >>
rect -17 1441 21819 1475
rect -17 17 17 1441
rect 21785 17 21819 1441
rect -17 -17 21819 17
<< metal1 >>
rect -23 1481 23 1487
rect 21779 1481 21825 1487
rect -29 1475 21831 1481
rect -29 1435 -17 1475
rect -23 23 -17 1435
rect -29 -17 -17 23
rect 17 1435 21785 1441
rect 17 23 23 1435
rect 119 1315 177 1435
rect 4327 1285 4467 1335
rect 8663 1285 8803 1335
rect 12999 1285 13139 1335
rect 17335 1285 17475 1335
rect 21625 1330 21683 1435
rect 119 1119 177 1169
rect 4327 1119 4467 1169
rect 8663 1119 8803 1169
rect 12999 1119 13139 1169
rect 17335 1119 17475 1169
rect 119 788 169 1004
rect 4327 953 4467 1003
rect 8663 953 8803 1003
rect 12999 953 13139 1003
rect 17335 953 17475 1003
rect 21633 953 21683 1169
rect 4327 787 4467 837
rect 8663 787 8803 837
rect 12999 787 13139 837
rect 17335 787 17475 837
rect 119 456 169 672
rect 4327 621 4467 671
rect 8663 621 8803 671
rect 12999 621 13139 671
rect 17335 621 17475 671
rect 21633 621 21683 837
rect 4327 455 4467 505
rect 8663 455 8803 505
rect 12999 455 13139 505
rect 17335 455 17475 505
rect 119 289 177 339
rect 4327 289 4467 339
rect 8663 289 8803 339
rect 12999 289 13139 339
rect 17335 289 17475 339
rect 21633 289 21683 505
rect 119 23 177 132
rect 4327 123 4467 173
rect 8663 123 8803 173
rect 12999 123 13139 173
rect 17335 123 17475 173
rect 21625 23 21684 128
rect 21779 23 21785 1435
rect 17 17 21785 23
rect 21819 1435 21831 1475
rect 21819 23 21825 1435
rect 21819 -17 21831 23
rect -29 -23 21831 -17
rect -23 -29 23 -23
rect 21779 -29 21825 -23
use sky130_fd_pr__res_high_po_0p35_9NXREG  sky130_fd_pr__res_high_po_0p35_9NXREG_0
timestamp 1717755416
transform 0 -1 10901 1 0 729
box -782 -10954 782 10954
<< labels >>
flabel metal1 124 314 124 314 0 FreeSans 1600 0 0 0 B
port 1 nsew
flabel metal1 125 1137 125 1137 0 FreeSans 1600 0 0 0 A
port 0 nsew
flabel metal1 21654 1388 21654 1388 0 FreeSans 1600 0 0 0 AVSS
port 3 nsew
<< end >>
