magic
tech sky130A
magscale 1 2
timestamp 1762701392
<< metal3 >>
rect -775 1694 528 1794
rect -766 -378 -666 32
rect 3732 -336 3832 74
rect -865 -2107 89 -2008
<< metal4 >>
rect -2810 -214 3990 -110
use sky130_fd_pr__cap_mim_m3_1_TVJG6P  sky130_fd_pr__cap_mim_m3_1_TVJG6P_0
timestamp 1762701392
transform 1 0 -333 0 1 -160
box -4165 -3800 4165 3800
<< labels >>
flabel metal4 3936 -161 3936 -161 0 FreeSans 160 0 0 0 A
port 0 nsew
flabel metal3 3777 -279 3777 -279 0 FreeSans 160 0 0 0 B
port 1 nsew
<< end >>
