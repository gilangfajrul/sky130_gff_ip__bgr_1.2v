magic
tech sky130A
magscale 1 2
timestamp 1716365683
<< metal3 >>
rect -7904 6492 -4132 6520
rect -7904 3468 -4216 6492
rect -4152 3468 -4132 6492
rect -7904 3440 -4132 3468
rect -3892 6492 -120 6520
rect -3892 3468 -204 6492
rect -140 3468 -120 6492
rect -3892 3440 -120 3468
rect 120 6492 3892 6520
rect 120 3468 3808 6492
rect 3872 3468 3892 6492
rect 120 3440 3892 3468
rect 4132 6492 7904 6520
rect 4132 3468 7820 6492
rect 7884 3468 7904 6492
rect 4132 3440 7904 3468
rect -7904 3172 -4132 3200
rect -7904 148 -4216 3172
rect -4152 148 -4132 3172
rect -7904 120 -4132 148
rect -3892 3172 -120 3200
rect -3892 148 -204 3172
rect -140 148 -120 3172
rect -3892 120 -120 148
rect 120 3172 3892 3200
rect 120 148 3808 3172
rect 3872 148 3892 3172
rect 120 120 3892 148
rect 4132 3172 7904 3200
rect 4132 148 7820 3172
rect 7884 148 7904 3172
rect 4132 120 7904 148
rect -7904 -148 -4132 -120
rect -7904 -3172 -4216 -148
rect -4152 -3172 -4132 -148
rect -7904 -3200 -4132 -3172
rect -3892 -148 -120 -120
rect -3892 -3172 -204 -148
rect -140 -3172 -120 -148
rect -3892 -3200 -120 -3172
rect 120 -148 3892 -120
rect 120 -3172 3808 -148
rect 3872 -3172 3892 -148
rect 120 -3200 3892 -3172
rect 4132 -148 7904 -120
rect 4132 -3172 7820 -148
rect 7884 -3172 7904 -148
rect 4132 -3200 7904 -3172
rect -7904 -3468 -4132 -3440
rect -7904 -6492 -4216 -3468
rect -4152 -6492 -4132 -3468
rect -7904 -6520 -4132 -6492
rect -3892 -3468 -120 -3440
rect -3892 -6492 -204 -3468
rect -140 -6492 -120 -3468
rect -3892 -6520 -120 -6492
rect 120 -3468 3892 -3440
rect 120 -6492 3808 -3468
rect 3872 -6492 3892 -3468
rect 120 -6520 3892 -6492
rect 4132 -3468 7904 -3440
rect 4132 -6492 7820 -3468
rect 7884 -6492 7904 -3468
rect 4132 -6520 7904 -6492
<< via3 >>
rect -4216 3468 -4152 6492
rect -204 3468 -140 6492
rect 3808 3468 3872 6492
rect 7820 3468 7884 6492
rect -4216 148 -4152 3172
rect -204 148 -140 3172
rect 3808 148 3872 3172
rect 7820 148 7884 3172
rect -4216 -3172 -4152 -148
rect -204 -3172 -140 -148
rect 3808 -3172 3872 -148
rect 7820 -3172 7884 -148
rect -4216 -6492 -4152 -3468
rect -204 -6492 -140 -3468
rect 3808 -6492 3872 -3468
rect 7820 -6492 7884 -3468
<< mimcap >>
rect -7864 6440 -4464 6480
rect -7864 3520 -7824 6440
rect -4504 3520 -4464 6440
rect -7864 3480 -4464 3520
rect -3852 6440 -452 6480
rect -3852 3520 -3812 6440
rect -492 3520 -452 6440
rect -3852 3480 -452 3520
rect 160 6440 3560 6480
rect 160 3520 200 6440
rect 3520 3520 3560 6440
rect 160 3480 3560 3520
rect 4172 6440 7572 6480
rect 4172 3520 4212 6440
rect 7532 3520 7572 6440
rect 4172 3480 7572 3520
rect -7864 3120 -4464 3160
rect -7864 200 -7824 3120
rect -4504 200 -4464 3120
rect -7864 160 -4464 200
rect -3852 3120 -452 3160
rect -3852 200 -3812 3120
rect -492 200 -452 3120
rect -3852 160 -452 200
rect 160 3120 3560 3160
rect 160 200 200 3120
rect 3520 200 3560 3120
rect 160 160 3560 200
rect 4172 3120 7572 3160
rect 4172 200 4212 3120
rect 7532 200 7572 3120
rect 4172 160 7572 200
rect -7864 -200 -4464 -160
rect -7864 -3120 -7824 -200
rect -4504 -3120 -4464 -200
rect -7864 -3160 -4464 -3120
rect -3852 -200 -452 -160
rect -3852 -3120 -3812 -200
rect -492 -3120 -452 -200
rect -3852 -3160 -452 -3120
rect 160 -200 3560 -160
rect 160 -3120 200 -200
rect 3520 -3120 3560 -200
rect 160 -3160 3560 -3120
rect 4172 -200 7572 -160
rect 4172 -3120 4212 -200
rect 7532 -3120 7572 -200
rect 4172 -3160 7572 -3120
rect -7864 -3520 -4464 -3480
rect -7864 -6440 -7824 -3520
rect -4504 -6440 -4464 -3520
rect -7864 -6480 -4464 -6440
rect -3852 -3520 -452 -3480
rect -3852 -6440 -3812 -3520
rect -492 -6440 -452 -3520
rect -3852 -6480 -452 -6440
rect 160 -3520 3560 -3480
rect 160 -6440 200 -3520
rect 3520 -6440 3560 -3520
rect 160 -6480 3560 -6440
rect 4172 -3520 7572 -3480
rect 4172 -6440 4212 -3520
rect 7532 -6440 7572 -3520
rect 4172 -6480 7572 -6440
<< mimcapcontact >>
rect -7824 3520 -4504 6440
rect -3812 3520 -492 6440
rect 200 3520 3520 6440
rect 4212 3520 7532 6440
rect -7824 200 -4504 3120
rect -3812 200 -492 3120
rect 200 200 3520 3120
rect 4212 200 7532 3120
rect -7824 -3120 -4504 -200
rect -3812 -3120 -492 -200
rect 200 -3120 3520 -200
rect 4212 -3120 7532 -200
rect -7824 -6440 -4504 -3520
rect -3812 -6440 -492 -3520
rect 200 -6440 3520 -3520
rect 4212 -6440 7532 -3520
<< metal4 >>
rect -4232 6492 -4136 6508
rect -7825 6440 -4503 6441
rect -7825 3520 -7824 6440
rect -4504 3520 -4503 6440
rect -7825 3519 -4503 3520
rect -4232 3468 -4216 6492
rect -4152 3468 -4136 6492
rect -220 6492 -124 6508
rect -3813 6440 -491 6441
rect -3813 3520 -3812 6440
rect -492 3520 -491 6440
rect -3813 3519 -491 3520
rect -4232 3452 -4136 3468
rect -220 3468 -204 6492
rect -140 3468 -124 6492
rect 3792 6492 3888 6508
rect 199 6440 3521 6441
rect 199 3520 200 6440
rect 3520 3520 3521 6440
rect 199 3519 3521 3520
rect -220 3452 -124 3468
rect 3792 3468 3808 6492
rect 3872 3468 3888 6492
rect 7804 6492 7900 6508
rect 4211 6440 7533 6441
rect 4211 3520 4212 6440
rect 7532 3520 7533 6440
rect 4211 3519 7533 3520
rect 3792 3452 3888 3468
rect 7804 3468 7820 6492
rect 7884 3468 7900 6492
rect 7804 3452 7900 3468
rect -4232 3172 -4136 3188
rect -7825 3120 -4503 3121
rect -7825 200 -7824 3120
rect -4504 200 -4503 3120
rect -7825 199 -4503 200
rect -4232 148 -4216 3172
rect -4152 148 -4136 3172
rect -220 3172 -124 3188
rect -3813 3120 -491 3121
rect -3813 200 -3812 3120
rect -492 200 -491 3120
rect -3813 199 -491 200
rect -4232 132 -4136 148
rect -220 148 -204 3172
rect -140 148 -124 3172
rect 3792 3172 3888 3188
rect 199 3120 3521 3121
rect 199 200 200 3120
rect 3520 200 3521 3120
rect 199 199 3521 200
rect -220 132 -124 148
rect 3792 148 3808 3172
rect 3872 148 3888 3172
rect 7804 3172 7900 3188
rect 4211 3120 7533 3121
rect 4211 200 4212 3120
rect 7532 200 7533 3120
rect 4211 199 7533 200
rect 3792 132 3888 148
rect 7804 148 7820 3172
rect 7884 148 7900 3172
rect 7804 132 7900 148
rect -4232 -148 -4136 -132
rect -7825 -200 -4503 -199
rect -7825 -3120 -7824 -200
rect -4504 -3120 -4503 -200
rect -7825 -3121 -4503 -3120
rect -4232 -3172 -4216 -148
rect -4152 -3172 -4136 -148
rect -220 -148 -124 -132
rect -3813 -200 -491 -199
rect -3813 -3120 -3812 -200
rect -492 -3120 -491 -200
rect -3813 -3121 -491 -3120
rect -4232 -3188 -4136 -3172
rect -220 -3172 -204 -148
rect -140 -3172 -124 -148
rect 3792 -148 3888 -132
rect 199 -200 3521 -199
rect 199 -3120 200 -200
rect 3520 -3120 3521 -200
rect 199 -3121 3521 -3120
rect -220 -3188 -124 -3172
rect 3792 -3172 3808 -148
rect 3872 -3172 3888 -148
rect 7804 -148 7900 -132
rect 4211 -200 7533 -199
rect 4211 -3120 4212 -200
rect 7532 -3120 7533 -200
rect 4211 -3121 7533 -3120
rect 3792 -3188 3888 -3172
rect 7804 -3172 7820 -148
rect 7884 -3172 7900 -148
rect 7804 -3188 7900 -3172
rect -4232 -3468 -4136 -3452
rect -7825 -3520 -4503 -3519
rect -7825 -6440 -7824 -3520
rect -4504 -6440 -4503 -3520
rect -7825 -6441 -4503 -6440
rect -4232 -6492 -4216 -3468
rect -4152 -6492 -4136 -3468
rect -220 -3468 -124 -3452
rect -3813 -3520 -491 -3519
rect -3813 -6440 -3812 -3520
rect -492 -6440 -491 -3520
rect -3813 -6441 -491 -6440
rect -4232 -6508 -4136 -6492
rect -220 -6492 -204 -3468
rect -140 -6492 -124 -3468
rect 3792 -3468 3888 -3452
rect 199 -3520 3521 -3519
rect 199 -6440 200 -3520
rect 3520 -6440 3521 -3520
rect 199 -6441 3521 -6440
rect -220 -6508 -124 -6492
rect 3792 -6492 3808 -3468
rect 3872 -6492 3888 -3468
rect 7804 -3468 7900 -3452
rect 4211 -3520 7533 -3519
rect 4211 -6440 4212 -3520
rect 7532 -6440 7533 -3520
rect 4211 -6441 7533 -6440
rect 3792 -6508 3888 -6492
rect 7804 -6492 7820 -3468
rect 7884 -6492 7900 -3468
rect 7804 -6508 7900 -6492
<< properties >>
string FIXED_BBOX 4132 3440 7612 6520
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 17 l 15 val 522.159 carea 2.00 cperi 0.19 nx 4 ny 4 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 0 tconnect 0 ccov 100
<< end >>
