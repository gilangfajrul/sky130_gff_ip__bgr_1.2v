magic
tech sky130A
magscale 1 2
timestamp 1717249874
<< psubdiff >>
rect -309 1533 -249 1567
rect 8527 1533 8587 1567
rect -309 1485 -275 1533
rect 8553 1485 8587 1533
rect -309 -95 -275 -69
rect 8553 -95 8587 -69
rect -309 -129 -249 -95
rect 8527 -129 8587 -95
<< psubdiffcont >>
rect -249 1533 8527 1567
rect -309 -69 -275 1485
rect 8553 -69 8587 1485
rect -249 -129 8527 -95
<< poly >>
rect -208 1483 -116 1499
rect -208 1449 -192 1483
rect -158 1449 -116 1483
rect -208 1433 -116 1449
rect 8394 1187 8424 1210
rect 54 1042 8224 1184
rect 8394 1171 8486 1187
rect 8394 1137 8436 1171
rect 8470 1137 8486 1171
rect 8394 1121 8486 1137
rect -146 793 -116 816
rect -208 777 -116 793
rect 8394 793 8424 816
rect -208 743 -192 777
rect -158 743 -116 777
rect -208 695 -116 743
rect -208 661 -192 695
rect -158 661 -116 695
rect -208 645 -116 661
rect 54 648 8224 790
rect 8394 777 8486 793
rect 8394 743 8436 777
rect 8470 743 8486 777
rect 8394 695 8486 743
rect 8394 661 8436 695
rect 8470 661 8486 695
rect -146 622 -116 645
rect 8394 645 8486 661
rect 8394 622 8424 645
rect 54 254 8224 396
rect -146 5 -116 28
rect -208 -11 -116 5
rect -208 -45 -192 -11
rect -158 -45 -116 -11
rect -208 -61 -116 -45
rect 8394 5 8424 28
rect 8394 -11 8486 5
rect 8394 -45 8436 -11
rect 8470 -45 8486 -11
rect 8394 -61 8486 -45
<< polycont >>
rect -192 1449 -158 1483
rect 8436 1137 8470 1171
rect -192 743 -158 777
rect -192 661 -158 695
rect 8436 743 8470 777
rect 8436 661 8470 695
rect -192 -45 -158 -11
rect 8436 -45 8470 -11
<< locali >>
rect -309 1533 -249 1567
rect 8527 1533 8587 1567
rect -309 1485 -275 1533
rect -192 1483 -158 1499
rect -192 1410 -158 1449
rect 8553 1485 8587 1533
rect 8436 1171 8470 1210
rect 8436 1121 8470 1137
rect -192 777 -158 816
rect -192 695 -158 743
rect -192 622 -158 661
rect 8436 777 8470 816
rect 8436 695 8470 743
rect 8436 622 8470 661
rect -192 -11 -158 28
rect -192 -61 -158 -45
rect 8436 -11 8470 28
rect 8436 -61 8470 -45
rect -309 -95 -275 -69
rect 8553 -95 8587 -69
rect -309 -129 -249 -95
rect 8527 -129 8587 -95
<< viali >>
rect 4178 1533 4212 1567
rect -309 1449 -275 1483
rect -192 1449 -158 1483
rect 8436 1137 8470 1171
rect 8553 1137 8587 1171
rect -309 702 -275 736
rect -192 743 -158 777
rect -192 661 -158 695
rect 8436 743 8470 777
rect 8436 661 8470 695
rect 8553 702 8587 736
rect -309 -45 -275 -11
rect -192 -45 -158 -11
rect 8436 -45 8470 -11
rect 8553 -45 8587 -11
rect 4066 -129 4100 -95
<< metal1 >>
rect 4172 1567 4218 1579
rect 4172 1533 4178 1567
rect 4212 1533 4218 1567
rect -315 1483 -152 1495
rect -315 1449 -309 1483
rect -275 1449 -192 1483
rect -158 1449 -152 1483
rect -315 1437 -152 1449
rect -198 1408 -152 1437
rect 8 1442 1089 1488
rect 8 1410 42 1442
rect -110 1210 48 1410
rect 4172 1407 4218 1533
rect 8230 1398 8388 1410
rect 4047 1222 4057 1398
rect 4109 1222 4119 1398
rect 8230 1222 8283 1398
rect 8335 1222 8388 1398
rect 4172 1016 4218 1222
rect 8230 1210 8388 1222
rect 8430 1183 8476 1210
rect 8430 1171 8593 1183
rect 8430 1137 8436 1171
rect 8470 1137 8553 1171
rect 8587 1137 8593 1171
rect 8430 1125 8593 1137
rect -110 1004 48 1016
rect -110 828 -57 1004
rect -5 828 48 1004
rect -110 816 48 828
rect -198 777 -152 816
rect -198 748 -192 777
rect -315 743 -192 748
rect -158 743 -152 777
rect -315 736 -152 743
rect -315 702 -309 736
rect -275 702 -152 736
rect -315 695 -152 702
rect -315 690 -192 695
rect -198 661 -192 690
rect -158 661 -152 695
rect -198 622 -152 661
rect -110 610 48 622
rect -110 434 -57 610
rect -5 434 48 610
rect -110 422 48 434
rect 4060 422 4218 1016
rect 8230 1004 8388 1016
rect 8230 828 8283 1004
rect 8335 828 8388 1004
rect 8230 820 8388 828
rect 8230 816 8387 820
rect 8430 777 8476 816
rect 8430 743 8436 777
rect 8470 748 8476 777
rect 8470 743 8593 748
rect 8430 736 8593 743
rect 8430 702 8553 736
rect 8587 702 8593 736
rect 8430 695 8593 702
rect 8430 661 8436 695
rect 8470 690 8593 695
rect 8470 661 8476 690
rect 8430 622 8476 661
rect 8230 610 8388 622
rect 8230 434 8283 610
rect 8335 434 8388 610
rect 8230 422 8388 434
rect -110 216 48 228
rect 4060 223 4106 422
rect -110 40 -57 216
rect -5 40 48 216
rect 4159 40 4169 216
rect 4221 40 4231 216
rect -110 28 48 40
rect -198 1 -152 28
rect -315 -11 -152 1
rect -315 -45 -309 -11
rect -275 -45 -192 -11
rect -158 -45 -152 -11
rect -315 -57 -152 -45
rect 4060 -95 4106 36
rect 8230 28 8388 228
rect 8236 -4 8270 28
rect 7161 -50 8270 -4
rect 8430 1 8476 28
rect 8430 -11 8593 1
rect 8430 -45 8436 -11
rect 8470 -45 8553 -11
rect 8587 -45 8593 -11
rect 8430 -57 8593 -45
rect 4060 -129 4066 -95
rect 4100 -129 4106 -95
rect 4060 -141 4106 -129
<< via1 >>
rect 4057 1222 4109 1398
rect 8283 1222 8335 1398
rect -57 828 -5 1004
rect -57 434 -5 610
rect 8283 828 8335 1004
rect 8283 434 8335 610
rect -57 40 -5 216
rect 4169 40 4221 216
<< metal2 >>
rect 4055 1398 4111 1408
rect 4055 1212 4111 1222
rect 8283 1398 8335 1408
rect 8283 1139 8335 1222
rect -270 1087 8548 1139
rect -270 351 -218 1087
rect -57 1004 -5 1014
rect -57 745 -5 828
rect 8281 1004 8337 1014
rect 8281 818 8337 828
rect -57 693 8335 745
rect -59 610 -3 620
rect -59 424 -3 434
rect 8283 610 8335 693
rect 8283 424 8335 434
rect 8496 351 8548 1087
rect -270 299 8548 351
rect -57 216 -5 299
rect -57 30 -5 40
rect 4167 216 4223 226
rect 4167 30 4223 40
<< via2 >>
rect 4055 1222 4057 1398
rect 4057 1222 4109 1398
rect 4109 1222 4111 1398
rect 8281 828 8283 1004
rect 8283 828 8335 1004
rect 8335 828 8337 1004
rect -59 434 -57 610
rect -57 434 -5 610
rect -5 434 -3 610
rect 4167 40 4169 216
rect 4169 40 4221 216
rect 4221 40 4223 216
<< metal3 >>
rect 4045 1398 4121 1403
rect 4041 1222 4051 1398
rect 4115 1222 4125 1398
rect 4045 1217 4121 1222
rect 8271 1004 8347 1009
rect 8271 828 8281 1004
rect 8337 828 8347 1004
rect 8271 823 8347 828
rect 8279 749 8339 823
rect -61 689 8339 749
rect -61 615 -1 689
rect -69 610 7 615
rect -69 434 -59 610
rect -3 434 7 610
rect -69 429 7 434
rect 4157 216 4233 221
rect 4153 40 4163 216
rect 4227 40 4237 216
rect 4157 35 4233 40
<< via3 >>
rect 4051 1222 4055 1398
rect 4055 1222 4111 1398
rect 4111 1222 4115 1398
rect 4163 40 4167 216
rect 4167 40 4223 216
rect 4223 40 4227 216
<< metal4 >>
rect 4050 1398 4170 1399
rect 4050 1222 4051 1398
rect 4115 1222 4170 1398
rect 4050 1221 4170 1222
rect 4108 217 4170 1221
rect 4108 216 4228 217
rect 4108 40 4163 216
rect 4227 40 4228 216
rect 4108 39 4228 40
use sky130_fd_pr__nfet_01v8_3KF9AC  sky130_fd_pr__nfet_01v8_3KF9AC_0
timestamp 1717076529
transform 1 0 2054 0 1 1341
box -2058 -157 2058 157
use sky130_fd_pr__nfet_01v8_3YKU97  sky130_fd_pr__nfet_01v8_3YKU97_0
timestamp 1717076529
transform 1 0 6224 0 1 97
box -2058 -157 2058 157
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_0
timestamp 1717248107
transform 1 0 -131 0 1 916
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_1
timestamp 1717248107
transform 1 0 -131 0 1 1308
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_2
timestamp 1717248107
transform 1 0 -131 0 1 522
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_3
timestamp 1717248107
transform 1 0 -131 0 1 128
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_4
timestamp 1717248107
transform 1 0 8409 0 1 128
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_5
timestamp 1717248107
transform 1 0 8409 0 1 522
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_6
timestamp 1717248107
transform 1 0 8409 0 1 916
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_7
timestamp 1717248107
transform 1 0 8409 0 1 1310
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_BSRS8Q  sky130_fd_pr__nfet_01v8_BSRS8Q_0
timestamp 1717249617
transform 1 0 6224 0 1 1310
box -2058 -126 2058 126
use sky130_fd_pr__nfet_01v8_P5G96Q  sky130_fd_pr__nfet_01v8_P5G96Q_1
timestamp 1716212328
transform 1 0 2054 0 1 128
box -2058 -126 2058 126
use sky130_fd_pr__nfet_01v8_P5G96Q  sky130_fd_pr__nfet_01v8_P5G96Q_4
timestamp 1716212328
transform 1 0 6224 0 1 522
box -2058 -126 2058 126
use sky130_fd_pr__nfet_01v8_P5G96Q  sky130_fd_pr__nfet_01v8_P5G96Q_5
timestamp 1716212328
transform 1 0 2054 0 1 522
box -2058 -126 2058 126
use sky130_fd_pr__nfet_01v8_P5G96Q  sky130_fd_pr__nfet_01v8_P5G96Q_6
timestamp 1716212328
transform 1 0 6224 0 1 916
box -2058 -126 2058 126
use sky130_fd_pr__nfet_01v8_P5G96Q  sky130_fd_pr__nfet_01v8_P5G96Q_7
timestamp 1716212328
transform 1 0 2054 0 1 916
box -2058 -126 2058 126
<< labels >>
flabel metal4 4130 186 4130 186 0 FreeSans 160 0 0 0 S2
port 6 nsew
flabel metal1 8516 -20 8516 -20 0 FreeSans 160 0 0 0 GND
port 4 nsew
flabel metal1 8310 134 8310 134 0 FreeSans 160 0 0 0 D2
port 3 nsew
flabel metal2 8302 652 8302 652 0 FreeSans 160 0 0 0 D3
port 2 nsew
flabel metal3 8310 784 8310 784 0 FreeSans 160 0 0 0 D4
port 1 nsew
flabel metal2 8306 1160 8306 1160 0 FreeSans 160 0 0 0 D1
port 0 nsew
<< end >>
