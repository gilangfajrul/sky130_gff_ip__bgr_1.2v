magic
tech sky130A
magscale 1 2
timestamp 1720284839
<< psubdiff >>
rect -405 6046 -345 6080
rect 695 6046 755 6080
rect -405 6020 -371 6046
rect -405 2266 -371 2292
rect 721 6020 755 6046
rect 721 2266 755 2292
rect -405 2232 -345 2266
rect 695 2232 755 2266
<< psubdiffcont >>
rect -345 6046 695 6080
rect -405 2292 -371 6020
rect 721 2292 755 6020
rect -345 2232 695 2266
<< viali >>
rect -405 6046 -345 6080
rect -345 6046 695 6080
rect 695 6046 755 6080
rect -405 6020 -371 6046
rect -405 2292 -371 6020
rect -405 2266 -371 2292
rect 721 6020 755 6046
rect 721 2292 755 6020
rect 721 2266 755 2292
rect -405 2232 -345 2266
rect -345 2232 695 2266
rect 695 2232 755 2266
<< metal1 >>
rect -411 6086 -365 6092
rect 715 6086 761 6092
rect -417 6080 767 6086
rect -417 6040 -405 6080
rect -411 2272 -405 6040
rect -417 2232 -405 2272
rect -371 6040 721 6046
rect -371 2272 -365 6040
rect -265 5919 -215 6040
rect 67 5962 283 6012
rect 67 5922 117 5962
rect 233 5922 283 5962
rect 565 5922 615 6040
rect -110 5870 -100 5922
rect -48 5870 -38 5922
rect 388 5870 398 5922
rect 450 5870 460 5922
rect -265 4096 -215 4250
rect 56 4226 66 4278
rect 118 4226 128 4278
rect 222 4226 232 4278
rect 284 4226 294 4278
rect -99 4181 -49 4224
rect 399 4181 449 4227
rect -99 4131 449 4181
rect -100 4086 -48 4096
rect 67 4095 117 4131
rect 233 4098 283 4131
rect 565 4092 615 4239
rect 388 4034 398 4086
rect 450 4034 460 4086
rect -100 4024 -48 4034
rect -100 2442 -48 2452
rect -265 2272 -215 2384
rect -100 2380 -48 2390
rect 67 2350 117 2400
rect 233 2350 283 2400
rect 388 2388 398 2440
rect 450 2388 460 2440
rect 67 2300 283 2350
rect 565 2272 615 2396
rect 715 2272 721 6040
rect -371 2266 721 2272
rect 755 6040 767 6080
rect 755 2272 761 6040
rect 755 2232 767 2272
rect -417 2226 767 2232
rect -411 2220 -365 2226
rect 715 2220 761 2226
<< via1 >>
rect -100 5870 -48 5922
rect 398 5870 450 5922
rect 66 4226 118 4278
rect 232 4226 284 4278
rect -100 4034 -48 4086
rect 398 4034 450 4086
rect -100 2390 -48 2442
rect 398 2388 450 2440
<< metal2 >>
rect -110 5960 460 6012
rect -110 5922 -38 5960
rect -110 5870 -100 5922
rect -48 5870 -38 5922
rect -110 5860 -38 5870
rect 388 5922 460 5960
rect 388 5870 398 5922
rect 450 5870 460 5922
rect 388 5860 460 5870
rect 66 4278 118 4288
rect 66 4182 118 4226
rect 232 4278 284 4288
rect 232 4182 284 4226
rect -110 4130 450 4182
rect -110 4086 -38 4130
rect -110 4034 -100 4086
rect -48 4034 -38 4086
rect 398 4086 450 4130
rect 398 4024 450 4034
rect -110 2390 -100 2442
rect -48 2390 -38 2442
rect -110 2352 -38 2390
rect 398 2440 450 2450
rect 398 2352 450 2388
rect -110 2300 450 2352
use sky130_fd_pr__res_high_po_0p35_RXTQM4  sky130_fd_pr__res_high_po_0p35_RXTQM4_0
timestamp 1720284156
transform 1 0 175 0 1 4156
box -450 -1784 450 1784
<< labels >>
flabel metal2 318 2324 318 2324 0 FreeSans 160 0 0 0 A
port 1 nsew
flabel metal1 252 2360 252 2360 0 FreeSans 160 0 0 0 C
port 2 nsew
flabel metal1 257 5949 257 5949 0 FreeSans 160 0 0 0 B
port 3 nsew
flabel metal2 327 5983 327 5983 0 FreeSans 160 0 0 0 D
port 4 nsew
flabel metal1 -245 2304 -245 2304 0 FreeSans 160 0 0 0 AVSS
port 5 nsew
<< end >>
