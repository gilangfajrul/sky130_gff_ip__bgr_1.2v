magic
tech sky130A
magscale 1 2
timestamp 1716365683
<< metal3 >>
rect -1886 212 1886 240
rect -1886 -212 1802 212
rect 1866 -212 1886 212
rect -1886 -240 1886 -212
<< via3 >>
rect 1802 -212 1866 212
<< mimcap >>
rect -1846 160 1554 200
rect -1846 -160 -1806 160
rect 1514 -160 1554 160
rect -1846 -200 1554 -160
<< mimcapcontact >>
rect -1806 -160 1514 160
<< metal4 >>
rect 1786 212 1882 228
rect -1807 160 1515 161
rect -1807 -160 -1806 160
rect 1514 -160 1515 160
rect -1807 -161 1515 -160
rect 1786 -212 1802 212
rect 1866 -212 1882 212
rect 1786 -228 1882 -212
<< properties >>
string FIXED_BBOX -1886 -240 1594 240
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 17 l 2.00 val 75.22 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
