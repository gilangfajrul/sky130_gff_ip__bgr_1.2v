magic
tech sky130A
magscale 1 2
timestamp 1717437593
<< nwell >>
rect -227 -1446 8585 509
<< nsubdiff >>
rect -191 439 -131 473
rect 8489 439 8549 473
rect -191 413 -157 439
rect 8515 413 8549 439
rect -191 -1376 -157 -1350
rect 8515 -1376 8549 -1350
rect -191 -1410 -131 -1376
rect 8489 -1410 8549 -1376
<< nsubdiffcont >>
rect -131 439 8489 473
rect -191 -1350 -157 413
rect 8515 -1350 8549 413
rect -131 -1410 8489 -1376
<< poly >>
rect -58 379 34 395
rect -58 345 -42 379
rect -8 345 34 379
rect -58 329 34 345
rect 4 321 34 329
rect 8324 379 8416 395
rect 8324 345 8366 379
rect 8400 345 8416 379
rect 8324 329 8416 345
rect 8324 298 8354 329
rect 4 -436 34 -348
rect -58 -452 34 -436
rect -58 -486 -42 -452
rect -8 -486 34 -452
rect -58 -502 34 -486
rect 4 -592 34 -502
rect 92 -540 8266 -398
rect 8324 -436 8354 -346
rect 8324 -452 8416 -436
rect 8324 -486 8366 -452
rect 8400 -486 8416 -452
rect 8324 -502 8416 -486
rect 8324 -578 8354 -502
rect 4 -1267 34 -1251
rect -58 -1283 34 -1267
rect -58 -1317 -42 -1283
rect -8 -1317 34 -1283
rect -58 -1333 34 -1317
rect 8324 -1267 8354 -1236
rect 8324 -1283 8416 -1267
rect 8324 -1317 8366 -1283
rect 8400 -1317 8416 -1283
rect 8324 -1333 8416 -1317
<< polycont >>
rect -42 345 -8 379
rect 8366 345 8400 379
rect -42 -486 -8 -452
rect 8366 -486 8400 -452
rect -42 -1317 -8 -1283
rect 8366 -1317 8400 -1283
<< locali >>
rect -191 439 -131 473
rect 8489 439 8549 473
rect -191 413 -157 439
rect 8515 413 8549 439
rect -42 379 -8 395
rect -42 296 -8 345
rect 8366 379 8400 395
rect 8366 298 8400 345
rect -42 -452 -8 -436
rect -42 -502 -8 -486
rect 8366 -452 8400 -436
rect 8366 -502 8400 -486
rect -42 -1283 -8 -1239
rect -42 -1333 -8 -1317
rect 8366 -1283 8400 -1236
rect 8366 -1333 8400 -1317
rect -191 -1376 -157 -1350
rect 8515 -1376 8549 -1350
rect -191 -1410 -131 -1376
rect 8489 -1410 8549 -1376
<< viali >>
rect -42 439 -8 473
rect 2104 439 2138 473
rect 4162 439 4196 473
rect 6220 439 6254 473
rect 8366 439 8400 473
rect -42 345 -8 379
rect 8366 345 8400 379
rect -191 -486 -157 -452
rect -42 -486 -8 -452
rect 8366 -486 8400 -452
rect 8515 -486 8549 -452
rect -42 -1317 -8 -1283
rect 8366 -1317 8400 -1283
rect -42 -1410 -8 -1376
rect 2104 -1410 2138 -1376
rect 4162 -1410 4196 -1376
rect 6220 -1410 6254 -1376
rect 8366 -1410 8400 -1376
<< metal1 >>
rect -48 473 -2 485
rect -48 439 -42 473
rect -8 439 -2 473
rect -48 379 -2 439
rect -48 345 -42 379
rect -8 345 -2 379
rect -48 295 -2 345
rect 2098 473 2144 485
rect 2098 439 2104 473
rect 2138 439 2144 473
rect 2098 286 2144 439
rect 4156 473 4202 485
rect 4156 439 4162 473
rect 4196 439 4202 473
rect 27 110 37 286
rect 89 110 99 286
rect 2085 110 2095 286
rect 2147 110 2157 286
rect 4156 280 4202 439
rect 6214 473 6260 485
rect 6214 439 6220 473
rect 6254 439 6260 473
rect 6214 286 6260 439
rect 8360 473 8406 485
rect 8360 439 8366 473
rect 8400 439 8406 473
rect 8360 379 8406 439
rect 8360 345 8366 379
rect 8400 345 8406 379
rect 8360 298 8406 345
rect 6201 110 6211 286
rect 6263 110 6273 286
rect 8259 110 8269 286
rect 8321 110 8331 286
rect 4156 57 4202 105
rect -152 -66 -142 -14
rect -90 -17 -80 -14
rect 588 -17 1596 20
rect 3633 11 4730 57
rect 6762 -17 7770 15
rect 8438 -17 8448 -14
rect -90 -63 8448 -17
rect -90 -66 -80 -63
rect 8438 -66 8448 -63
rect 8500 -66 8510 -14
rect -48 -440 -2 -313
rect -197 -452 -2 -440
rect 40 -443 86 -320
rect 2085 -322 2095 -146
rect 2147 -322 2157 -146
rect 4143 -322 4153 -146
rect 4205 -322 4215 -146
rect 6201 -322 6211 -146
rect 6263 -322 6273 -146
rect -197 -486 -191 -452
rect -157 -486 -42 -452
rect -8 -486 -2 -452
rect -197 -498 -2 -486
rect 27 -495 37 -443
rect 89 -495 99 -443
rect 588 -452 1596 -414
rect 6762 -452 7770 -419
rect 8272 -443 8318 -316
rect 8360 -440 8406 -309
rect 588 -486 7770 -452
rect -48 -614 -2 -498
rect 40 -618 86 -495
rect 588 -523 1596 -486
rect 6762 -528 7770 -486
rect 8259 -495 8269 -443
rect 8321 -495 8331 -443
rect 8360 -452 8555 -440
rect 8360 -486 8366 -452
rect 8400 -486 8515 -452
rect 8549 -486 8555 -452
rect 8272 -614 8318 -495
rect 8360 -498 8555 -486
rect 8360 -610 8406 -498
rect 2085 -792 2095 -616
rect 2147 -792 2157 -616
rect 4143 -792 4153 -616
rect 4205 -792 4215 -616
rect 6201 -792 6211 -616
rect 6263 -792 6273 -616
rect -152 -924 -142 -872
rect -90 -875 -80 -872
rect 8438 -875 8448 -872
rect -90 -921 8448 -875
rect -90 -924 -80 -921
rect 588 -962 1596 -921
rect 3639 -995 4736 -949
rect 6762 -954 7770 -921
rect 8438 -924 8448 -921
rect 8500 -924 8510 -872
rect -48 -1283 -2 -1203
rect 27 -1224 37 -1048
rect 89 -1224 99 -1048
rect 2085 -1224 2095 -1048
rect 2147 -1224 2157 -1048
rect 4156 -1050 4202 -995
rect -48 -1317 -42 -1283
rect -8 -1317 -2 -1283
rect -48 -1376 -2 -1317
rect -48 -1410 -42 -1376
rect -8 -1410 -2 -1376
rect -48 -1422 -2 -1410
rect 2098 -1376 2144 -1224
rect 2098 -1410 2104 -1376
rect 2138 -1410 2144 -1376
rect 2098 -1422 2144 -1410
rect 4156 -1376 4202 -1204
rect 6201 -1224 6211 -1048
rect 6263 -1224 6273 -1048
rect 8259 -1224 8269 -1048
rect 8321 -1224 8331 -1048
rect 4156 -1410 4162 -1376
rect 4196 -1410 4202 -1376
rect 4156 -1422 4202 -1410
rect 6214 -1376 6260 -1224
rect 6214 -1410 6220 -1376
rect 6254 -1410 6260 -1376
rect 6214 -1422 6260 -1410
rect 8360 -1283 8406 -1236
rect 8360 -1317 8366 -1283
rect 8400 -1317 8406 -1283
rect 8360 -1376 8406 -1317
rect 8360 -1410 8366 -1376
rect 8400 -1410 8406 -1376
rect 8360 -1422 8406 -1410
<< via1 >>
rect 37 110 89 286
rect 2095 110 2147 286
rect 6211 110 6263 286
rect 8269 110 8321 286
rect -142 -66 -90 -14
rect 8448 -66 8500 -14
rect 2095 -322 2147 -146
rect 4153 -322 4205 -146
rect 6211 -322 6263 -146
rect 37 -495 89 -443
rect 8269 -495 8321 -443
rect 2095 -792 2147 -616
rect 4153 -792 4205 -616
rect 6211 -792 6263 -616
rect -142 -924 -90 -872
rect 8448 -924 8500 -872
rect 37 -1224 89 -1048
rect 2095 -1224 2147 -1048
rect 6211 -1224 6263 -1048
rect 8269 -1224 8321 -1048
<< metal2 >>
rect 37 336 8321 388
rect 37 296 89 336
rect 8269 296 8321 336
rect 35 286 91 296
rect 35 100 91 110
rect 2095 286 2147 296
rect -142 -14 -90 -4
rect -142 -872 -90 -66
rect 2095 -146 2147 110
rect 6211 286 6263 296
rect 35 -441 91 -431
rect 35 -507 91 -497
rect -142 -934 -90 -924
rect 2095 -616 2147 -322
rect 35 -1048 91 -1038
rect 35 -1234 91 -1224
rect 2095 -1048 2147 -792
rect 4153 -146 4205 -136
rect 4153 -616 4205 -322
rect 4153 -802 4205 -792
rect 6211 -146 6263 110
rect 8267 286 8323 296
rect 8267 100 8323 110
rect 6211 -616 6263 -322
rect 8448 -14 8500 -4
rect 8267 -441 8323 -431
rect 8267 -507 8323 -497
rect 2095 -1234 2147 -1224
rect 6211 -1048 6263 -792
rect 8448 -872 8500 -66
rect 8448 -934 8500 -924
rect 6211 -1234 6263 -1224
rect 8267 -1048 8323 -1038
rect 8267 -1234 8323 -1224
rect 37 -1274 89 -1234
rect 8269 -1274 8321 -1234
rect 37 -1326 8321 -1274
<< via2 >>
rect 35 110 37 286
rect 37 110 89 286
rect 89 110 91 286
rect 35 -443 91 -441
rect 35 -495 37 -443
rect 37 -495 89 -443
rect 89 -495 91 -443
rect 35 -497 91 -495
rect 35 -1224 37 -1048
rect 37 -1224 89 -1048
rect 89 -1224 91 -1048
rect 8267 110 8269 286
rect 8269 110 8321 286
rect 8321 110 8323 286
rect 8267 -443 8323 -441
rect 8267 -495 8269 -443
rect 8269 -495 8321 -443
rect 8321 -495 8323 -443
rect 8267 -497 8323 -495
rect 8267 -1224 8269 -1048
rect 8269 -1224 8321 -1048
rect 8321 -1224 8323 -1048
<< metal3 >>
rect 25 286 101 291
rect 25 110 35 286
rect 91 110 101 286
rect 25 105 101 110
rect 8257 286 8333 291
rect 8257 110 8267 286
rect 8323 110 8333 286
rect 8257 105 8333 110
rect 33 -4 93 105
rect -142 -64 93 -4
rect 8265 -4 8325 105
rect 8265 -64 8500 -4
rect -142 -874 -82 -64
rect 25 -439 101 -436
rect 8257 -439 8333 -436
rect 25 -441 8333 -439
rect 25 -497 35 -441
rect 91 -497 8267 -441
rect 8323 -497 8333 -441
rect 25 -499 8333 -497
rect 25 -502 101 -499
rect 8257 -502 8333 -499
rect 8440 -874 8500 -64
rect -142 -934 93 -874
rect 33 -1043 93 -934
rect 8265 -934 8500 -874
rect 8265 -1043 8325 -934
rect 25 -1048 101 -1043
rect 25 -1224 35 -1048
rect 91 -1224 101 -1048
rect 25 -1229 101 -1224
rect 8257 -1048 8333 -1043
rect 8257 -1224 8267 -1048
rect 8323 -1224 8333 -1048
rect 8257 -1229 8333 -1224
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_0
timestamp 1717421032
transform 1 0 19 0 1 -704
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_1
timestamp 1717421032
transform 1 0 8339 0 1 -1136
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_2
timestamp 1717421032
transform 1 0 8339 0 1 -704
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_3
timestamp 1717421032
transform 1 0 8339 0 1 -234
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_4
timestamp 1717421032
transform 1 0 8339 0 1 198
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_5
timestamp 1717421032
transform 1 0 19 0 1 198
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_6
timestamp 1717421032
transform 1 0 19 0 1 -234
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_8
timestamp 1717421032
transform 1 0 19 0 1 -1136
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_8WJJP2  sky130_fd_pr__pfet_01v8_8WJJP2_0
timestamp 1717408091
transform 1 0 4179 0 1 -668
box -4181 -198 4181 164
use sky130_fd_pr__pfet_01v8_8WJJP2  sky130_fd_pr__pfet_01v8_8WJJP2_1
timestamp 1717408091
transform 1 0 4179 0 1 -1100
box -4181 -198 4181 164
use sky130_fd_pr__pfet_01v8_C2SJBD  sky130_fd_pr__pfet_01v8_C2SJBD_0
timestamp 1717408091
transform 1 0 4179 0 1 162
box -4181 -164 4181 198
use sky130_fd_pr__pfet_01v8_C2SJBD  sky130_fd_pr__pfet_01v8_C2SJBD_1
timestamp 1717408091
transform 1 0 4179 0 1 -270
box -4181 -164 4181 198
<< labels >>
flabel metal1 4175 418 4175 418 0 FreeSans 160 0 0 0 vdde
port 1 nsew
flabel metal2 8473 -217 8473 -217 0 FreeSans 160 0 0 0 G10
port 2 nsew
flabel metal1 8294 -385 8294 -385 0 FreeSans 160 0 0 0 D2
port 4 nsew
flabel metal1 6783 -505 6783 -505 0 FreeSans 160 0 0 0 G
port 6 nsew
flabel metal3 8274 8 8274 8 0 FreeSans 160 0 0 0 D10
port 7 nsew
flabel metal2 4175 -374 4175 -374 0 FreeSans 160 0 0 0 D1
port 9 nsew
<< end >>
