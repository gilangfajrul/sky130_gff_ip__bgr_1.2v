magic
tech sky130A
magscale 1 2
timestamp 1717356610
<< nwell >>
rect -3381 -198 3381 164
<< pmos >>
rect -3287 -136 -1687 64
rect -1629 -136 -29 64
rect 29 -136 1629 64
rect 1687 -136 3287 64
<< pdiff >>
rect -3345 52 -3287 64
rect -3345 -124 -3333 52
rect -3299 -124 -3287 52
rect -3345 -136 -3287 -124
rect -1687 52 -1629 64
rect -1687 -124 -1675 52
rect -1641 -124 -1629 52
rect -1687 -136 -1629 -124
rect -29 52 29 64
rect -29 -124 -17 52
rect 17 -124 29 52
rect -29 -136 29 -124
rect 1629 52 1687 64
rect 1629 -124 1641 52
rect 1675 -124 1687 52
rect 1629 -136 1687 -124
rect 3287 52 3345 64
rect 3287 -124 3299 52
rect 3333 -124 3345 52
rect 3287 -136 3345 -124
<< pdiffc >>
rect -3333 -124 -3299 52
rect -1675 -124 -1641 52
rect -17 -124 17 52
rect 1641 -124 1675 52
rect 3299 -124 3333 52
<< poly >>
rect -2895 145 -2079 161
rect -2895 128 -2879 145
rect -3287 111 -2879 128
rect -2095 128 -2079 145
rect -1237 145 -421 161
rect -1237 128 -1221 145
rect -2095 111 -1687 128
rect -3287 64 -1687 111
rect -1629 111 -1221 128
rect -437 128 -421 145
rect 421 145 1237 161
rect 421 128 437 145
rect -437 111 -29 128
rect -1629 64 -29 111
rect 29 111 437 128
rect 1221 128 1237 145
rect 2079 145 2895 161
rect 2079 128 2095 145
rect 1221 111 1629 128
rect 29 64 1629 111
rect 1687 111 2095 128
rect 2879 128 2895 145
rect 2879 111 3287 128
rect 1687 64 3287 111
rect -3287 -162 -1687 -136
rect -1629 -162 -29 -136
rect 29 -162 1629 -136
rect 1687 -162 3287 -136
<< polycont >>
rect -2879 111 -2095 145
rect -1221 111 -437 145
rect 437 111 1221 145
rect 2095 111 2879 145
<< locali >>
rect -2895 111 -2879 145
rect -2095 111 -2079 145
rect -1237 111 -1221 145
rect -437 111 -421 145
rect 421 111 437 145
rect 1221 111 1237 145
rect 2079 111 2095 145
rect 2879 111 2895 145
rect -3333 52 -3299 68
rect -3333 -140 -3299 -124
rect -1675 52 -1641 68
rect -1675 -140 -1641 -124
rect -17 52 17 68
rect -17 -140 17 -124
rect 1641 52 1675 68
rect 1641 -140 1675 -124
rect 3299 52 3333 68
rect 3299 -140 3333 -124
<< viali >>
rect -2879 111 -2095 145
rect -1221 111 -437 145
rect 437 111 1221 145
rect 2095 111 2879 145
rect -3333 -124 -3299 52
rect -1675 -124 -1641 52
rect -17 -124 17 52
rect 1641 -124 1675 52
rect 3299 -124 3333 52
<< metal1 >>
rect -2891 145 -2083 151
rect -2891 111 -2879 145
rect -2095 111 -2083 145
rect -2891 105 -2083 111
rect -1233 145 -425 151
rect -1233 111 -1221 145
rect -437 111 -425 145
rect -1233 105 -425 111
rect 425 145 1233 151
rect 425 111 437 145
rect 1221 111 1233 145
rect 425 105 1233 111
rect 2083 145 2891 151
rect 2083 111 2095 145
rect 2879 111 2891 145
rect 2083 105 2891 111
rect -3339 52 -3293 64
rect -3339 -124 -3333 52
rect -3299 -124 -3293 52
rect -3339 -136 -3293 -124
rect -1681 52 -1635 64
rect -1681 -124 -1675 52
rect -1641 -124 -1635 52
rect -1681 -136 -1635 -124
rect -23 52 23 64
rect -23 -124 -17 52
rect 17 -124 23 52
rect -23 -136 23 -124
rect 1635 52 1681 64
rect 1635 -124 1641 52
rect 1675 -124 1681 52
rect 1635 -136 1681 -124
rect 3293 52 3339 64
rect 3293 -124 3299 52
rect 3333 -124 3339 52
rect 3293 -136 3339 -124
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 8 m 1 nf 4 diffcov 100 polycov 50 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
