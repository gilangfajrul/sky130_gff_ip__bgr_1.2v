magic
tech sky130A
magscale 1 2
timestamp 1716999520
<< pwell >>
rect -425 -519 425 519
<< nmos >>
rect -229 109 -29 309
rect 29 109 229 309
rect -229 -309 -29 -109
rect 29 -309 229 -109
<< ndiff >>
rect -287 297 -229 309
rect -287 121 -275 297
rect -241 121 -229 297
rect -287 109 -229 121
rect -29 297 29 309
rect -29 121 -17 297
rect 17 121 29 297
rect -29 109 29 121
rect 229 297 287 309
rect 229 121 241 297
rect 275 121 287 297
rect 229 109 287 121
rect -287 -121 -229 -109
rect -287 -297 -275 -121
rect -241 -297 -229 -121
rect -287 -309 -229 -297
rect -29 -121 29 -109
rect -29 -297 -17 -121
rect 17 -297 29 -121
rect -29 -309 29 -297
rect 229 -121 287 -109
rect 229 -297 241 -121
rect 275 -297 287 -121
rect 229 -309 287 -297
<< ndiffc >>
rect -275 121 -241 297
rect -17 121 17 297
rect 241 121 275 297
rect -275 -297 -241 -121
rect -17 -297 17 -121
rect 241 -297 275 -121
<< psubdiff >>
rect -389 449 -293 483
rect 293 449 389 483
rect -389 387 -355 449
rect 355 387 389 449
rect -389 -449 -355 -387
rect 355 -449 389 -387
rect -389 -483 -293 -449
rect 293 -483 389 -449
<< psubdiffcont >>
rect -293 449 293 483
rect -389 -387 -355 387
rect 355 -387 389 387
rect -293 -483 293 -449
<< poly >>
rect -229 381 -29 397
rect -229 347 -213 381
rect -45 347 -29 381
rect -229 309 -29 347
rect 29 381 229 397
rect 29 347 45 381
rect 213 347 229 381
rect 29 309 229 347
rect -229 71 -29 109
rect -229 37 -213 71
rect -45 37 -29 71
rect -229 21 -29 37
rect 29 71 229 109
rect 29 37 45 71
rect 213 37 229 71
rect 29 21 229 37
rect -229 -37 -29 -21
rect -229 -71 -213 -37
rect -45 -71 -29 -37
rect -229 -109 -29 -71
rect 29 -37 229 -21
rect 29 -71 45 -37
rect 213 -71 229 -37
rect 29 -109 229 -71
rect -229 -347 -29 -309
rect -229 -381 -213 -347
rect -45 -381 -29 -347
rect -229 -397 -29 -381
rect 29 -347 229 -309
rect 29 -381 45 -347
rect 213 -381 229 -347
rect 29 -397 229 -381
<< polycont >>
rect -213 347 -45 381
rect 45 347 213 381
rect -213 37 -45 71
rect 45 37 213 71
rect -213 -71 -45 -37
rect 45 -71 213 -37
rect -213 -381 -45 -347
rect 45 -381 213 -347
<< locali >>
rect -389 449 -293 483
rect 293 449 389 483
rect -389 387 -355 449
rect 355 387 389 449
rect -229 347 -213 381
rect -45 347 -29 381
rect 29 347 45 381
rect 213 347 229 381
rect -275 297 -241 313
rect -275 105 -241 121
rect -17 297 17 313
rect -17 105 17 121
rect 241 297 275 313
rect 241 105 275 121
rect -229 37 -213 71
rect -45 37 -29 71
rect 29 37 45 71
rect 213 37 229 71
rect -229 -71 -213 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 213 -71 229 -37
rect -275 -121 -241 -105
rect -275 -313 -241 -297
rect -17 -121 17 -105
rect -17 -313 17 -297
rect 241 -121 275 -105
rect 241 -313 275 -297
rect -229 -381 -213 -347
rect -45 -381 -29 -347
rect 29 -381 45 -347
rect 213 -381 229 -347
rect -389 -449 -355 -387
rect 355 -449 389 -387
rect -389 -483 -293 -449
rect 293 -483 389 -449
<< viali >>
rect -213 347 -45 381
rect 45 347 213 381
rect -275 121 -241 297
rect -17 121 17 297
rect 241 121 275 297
rect -213 37 -45 71
rect 45 37 213 71
rect -213 -71 -45 -37
rect 45 -71 213 -37
rect -275 -297 -241 -121
rect -17 -297 17 -121
rect 241 -297 275 -121
rect -213 -381 -45 -347
rect 45 -381 213 -347
<< metal1 >>
rect -225 381 -33 387
rect -225 347 -213 381
rect -45 347 -33 381
rect -225 341 -33 347
rect 33 381 225 387
rect 33 347 45 381
rect 213 347 225 381
rect 33 341 225 347
rect -281 297 -235 309
rect -281 121 -275 297
rect -241 121 -235 297
rect -281 109 -235 121
rect -23 297 23 309
rect -23 121 -17 297
rect 17 121 23 297
rect -23 109 23 121
rect 235 297 281 309
rect 235 121 241 297
rect 275 121 281 297
rect 235 109 281 121
rect -225 71 -33 77
rect -225 37 -213 71
rect -45 37 -33 71
rect -225 31 -33 37
rect 33 71 225 77
rect 33 37 45 71
rect 213 37 225 71
rect 33 31 225 37
rect -225 -37 -33 -31
rect -225 -71 -213 -37
rect -45 -71 -33 -37
rect -225 -77 -33 -71
rect 33 -37 225 -31
rect 33 -71 45 -37
rect 213 -71 225 -37
rect 33 -77 225 -71
rect -281 -121 -235 -109
rect -281 -297 -275 -121
rect -241 -297 -235 -121
rect -281 -309 -235 -297
rect -23 -121 23 -109
rect -23 -297 -17 -121
rect 17 -297 23 -121
rect -23 -309 23 -297
rect 235 -121 281 -109
rect 235 -297 241 -121
rect 275 -297 281 -121
rect 235 -309 281 -297
rect -225 -347 -33 -341
rect -225 -381 -213 -347
rect -45 -381 -33 -347
rect -225 -387 -33 -381
rect 33 -347 225 -341
rect 33 -381 45 -347
rect 213 -381 225 -347
rect 33 -387 225 -381
<< properties >>
string FIXED_BBOX -372 -466 372 466
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 1 m 2 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
