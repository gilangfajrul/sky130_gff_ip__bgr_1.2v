magic
tech sky130A
magscale 1 2
timestamp 1716351939
<< xpolycontact >>
rect -284 1608 -214 2040
rect -284 1098 -214 1530
rect -118 1608 -48 2040
rect -118 1098 -48 1530
rect 48 1608 118 2040
rect 48 1098 118 1530
rect 214 1608 284 2040
rect 214 1098 284 1530
rect -284 562 -214 994
rect -284 52 -214 484
rect -118 562 -48 994
rect -118 52 -48 484
rect 48 562 118 994
rect 48 52 118 484
rect 214 562 284 994
rect 214 52 284 484
rect -284 -484 -214 -52
rect -284 -994 -214 -562
rect -118 -484 -48 -52
rect -118 -994 -48 -562
rect 48 -484 118 -52
rect 48 -994 118 -562
rect 214 -484 284 -52
rect 214 -994 284 -562
rect -284 -1530 -214 -1098
rect -284 -2040 -214 -1608
rect -118 -1530 -48 -1098
rect -118 -2040 -48 -1608
rect 48 -1530 118 -1098
rect 48 -2040 118 -1608
rect 214 -1530 284 -1098
rect 214 -2040 284 -1608
<< ppolyres >>
rect -284 1530 -214 1608
rect -118 1530 -48 1608
rect 48 1530 118 1608
rect 214 1530 284 1608
rect -284 484 -214 562
rect -118 484 -48 562
rect 48 484 118 562
rect 214 484 284 562
rect -284 -562 -214 -484
rect -118 -562 -48 -484
rect 48 -562 118 -484
rect 214 -562 284 -484
rect -284 -1608 -214 -1530
rect -118 -1608 -48 -1530
rect 48 -1608 118 -1530
rect 214 -1608 284 -1530
<< viali >>
rect -268 1625 -230 2022
rect -102 1625 -64 2022
rect 64 1625 102 2022
rect 230 1625 268 2022
rect -268 1116 -230 1513
rect -102 1116 -64 1513
rect 64 1116 102 1513
rect 230 1116 268 1513
rect -268 579 -230 976
rect -102 579 -64 976
rect 64 579 102 976
rect 230 579 268 976
rect -268 70 -230 467
rect -102 70 -64 467
rect 64 70 102 467
rect 230 70 268 467
rect -268 -467 -230 -70
rect -102 -467 -64 -70
rect 64 -467 102 -70
rect 230 -467 268 -70
rect -268 -976 -230 -579
rect -102 -976 -64 -579
rect 64 -976 102 -579
rect 230 -976 268 -579
rect -268 -1513 -230 -1116
rect -102 -1513 -64 -1116
rect 64 -1513 102 -1116
rect 230 -1513 268 -1116
rect -268 -2022 -230 -1625
rect -102 -2022 -64 -1625
rect 64 -2022 102 -1625
rect 230 -2022 268 -1625
<< metal1 >>
rect -274 2022 -224 2034
rect -274 1625 -268 2022
rect -230 1625 -224 2022
rect -274 1613 -224 1625
rect -108 2022 -58 2034
rect -108 1625 -102 2022
rect -64 1625 -58 2022
rect -108 1613 -58 1625
rect 58 2022 108 2034
rect 58 1625 64 2022
rect 102 1625 108 2022
rect 58 1613 108 1625
rect 224 2022 274 2034
rect 224 1625 230 2022
rect 268 1625 274 2022
rect 224 1613 274 1625
rect -274 1513 -224 1525
rect -274 1116 -268 1513
rect -230 1116 -224 1513
rect -274 1104 -224 1116
rect -108 1513 -58 1525
rect -108 1116 -102 1513
rect -64 1116 -58 1513
rect -108 1104 -58 1116
rect 58 1513 108 1525
rect 58 1116 64 1513
rect 102 1116 108 1513
rect 58 1104 108 1116
rect 224 1513 274 1525
rect 224 1116 230 1513
rect 268 1116 274 1513
rect 224 1104 274 1116
rect -274 976 -224 988
rect -274 579 -268 976
rect -230 579 -224 976
rect -274 567 -224 579
rect -108 976 -58 988
rect -108 579 -102 976
rect -64 579 -58 976
rect -108 567 -58 579
rect 58 976 108 988
rect 58 579 64 976
rect 102 579 108 976
rect 58 567 108 579
rect 224 976 274 988
rect 224 579 230 976
rect 268 579 274 976
rect 224 567 274 579
rect -274 467 -224 479
rect -274 70 -268 467
rect -230 70 -224 467
rect -274 58 -224 70
rect -108 467 -58 479
rect -108 70 -102 467
rect -64 70 -58 467
rect -108 58 -58 70
rect 58 467 108 479
rect 58 70 64 467
rect 102 70 108 467
rect 58 58 108 70
rect 224 467 274 479
rect 224 70 230 467
rect 268 70 274 467
rect 224 58 274 70
rect -274 -70 -224 -58
rect -274 -467 -268 -70
rect -230 -467 -224 -70
rect -274 -479 -224 -467
rect -108 -70 -58 -58
rect -108 -467 -102 -70
rect -64 -467 -58 -70
rect -108 -479 -58 -467
rect 58 -70 108 -58
rect 58 -467 64 -70
rect 102 -467 108 -70
rect 58 -479 108 -467
rect 224 -70 274 -58
rect 224 -467 230 -70
rect 268 -467 274 -70
rect 224 -479 274 -467
rect -274 -579 -224 -567
rect -274 -976 -268 -579
rect -230 -976 -224 -579
rect -274 -988 -224 -976
rect -108 -579 -58 -567
rect -108 -976 -102 -579
rect -64 -976 -58 -579
rect -108 -988 -58 -976
rect 58 -579 108 -567
rect 58 -976 64 -579
rect 102 -976 108 -579
rect 58 -988 108 -976
rect 224 -579 274 -567
rect 224 -976 230 -579
rect 268 -976 274 -579
rect 224 -988 274 -976
rect -274 -1116 -224 -1104
rect -274 -1513 -268 -1116
rect -230 -1513 -224 -1116
rect -274 -1525 -224 -1513
rect -108 -1116 -58 -1104
rect -108 -1513 -102 -1116
rect -64 -1513 -58 -1116
rect -108 -1525 -58 -1513
rect 58 -1116 108 -1104
rect 58 -1513 64 -1116
rect 102 -1513 108 -1116
rect 58 -1525 108 -1513
rect 224 -1116 274 -1104
rect 224 -1513 230 -1116
rect 268 -1513 274 -1116
rect 224 -1525 274 -1513
rect -274 -1625 -224 -1613
rect -274 -2022 -268 -1625
rect -230 -2022 -224 -1625
rect -274 -2034 -224 -2022
rect -108 -1625 -58 -1613
rect -108 -2022 -102 -1625
rect -64 -2022 -58 -1625
rect -108 -2034 -58 -2022
rect 58 -1625 108 -1613
rect 58 -2022 64 -1625
rect 102 -2022 108 -1625
rect 58 -2034 108 -2022
rect 224 -1625 274 -1613
rect 224 -2022 230 -1625
rect 268 -2022 274 -1625
rect 224 -2034 274 -2022
<< properties >>
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.350 l 0.55 m 4 nx 4 wmin 0.350 lmin 0.50 rho 319.8 val 1.615k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
