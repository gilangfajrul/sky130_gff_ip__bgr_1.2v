** sch_path: /foss/designs/sky130_gff_ip__bgr_1.2v/xschem/op_tb.sch
**.subckt op_tb
V1 Vvdd GND 1.8
V2 vp GND 0.67
V3 vn GND ac 1 sin(0.671 1) dc 0.67
x1 out Vvdd Vgnd vp vn Vgnd Vvdd op
V4 Vgnd GND 0
C1 out Vgnd 1p m=1
**** begin user architecture code
.lib /foss/pdks/sky130A/libs.tech/combined/sky130.lib.spice tt


.temp 27
.control
option sparse
save all
op
write ota-5t_tb-ac.raw
set appendwrite

ac dec 101 1k 100MEG
write ota-5t_tb-ac.raw
plot 20*log10(v_out)

meas ac dcgain MAX vmag(v_out) FROM=10 TO=10k
let f3db = dcgain/sqrt(2)
meas ac fbw WHEN vmag(v_out)=f3db FALL=1
let gainerror=(dcgain-1)/1
print dcgain
print fbw
print gainerror

noise v(v_out) Vin dec 101 1k 100MEG
print onoise_total

.endc


**** end user architecture code
**.ends

* expanding   symbol:  op.sym # of pins=7
** sym_path: /foss/designs/sky130_gff_ip__bgr_1.2v/xschem/op.sym
** sch_path: /foss/designs/sky130_gff_ip__bgr_1.2v/xschem/op.sch
.subckt op vo_out vdd vss vi_p vi_n psubs nwell
*.iopin vss
*.iopin vdd
*.opin vo_out
*.ipin vi_p
*.ipin vi_n
*.iopin psubs
*.iopin nwell
XM1a net3 vi_p net1 psubs sky130_fd_pr__nfet_01v8 L=5 W=1.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
**** begin user architecture code


.include ./sizing_opamp.spice


**** end user architecture code
XM2a net3 net3 vdd nwell sky130_fd_pr__pfet_01v8 L=5 W=2.5 nf=1 ad=0.725 as=0.725 pd=5.58 ps=5.58 nrd=0.116 nrs=0.116 sa=0 sb=0
+ sd=0 mult=1 m=1
XM0a net4 net4 vss psubs sky130_fd_pr__nfet_01v8 L=1.5 W=6 nf=1 ad=1.74 as=1.74 pd=12.58 ps=12.58 nrd=0.0483333333333333
+ nrs=0.0483333333333333 sa=0 sb=0 sd=0 mult=1 m=1
I0 vdd net4 20e-6
XM3 net1 net4 vss psubs sky130_fd_pr__nfet_01v8 L=5 W=1.5 nf=1 ad=0.435 as=0.435 pd=3.58 ps=3.58 nrd=0.193333333333333
+ nrs=0.193333333333333 sa=0 sb=0 sd=0 mult=1 m=1
XM7 vo_out net2 vdd nwell sky130_fd_pr__pfet_01v8 L=5 W=4.5 nf=1 ad=1.305 as=1.305 pd=9.58 ps=9.58 nrd=0.0644444444444444
+ nrs=0.0644444444444444 sa=0 sb=0 sd=0 mult=1 m=1
XM8 vo_out net4 vss psubs sky130_fd_pr__nfet_01v8 L=5 W=0.5 nf={nf3} ad='int(({nf3} + 1)/2) * 0.5 / {nf3} * 0.29' as='int(({nf3} + 2)/2) * 0.5 / {nf3} * 0.29'
+ pd='2*int(({nf3} + 1)/2) * (0.5 / {nf3} + 0.29)' ps='2*int(({nf3} + 2)/2) * (0.5 / {nf3} + 0.29)' nrd=0.58 nrs=0.58 sa=0 sb=0 sd=0
+ mult=1 m=1
XR1 vo_out net5 vss sky130_fd_pr__res_high_po_0p35 L=32 mult=1 m=1
XC1 net2 net5 sky130_fd_pr__cap_mim_m3_1 W=128 L=128 MF=1 m=1
XM4 net2 vi_n net1 psubs sky130_fd_pr__nfet_01v8 L=5 W=1.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 net2 net3 vdd nwell sky130_fd_pr__pfet_01v8 L=5 W=2.5 nf=1 ad=0.725 as=0.725 pd=5.58 ps=5.58 nrd=0.116 nrs=0.116 sa=0 sb=0
+ sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
