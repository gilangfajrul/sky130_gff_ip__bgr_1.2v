magic
tech sky130A
magscale 1 2
timestamp 1717437593
<< pwell >>
rect -948 -17458 948 17458
<< psubdiff >>
rect -912 17388 -816 17422
rect 816 17388 912 17422
rect -912 17326 -878 17388
rect 878 17326 912 17388
rect -912 -17388 -878 -17326
rect 878 -17388 912 -17326
rect -912 -17422 -816 -17388
rect 816 -17422 912 -17388
<< psubdiffcont >>
rect -816 17388 816 17422
rect -912 -17326 -878 17326
rect 878 -17326 912 17326
rect -816 -17422 816 -17388
<< xpolycontact >>
rect -782 16860 -712 17292
rect -782 13060 -712 13492
rect -616 16860 -546 17292
rect -616 13060 -546 13492
rect -450 16860 -380 17292
rect -450 13060 -380 13492
rect -284 16860 -214 17292
rect -284 13060 -214 13492
rect -118 16860 -48 17292
rect -118 13060 -48 13492
rect 48 16860 118 17292
rect 48 13060 118 13492
rect 214 16860 284 17292
rect 214 13060 284 13492
rect 380 16860 450 17292
rect 380 13060 450 13492
rect 546 16860 616 17292
rect 546 13060 616 13492
rect 712 16860 782 17292
rect 712 13060 782 13492
rect -782 12524 -712 12956
rect -782 8724 -712 9156
rect -616 12524 -546 12956
rect -616 8724 -546 9156
rect -450 12524 -380 12956
rect -450 8724 -380 9156
rect -284 12524 -214 12956
rect -284 8724 -214 9156
rect -118 12524 -48 12956
rect -118 8724 -48 9156
rect 48 12524 118 12956
rect 48 8724 118 9156
rect 214 12524 284 12956
rect 214 8724 284 9156
rect 380 12524 450 12956
rect 380 8724 450 9156
rect 546 12524 616 12956
rect 546 8724 616 9156
rect 712 12524 782 12956
rect 712 8724 782 9156
rect -782 8188 -712 8620
rect -782 4388 -712 4820
rect -616 8188 -546 8620
rect -616 4388 -546 4820
rect -450 8188 -380 8620
rect -450 4388 -380 4820
rect -284 8188 -214 8620
rect -284 4388 -214 4820
rect -118 8188 -48 8620
rect -118 4388 -48 4820
rect 48 8188 118 8620
rect 48 4388 118 4820
rect 214 8188 284 8620
rect 214 4388 284 4820
rect 380 8188 450 8620
rect 380 4388 450 4820
rect 546 8188 616 8620
rect 546 4388 616 4820
rect 712 8188 782 8620
rect 712 4388 782 4820
rect -782 3852 -712 4284
rect -782 52 -712 484
rect -616 3852 -546 4284
rect -616 52 -546 484
rect -450 3852 -380 4284
rect -450 52 -380 484
rect -284 3852 -214 4284
rect -284 52 -214 484
rect -118 3852 -48 4284
rect -118 52 -48 484
rect 48 3852 118 4284
rect 48 52 118 484
rect 214 3852 284 4284
rect 214 52 284 484
rect 380 3852 450 4284
rect 380 52 450 484
rect 546 3852 616 4284
rect 546 52 616 484
rect 712 3852 782 4284
rect 712 52 782 484
rect -782 -484 -712 -52
rect -782 -4284 -712 -3852
rect -616 -484 -546 -52
rect -616 -4284 -546 -3852
rect -450 -484 -380 -52
rect -450 -4284 -380 -3852
rect -284 -484 -214 -52
rect -284 -4284 -214 -3852
rect -118 -484 -48 -52
rect -118 -4284 -48 -3852
rect 48 -484 118 -52
rect 48 -4284 118 -3852
rect 214 -484 284 -52
rect 214 -4284 284 -3852
rect 380 -484 450 -52
rect 380 -4284 450 -3852
rect 546 -484 616 -52
rect 546 -4284 616 -3852
rect 712 -484 782 -52
rect 712 -4284 782 -3852
rect -782 -4820 -712 -4388
rect -782 -8620 -712 -8188
rect -616 -4820 -546 -4388
rect -616 -8620 -546 -8188
rect -450 -4820 -380 -4388
rect -450 -8620 -380 -8188
rect -284 -4820 -214 -4388
rect -284 -8620 -214 -8188
rect -118 -4820 -48 -4388
rect -118 -8620 -48 -8188
rect 48 -4820 118 -4388
rect 48 -8620 118 -8188
rect 214 -4820 284 -4388
rect 214 -8620 284 -8188
rect 380 -4820 450 -4388
rect 380 -8620 450 -8188
rect 546 -4820 616 -4388
rect 546 -8620 616 -8188
rect 712 -4820 782 -4388
rect 712 -8620 782 -8188
rect -782 -9156 -712 -8724
rect -782 -12956 -712 -12524
rect -616 -9156 -546 -8724
rect -616 -12956 -546 -12524
rect -450 -9156 -380 -8724
rect -450 -12956 -380 -12524
rect -284 -9156 -214 -8724
rect -284 -12956 -214 -12524
rect -118 -9156 -48 -8724
rect -118 -12956 -48 -12524
rect 48 -9156 118 -8724
rect 48 -12956 118 -12524
rect 214 -9156 284 -8724
rect 214 -12956 284 -12524
rect 380 -9156 450 -8724
rect 380 -12956 450 -12524
rect 546 -9156 616 -8724
rect 546 -12956 616 -12524
rect 712 -9156 782 -8724
rect 712 -12956 782 -12524
rect -782 -13492 -712 -13060
rect -782 -17292 -712 -16860
rect -616 -13492 -546 -13060
rect -616 -17292 -546 -16860
rect -450 -13492 -380 -13060
rect -450 -17292 -380 -16860
rect -284 -13492 -214 -13060
rect -284 -17292 -214 -16860
rect -118 -13492 -48 -13060
rect -118 -17292 -48 -16860
rect 48 -13492 118 -13060
rect 48 -17292 118 -16860
rect 214 -13492 284 -13060
rect 214 -17292 284 -16860
rect 380 -13492 450 -13060
rect 380 -17292 450 -16860
rect 546 -13492 616 -13060
rect 546 -17292 616 -16860
rect 712 -13492 782 -13060
rect 712 -17292 782 -16860
<< ppolyres >>
rect -782 13492 -712 16860
rect -616 13492 -546 16860
rect -450 13492 -380 16860
rect -284 13492 -214 16860
rect -118 13492 -48 16860
rect 48 13492 118 16860
rect 214 13492 284 16860
rect 380 13492 450 16860
rect 546 13492 616 16860
rect 712 13492 782 16860
rect -782 9156 -712 12524
rect -616 9156 -546 12524
rect -450 9156 -380 12524
rect -284 9156 -214 12524
rect -118 9156 -48 12524
rect 48 9156 118 12524
rect 214 9156 284 12524
rect 380 9156 450 12524
rect 546 9156 616 12524
rect 712 9156 782 12524
rect -782 4820 -712 8188
rect -616 4820 -546 8188
rect -450 4820 -380 8188
rect -284 4820 -214 8188
rect -118 4820 -48 8188
rect 48 4820 118 8188
rect 214 4820 284 8188
rect 380 4820 450 8188
rect 546 4820 616 8188
rect 712 4820 782 8188
rect -782 484 -712 3852
rect -616 484 -546 3852
rect -450 484 -380 3852
rect -284 484 -214 3852
rect -118 484 -48 3852
rect 48 484 118 3852
rect 214 484 284 3852
rect 380 484 450 3852
rect 546 484 616 3852
rect 712 484 782 3852
rect -782 -3852 -712 -484
rect -616 -3852 -546 -484
rect -450 -3852 -380 -484
rect -284 -3852 -214 -484
rect -118 -3852 -48 -484
rect 48 -3852 118 -484
rect 214 -3852 284 -484
rect 380 -3852 450 -484
rect 546 -3852 616 -484
rect 712 -3852 782 -484
rect -782 -8188 -712 -4820
rect -616 -8188 -546 -4820
rect -450 -8188 -380 -4820
rect -284 -8188 -214 -4820
rect -118 -8188 -48 -4820
rect 48 -8188 118 -4820
rect 214 -8188 284 -4820
rect 380 -8188 450 -4820
rect 546 -8188 616 -4820
rect 712 -8188 782 -4820
rect -782 -12524 -712 -9156
rect -616 -12524 -546 -9156
rect -450 -12524 -380 -9156
rect -284 -12524 -214 -9156
rect -118 -12524 -48 -9156
rect 48 -12524 118 -9156
rect 214 -12524 284 -9156
rect 380 -12524 450 -9156
rect 546 -12524 616 -9156
rect 712 -12524 782 -9156
rect -782 -16860 -712 -13492
rect -616 -16860 -546 -13492
rect -450 -16860 -380 -13492
rect -284 -16860 -214 -13492
rect -118 -16860 -48 -13492
rect 48 -16860 118 -13492
rect 214 -16860 284 -13492
rect 380 -16860 450 -13492
rect 546 -16860 616 -13492
rect 712 -16860 782 -13492
<< locali >>
rect -912 17388 -816 17422
rect 816 17388 912 17422
rect -912 17326 -878 17388
rect 878 17326 912 17388
rect -912 -17388 -878 -17326
rect 878 -17388 912 -17326
rect -912 -17422 -816 -17388
rect 816 -17422 912 -17388
<< viali >>
rect -766 16877 -728 17274
rect -600 16877 -562 17274
rect -434 16877 -396 17274
rect -268 16877 -230 17274
rect -102 16877 -64 17274
rect 64 16877 102 17274
rect 230 16877 268 17274
rect 396 16877 434 17274
rect 562 16877 600 17274
rect 728 16877 766 17274
rect -766 13078 -728 13475
rect -600 13078 -562 13475
rect -434 13078 -396 13475
rect -268 13078 -230 13475
rect -102 13078 -64 13475
rect 64 13078 102 13475
rect 230 13078 268 13475
rect 396 13078 434 13475
rect 562 13078 600 13475
rect 728 13078 766 13475
rect -766 12541 -728 12938
rect -600 12541 -562 12938
rect -434 12541 -396 12938
rect -268 12541 -230 12938
rect -102 12541 -64 12938
rect 64 12541 102 12938
rect 230 12541 268 12938
rect 396 12541 434 12938
rect 562 12541 600 12938
rect 728 12541 766 12938
rect -766 8742 -728 9139
rect -600 8742 -562 9139
rect -434 8742 -396 9139
rect -268 8742 -230 9139
rect -102 8742 -64 9139
rect 64 8742 102 9139
rect 230 8742 268 9139
rect 396 8742 434 9139
rect 562 8742 600 9139
rect 728 8742 766 9139
rect -766 8205 -728 8602
rect -600 8205 -562 8602
rect -434 8205 -396 8602
rect -268 8205 -230 8602
rect -102 8205 -64 8602
rect 64 8205 102 8602
rect 230 8205 268 8602
rect 396 8205 434 8602
rect 562 8205 600 8602
rect 728 8205 766 8602
rect -766 4406 -728 4803
rect -600 4406 -562 4803
rect -434 4406 -396 4803
rect -268 4406 -230 4803
rect -102 4406 -64 4803
rect 64 4406 102 4803
rect 230 4406 268 4803
rect 396 4406 434 4803
rect 562 4406 600 4803
rect 728 4406 766 4803
rect -766 3869 -728 4266
rect -600 3869 -562 4266
rect -434 3869 -396 4266
rect -268 3869 -230 4266
rect -102 3869 -64 4266
rect 64 3869 102 4266
rect 230 3869 268 4266
rect 396 3869 434 4266
rect 562 3869 600 4266
rect 728 3869 766 4266
rect -766 70 -728 467
rect -600 70 -562 467
rect -434 70 -396 467
rect -268 70 -230 467
rect -102 70 -64 467
rect 64 70 102 467
rect 230 70 268 467
rect 396 70 434 467
rect 562 70 600 467
rect 728 70 766 467
rect -766 -467 -728 -70
rect -600 -467 -562 -70
rect -434 -467 -396 -70
rect -268 -467 -230 -70
rect -102 -467 -64 -70
rect 64 -467 102 -70
rect 230 -467 268 -70
rect 396 -467 434 -70
rect 562 -467 600 -70
rect 728 -467 766 -70
rect -766 -4266 -728 -3869
rect -600 -4266 -562 -3869
rect -434 -4266 -396 -3869
rect -268 -4266 -230 -3869
rect -102 -4266 -64 -3869
rect 64 -4266 102 -3869
rect 230 -4266 268 -3869
rect 396 -4266 434 -3869
rect 562 -4266 600 -3869
rect 728 -4266 766 -3869
rect -766 -4803 -728 -4406
rect -600 -4803 -562 -4406
rect -434 -4803 -396 -4406
rect -268 -4803 -230 -4406
rect -102 -4803 -64 -4406
rect 64 -4803 102 -4406
rect 230 -4803 268 -4406
rect 396 -4803 434 -4406
rect 562 -4803 600 -4406
rect 728 -4803 766 -4406
rect -766 -8602 -728 -8205
rect -600 -8602 -562 -8205
rect -434 -8602 -396 -8205
rect -268 -8602 -230 -8205
rect -102 -8602 -64 -8205
rect 64 -8602 102 -8205
rect 230 -8602 268 -8205
rect 396 -8602 434 -8205
rect 562 -8602 600 -8205
rect 728 -8602 766 -8205
rect -766 -9139 -728 -8742
rect -600 -9139 -562 -8742
rect -434 -9139 -396 -8742
rect -268 -9139 -230 -8742
rect -102 -9139 -64 -8742
rect 64 -9139 102 -8742
rect 230 -9139 268 -8742
rect 396 -9139 434 -8742
rect 562 -9139 600 -8742
rect 728 -9139 766 -8742
rect -766 -12938 -728 -12541
rect -600 -12938 -562 -12541
rect -434 -12938 -396 -12541
rect -268 -12938 -230 -12541
rect -102 -12938 -64 -12541
rect 64 -12938 102 -12541
rect 230 -12938 268 -12541
rect 396 -12938 434 -12541
rect 562 -12938 600 -12541
rect 728 -12938 766 -12541
rect -766 -13475 -728 -13078
rect -600 -13475 -562 -13078
rect -434 -13475 -396 -13078
rect -268 -13475 -230 -13078
rect -102 -13475 -64 -13078
rect 64 -13475 102 -13078
rect 230 -13475 268 -13078
rect 396 -13475 434 -13078
rect 562 -13475 600 -13078
rect 728 -13475 766 -13078
rect -766 -17274 -728 -16877
rect -600 -17274 -562 -16877
rect -434 -17274 -396 -16877
rect -268 -17274 -230 -16877
rect -102 -17274 -64 -16877
rect 64 -17274 102 -16877
rect 230 -17274 268 -16877
rect 396 -17274 434 -16877
rect 562 -17274 600 -16877
rect 728 -17274 766 -16877
<< metal1 >>
rect -772 17274 -722 17286
rect -772 16877 -766 17274
rect -728 16877 -722 17274
rect -772 16865 -722 16877
rect -606 17274 -556 17286
rect -606 16877 -600 17274
rect -562 16877 -556 17274
rect -606 16865 -556 16877
rect -440 17274 -390 17286
rect -440 16877 -434 17274
rect -396 16877 -390 17274
rect -440 16865 -390 16877
rect -274 17274 -224 17286
rect -274 16877 -268 17274
rect -230 16877 -224 17274
rect -274 16865 -224 16877
rect -108 17274 -58 17286
rect -108 16877 -102 17274
rect -64 16877 -58 17274
rect -108 16865 -58 16877
rect 58 17274 108 17286
rect 58 16877 64 17274
rect 102 16877 108 17274
rect 58 16865 108 16877
rect 224 17274 274 17286
rect 224 16877 230 17274
rect 268 16877 274 17274
rect 224 16865 274 16877
rect 390 17274 440 17286
rect 390 16877 396 17274
rect 434 16877 440 17274
rect 390 16865 440 16877
rect 556 17274 606 17286
rect 556 16877 562 17274
rect 600 16877 606 17274
rect 556 16865 606 16877
rect 722 17274 772 17286
rect 722 16877 728 17274
rect 766 16877 772 17274
rect 722 16865 772 16877
rect -772 13475 -722 13487
rect -772 13078 -766 13475
rect -728 13078 -722 13475
rect -772 13066 -722 13078
rect -606 13475 -556 13487
rect -606 13078 -600 13475
rect -562 13078 -556 13475
rect -606 13066 -556 13078
rect -440 13475 -390 13487
rect -440 13078 -434 13475
rect -396 13078 -390 13475
rect -440 13066 -390 13078
rect -274 13475 -224 13487
rect -274 13078 -268 13475
rect -230 13078 -224 13475
rect -274 13066 -224 13078
rect -108 13475 -58 13487
rect -108 13078 -102 13475
rect -64 13078 -58 13475
rect -108 13066 -58 13078
rect 58 13475 108 13487
rect 58 13078 64 13475
rect 102 13078 108 13475
rect 58 13066 108 13078
rect 224 13475 274 13487
rect 224 13078 230 13475
rect 268 13078 274 13475
rect 224 13066 274 13078
rect 390 13475 440 13487
rect 390 13078 396 13475
rect 434 13078 440 13475
rect 390 13066 440 13078
rect 556 13475 606 13487
rect 556 13078 562 13475
rect 600 13078 606 13475
rect 556 13066 606 13078
rect 722 13475 772 13487
rect 722 13078 728 13475
rect 766 13078 772 13475
rect 722 13066 772 13078
rect -772 12938 -722 12950
rect -772 12541 -766 12938
rect -728 12541 -722 12938
rect -772 12529 -722 12541
rect -606 12938 -556 12950
rect -606 12541 -600 12938
rect -562 12541 -556 12938
rect -606 12529 -556 12541
rect -440 12938 -390 12950
rect -440 12541 -434 12938
rect -396 12541 -390 12938
rect -440 12529 -390 12541
rect -274 12938 -224 12950
rect -274 12541 -268 12938
rect -230 12541 -224 12938
rect -274 12529 -224 12541
rect -108 12938 -58 12950
rect -108 12541 -102 12938
rect -64 12541 -58 12938
rect -108 12529 -58 12541
rect 58 12938 108 12950
rect 58 12541 64 12938
rect 102 12541 108 12938
rect 58 12529 108 12541
rect 224 12938 274 12950
rect 224 12541 230 12938
rect 268 12541 274 12938
rect 224 12529 274 12541
rect 390 12938 440 12950
rect 390 12541 396 12938
rect 434 12541 440 12938
rect 390 12529 440 12541
rect 556 12938 606 12950
rect 556 12541 562 12938
rect 600 12541 606 12938
rect 556 12529 606 12541
rect 722 12938 772 12950
rect 722 12541 728 12938
rect 766 12541 772 12938
rect 722 12529 772 12541
rect -772 9139 -722 9151
rect -772 8742 -766 9139
rect -728 8742 -722 9139
rect -772 8730 -722 8742
rect -606 9139 -556 9151
rect -606 8742 -600 9139
rect -562 8742 -556 9139
rect -606 8730 -556 8742
rect -440 9139 -390 9151
rect -440 8742 -434 9139
rect -396 8742 -390 9139
rect -440 8730 -390 8742
rect -274 9139 -224 9151
rect -274 8742 -268 9139
rect -230 8742 -224 9139
rect -274 8730 -224 8742
rect -108 9139 -58 9151
rect -108 8742 -102 9139
rect -64 8742 -58 9139
rect -108 8730 -58 8742
rect 58 9139 108 9151
rect 58 8742 64 9139
rect 102 8742 108 9139
rect 58 8730 108 8742
rect 224 9139 274 9151
rect 224 8742 230 9139
rect 268 8742 274 9139
rect 224 8730 274 8742
rect 390 9139 440 9151
rect 390 8742 396 9139
rect 434 8742 440 9139
rect 390 8730 440 8742
rect 556 9139 606 9151
rect 556 8742 562 9139
rect 600 8742 606 9139
rect 556 8730 606 8742
rect 722 9139 772 9151
rect 722 8742 728 9139
rect 766 8742 772 9139
rect 722 8730 772 8742
rect -772 8602 -722 8614
rect -772 8205 -766 8602
rect -728 8205 -722 8602
rect -772 8193 -722 8205
rect -606 8602 -556 8614
rect -606 8205 -600 8602
rect -562 8205 -556 8602
rect -606 8193 -556 8205
rect -440 8602 -390 8614
rect -440 8205 -434 8602
rect -396 8205 -390 8602
rect -440 8193 -390 8205
rect -274 8602 -224 8614
rect -274 8205 -268 8602
rect -230 8205 -224 8602
rect -274 8193 -224 8205
rect -108 8602 -58 8614
rect -108 8205 -102 8602
rect -64 8205 -58 8602
rect -108 8193 -58 8205
rect 58 8602 108 8614
rect 58 8205 64 8602
rect 102 8205 108 8602
rect 58 8193 108 8205
rect 224 8602 274 8614
rect 224 8205 230 8602
rect 268 8205 274 8602
rect 224 8193 274 8205
rect 390 8602 440 8614
rect 390 8205 396 8602
rect 434 8205 440 8602
rect 390 8193 440 8205
rect 556 8602 606 8614
rect 556 8205 562 8602
rect 600 8205 606 8602
rect 556 8193 606 8205
rect 722 8602 772 8614
rect 722 8205 728 8602
rect 766 8205 772 8602
rect 722 8193 772 8205
rect -772 4803 -722 4815
rect -772 4406 -766 4803
rect -728 4406 -722 4803
rect -772 4394 -722 4406
rect -606 4803 -556 4815
rect -606 4406 -600 4803
rect -562 4406 -556 4803
rect -606 4394 -556 4406
rect -440 4803 -390 4815
rect -440 4406 -434 4803
rect -396 4406 -390 4803
rect -440 4394 -390 4406
rect -274 4803 -224 4815
rect -274 4406 -268 4803
rect -230 4406 -224 4803
rect -274 4394 -224 4406
rect -108 4803 -58 4815
rect -108 4406 -102 4803
rect -64 4406 -58 4803
rect -108 4394 -58 4406
rect 58 4803 108 4815
rect 58 4406 64 4803
rect 102 4406 108 4803
rect 58 4394 108 4406
rect 224 4803 274 4815
rect 224 4406 230 4803
rect 268 4406 274 4803
rect 224 4394 274 4406
rect 390 4803 440 4815
rect 390 4406 396 4803
rect 434 4406 440 4803
rect 390 4394 440 4406
rect 556 4803 606 4815
rect 556 4406 562 4803
rect 600 4406 606 4803
rect 556 4394 606 4406
rect 722 4803 772 4815
rect 722 4406 728 4803
rect 766 4406 772 4803
rect 722 4394 772 4406
rect -772 4266 -722 4278
rect -772 3869 -766 4266
rect -728 3869 -722 4266
rect -772 3857 -722 3869
rect -606 4266 -556 4278
rect -606 3869 -600 4266
rect -562 3869 -556 4266
rect -606 3857 -556 3869
rect -440 4266 -390 4278
rect -440 3869 -434 4266
rect -396 3869 -390 4266
rect -440 3857 -390 3869
rect -274 4266 -224 4278
rect -274 3869 -268 4266
rect -230 3869 -224 4266
rect -274 3857 -224 3869
rect -108 4266 -58 4278
rect -108 3869 -102 4266
rect -64 3869 -58 4266
rect -108 3857 -58 3869
rect 58 4266 108 4278
rect 58 3869 64 4266
rect 102 3869 108 4266
rect 58 3857 108 3869
rect 224 4266 274 4278
rect 224 3869 230 4266
rect 268 3869 274 4266
rect 224 3857 274 3869
rect 390 4266 440 4278
rect 390 3869 396 4266
rect 434 3869 440 4266
rect 390 3857 440 3869
rect 556 4266 606 4278
rect 556 3869 562 4266
rect 600 3869 606 4266
rect 556 3857 606 3869
rect 722 4266 772 4278
rect 722 3869 728 4266
rect 766 3869 772 4266
rect 722 3857 772 3869
rect -772 467 -722 479
rect -772 70 -766 467
rect -728 70 -722 467
rect -772 58 -722 70
rect -606 467 -556 479
rect -606 70 -600 467
rect -562 70 -556 467
rect -606 58 -556 70
rect -440 467 -390 479
rect -440 70 -434 467
rect -396 70 -390 467
rect -440 58 -390 70
rect -274 467 -224 479
rect -274 70 -268 467
rect -230 70 -224 467
rect -274 58 -224 70
rect -108 467 -58 479
rect -108 70 -102 467
rect -64 70 -58 467
rect -108 58 -58 70
rect 58 467 108 479
rect 58 70 64 467
rect 102 70 108 467
rect 58 58 108 70
rect 224 467 274 479
rect 224 70 230 467
rect 268 70 274 467
rect 224 58 274 70
rect 390 467 440 479
rect 390 70 396 467
rect 434 70 440 467
rect 390 58 440 70
rect 556 467 606 479
rect 556 70 562 467
rect 600 70 606 467
rect 556 58 606 70
rect 722 467 772 479
rect 722 70 728 467
rect 766 70 772 467
rect 722 58 772 70
rect -772 -70 -722 -58
rect -772 -467 -766 -70
rect -728 -467 -722 -70
rect -772 -479 -722 -467
rect -606 -70 -556 -58
rect -606 -467 -600 -70
rect -562 -467 -556 -70
rect -606 -479 -556 -467
rect -440 -70 -390 -58
rect -440 -467 -434 -70
rect -396 -467 -390 -70
rect -440 -479 -390 -467
rect -274 -70 -224 -58
rect -274 -467 -268 -70
rect -230 -467 -224 -70
rect -274 -479 -224 -467
rect -108 -70 -58 -58
rect -108 -467 -102 -70
rect -64 -467 -58 -70
rect -108 -479 -58 -467
rect 58 -70 108 -58
rect 58 -467 64 -70
rect 102 -467 108 -70
rect 58 -479 108 -467
rect 224 -70 274 -58
rect 224 -467 230 -70
rect 268 -467 274 -70
rect 224 -479 274 -467
rect 390 -70 440 -58
rect 390 -467 396 -70
rect 434 -467 440 -70
rect 390 -479 440 -467
rect 556 -70 606 -58
rect 556 -467 562 -70
rect 600 -467 606 -70
rect 556 -479 606 -467
rect 722 -70 772 -58
rect 722 -467 728 -70
rect 766 -467 772 -70
rect 722 -479 772 -467
rect -772 -3869 -722 -3857
rect -772 -4266 -766 -3869
rect -728 -4266 -722 -3869
rect -772 -4278 -722 -4266
rect -606 -3869 -556 -3857
rect -606 -4266 -600 -3869
rect -562 -4266 -556 -3869
rect -606 -4278 -556 -4266
rect -440 -3869 -390 -3857
rect -440 -4266 -434 -3869
rect -396 -4266 -390 -3869
rect -440 -4278 -390 -4266
rect -274 -3869 -224 -3857
rect -274 -4266 -268 -3869
rect -230 -4266 -224 -3869
rect -274 -4278 -224 -4266
rect -108 -3869 -58 -3857
rect -108 -4266 -102 -3869
rect -64 -4266 -58 -3869
rect -108 -4278 -58 -4266
rect 58 -3869 108 -3857
rect 58 -4266 64 -3869
rect 102 -4266 108 -3869
rect 58 -4278 108 -4266
rect 224 -3869 274 -3857
rect 224 -4266 230 -3869
rect 268 -4266 274 -3869
rect 224 -4278 274 -4266
rect 390 -3869 440 -3857
rect 390 -4266 396 -3869
rect 434 -4266 440 -3869
rect 390 -4278 440 -4266
rect 556 -3869 606 -3857
rect 556 -4266 562 -3869
rect 600 -4266 606 -3869
rect 556 -4278 606 -4266
rect 722 -3869 772 -3857
rect 722 -4266 728 -3869
rect 766 -4266 772 -3869
rect 722 -4278 772 -4266
rect -772 -4406 -722 -4394
rect -772 -4803 -766 -4406
rect -728 -4803 -722 -4406
rect -772 -4815 -722 -4803
rect -606 -4406 -556 -4394
rect -606 -4803 -600 -4406
rect -562 -4803 -556 -4406
rect -606 -4815 -556 -4803
rect -440 -4406 -390 -4394
rect -440 -4803 -434 -4406
rect -396 -4803 -390 -4406
rect -440 -4815 -390 -4803
rect -274 -4406 -224 -4394
rect -274 -4803 -268 -4406
rect -230 -4803 -224 -4406
rect -274 -4815 -224 -4803
rect -108 -4406 -58 -4394
rect -108 -4803 -102 -4406
rect -64 -4803 -58 -4406
rect -108 -4815 -58 -4803
rect 58 -4406 108 -4394
rect 58 -4803 64 -4406
rect 102 -4803 108 -4406
rect 58 -4815 108 -4803
rect 224 -4406 274 -4394
rect 224 -4803 230 -4406
rect 268 -4803 274 -4406
rect 224 -4815 274 -4803
rect 390 -4406 440 -4394
rect 390 -4803 396 -4406
rect 434 -4803 440 -4406
rect 390 -4815 440 -4803
rect 556 -4406 606 -4394
rect 556 -4803 562 -4406
rect 600 -4803 606 -4406
rect 556 -4815 606 -4803
rect 722 -4406 772 -4394
rect 722 -4803 728 -4406
rect 766 -4803 772 -4406
rect 722 -4815 772 -4803
rect -772 -8205 -722 -8193
rect -772 -8602 -766 -8205
rect -728 -8602 -722 -8205
rect -772 -8614 -722 -8602
rect -606 -8205 -556 -8193
rect -606 -8602 -600 -8205
rect -562 -8602 -556 -8205
rect -606 -8614 -556 -8602
rect -440 -8205 -390 -8193
rect -440 -8602 -434 -8205
rect -396 -8602 -390 -8205
rect -440 -8614 -390 -8602
rect -274 -8205 -224 -8193
rect -274 -8602 -268 -8205
rect -230 -8602 -224 -8205
rect -274 -8614 -224 -8602
rect -108 -8205 -58 -8193
rect -108 -8602 -102 -8205
rect -64 -8602 -58 -8205
rect -108 -8614 -58 -8602
rect 58 -8205 108 -8193
rect 58 -8602 64 -8205
rect 102 -8602 108 -8205
rect 58 -8614 108 -8602
rect 224 -8205 274 -8193
rect 224 -8602 230 -8205
rect 268 -8602 274 -8205
rect 224 -8614 274 -8602
rect 390 -8205 440 -8193
rect 390 -8602 396 -8205
rect 434 -8602 440 -8205
rect 390 -8614 440 -8602
rect 556 -8205 606 -8193
rect 556 -8602 562 -8205
rect 600 -8602 606 -8205
rect 556 -8614 606 -8602
rect 722 -8205 772 -8193
rect 722 -8602 728 -8205
rect 766 -8602 772 -8205
rect 722 -8614 772 -8602
rect -772 -8742 -722 -8730
rect -772 -9139 -766 -8742
rect -728 -9139 -722 -8742
rect -772 -9151 -722 -9139
rect -606 -8742 -556 -8730
rect -606 -9139 -600 -8742
rect -562 -9139 -556 -8742
rect -606 -9151 -556 -9139
rect -440 -8742 -390 -8730
rect -440 -9139 -434 -8742
rect -396 -9139 -390 -8742
rect -440 -9151 -390 -9139
rect -274 -8742 -224 -8730
rect -274 -9139 -268 -8742
rect -230 -9139 -224 -8742
rect -274 -9151 -224 -9139
rect -108 -8742 -58 -8730
rect -108 -9139 -102 -8742
rect -64 -9139 -58 -8742
rect -108 -9151 -58 -9139
rect 58 -8742 108 -8730
rect 58 -9139 64 -8742
rect 102 -9139 108 -8742
rect 58 -9151 108 -9139
rect 224 -8742 274 -8730
rect 224 -9139 230 -8742
rect 268 -9139 274 -8742
rect 224 -9151 274 -9139
rect 390 -8742 440 -8730
rect 390 -9139 396 -8742
rect 434 -9139 440 -8742
rect 390 -9151 440 -9139
rect 556 -8742 606 -8730
rect 556 -9139 562 -8742
rect 600 -9139 606 -8742
rect 556 -9151 606 -9139
rect 722 -8742 772 -8730
rect 722 -9139 728 -8742
rect 766 -9139 772 -8742
rect 722 -9151 772 -9139
rect -772 -12541 -722 -12529
rect -772 -12938 -766 -12541
rect -728 -12938 -722 -12541
rect -772 -12950 -722 -12938
rect -606 -12541 -556 -12529
rect -606 -12938 -600 -12541
rect -562 -12938 -556 -12541
rect -606 -12950 -556 -12938
rect -440 -12541 -390 -12529
rect -440 -12938 -434 -12541
rect -396 -12938 -390 -12541
rect -440 -12950 -390 -12938
rect -274 -12541 -224 -12529
rect -274 -12938 -268 -12541
rect -230 -12938 -224 -12541
rect -274 -12950 -224 -12938
rect -108 -12541 -58 -12529
rect -108 -12938 -102 -12541
rect -64 -12938 -58 -12541
rect -108 -12950 -58 -12938
rect 58 -12541 108 -12529
rect 58 -12938 64 -12541
rect 102 -12938 108 -12541
rect 58 -12950 108 -12938
rect 224 -12541 274 -12529
rect 224 -12938 230 -12541
rect 268 -12938 274 -12541
rect 224 -12950 274 -12938
rect 390 -12541 440 -12529
rect 390 -12938 396 -12541
rect 434 -12938 440 -12541
rect 390 -12950 440 -12938
rect 556 -12541 606 -12529
rect 556 -12938 562 -12541
rect 600 -12938 606 -12541
rect 556 -12950 606 -12938
rect 722 -12541 772 -12529
rect 722 -12938 728 -12541
rect 766 -12938 772 -12541
rect 722 -12950 772 -12938
rect -772 -13078 -722 -13066
rect -772 -13475 -766 -13078
rect -728 -13475 -722 -13078
rect -772 -13487 -722 -13475
rect -606 -13078 -556 -13066
rect -606 -13475 -600 -13078
rect -562 -13475 -556 -13078
rect -606 -13487 -556 -13475
rect -440 -13078 -390 -13066
rect -440 -13475 -434 -13078
rect -396 -13475 -390 -13078
rect -440 -13487 -390 -13475
rect -274 -13078 -224 -13066
rect -274 -13475 -268 -13078
rect -230 -13475 -224 -13078
rect -274 -13487 -224 -13475
rect -108 -13078 -58 -13066
rect -108 -13475 -102 -13078
rect -64 -13475 -58 -13078
rect -108 -13487 -58 -13475
rect 58 -13078 108 -13066
rect 58 -13475 64 -13078
rect 102 -13475 108 -13078
rect 58 -13487 108 -13475
rect 224 -13078 274 -13066
rect 224 -13475 230 -13078
rect 268 -13475 274 -13078
rect 224 -13487 274 -13475
rect 390 -13078 440 -13066
rect 390 -13475 396 -13078
rect 434 -13475 440 -13078
rect 390 -13487 440 -13475
rect 556 -13078 606 -13066
rect 556 -13475 562 -13078
rect 600 -13475 606 -13078
rect 556 -13487 606 -13475
rect 722 -13078 772 -13066
rect 722 -13475 728 -13078
rect 766 -13475 772 -13078
rect 722 -13487 772 -13475
rect -772 -16877 -722 -16865
rect -772 -17274 -766 -16877
rect -728 -17274 -722 -16877
rect -772 -17286 -722 -17274
rect -606 -16877 -556 -16865
rect -606 -17274 -600 -16877
rect -562 -17274 -556 -16877
rect -606 -17286 -556 -17274
rect -440 -16877 -390 -16865
rect -440 -17274 -434 -16877
rect -396 -17274 -390 -16877
rect -440 -17286 -390 -17274
rect -274 -16877 -224 -16865
rect -274 -17274 -268 -16877
rect -230 -17274 -224 -16877
rect -274 -17286 -224 -17274
rect -108 -16877 -58 -16865
rect -108 -17274 -102 -16877
rect -64 -17274 -58 -16877
rect -108 -17286 -58 -17274
rect 58 -16877 108 -16865
rect 58 -17274 64 -16877
rect 102 -17274 108 -16877
rect 58 -17286 108 -17274
rect 224 -16877 274 -16865
rect 224 -17274 230 -16877
rect 268 -17274 274 -16877
rect 224 -17286 274 -17274
rect 390 -16877 440 -16865
rect 390 -17274 396 -16877
rect 434 -17274 440 -16877
rect 390 -17286 440 -17274
rect 556 -16877 606 -16865
rect 556 -17274 562 -16877
rect 600 -17274 606 -16877
rect 556 -17286 606 -17274
rect 722 -16877 772 -16865
rect 722 -17274 728 -16877
rect 766 -17274 772 -16877
rect 722 -17286 772 -17274
<< properties >>
string FIXED_BBOX -895 -17405 895 17405
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.350 l 17 m 8 nx 10 wmin 0.350 lmin 0.50 rho 319.8 val 16.646k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
