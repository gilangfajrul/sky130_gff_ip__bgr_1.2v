magic
tech sky130A
magscale 1 2
timestamp 1717437593
<< pwell >>
rect -616 -26130 616 26130
<< psubdiff >>
rect -580 26060 -484 26094
rect 484 26060 580 26094
rect -580 25998 -546 26060
rect 546 25998 580 26060
rect -580 -26060 -546 -25998
rect 546 -26060 580 -25998
rect -580 -26094 -484 -26060
rect 484 -26094 580 -26060
<< psubdiffcont >>
rect -484 26060 484 26094
rect -580 -25998 -546 25998
rect 546 -25998 580 25998
rect -484 -26094 484 -26060
<< xpolycontact >>
rect -450 25532 -380 25964
rect -450 21732 -380 22164
rect -284 25532 -214 25964
rect -284 21732 -214 22164
rect -118 25532 -48 25964
rect -118 21732 -48 22164
rect 48 25532 118 25964
rect 48 21732 118 22164
rect 214 25532 284 25964
rect 214 21732 284 22164
rect 380 25532 450 25964
rect 380 21732 450 22164
rect -450 21196 -380 21628
rect -450 17396 -380 17828
rect -284 21196 -214 21628
rect -284 17396 -214 17828
rect -118 21196 -48 21628
rect -118 17396 -48 17828
rect 48 21196 118 21628
rect 48 17396 118 17828
rect 214 21196 284 21628
rect 214 17396 284 17828
rect 380 21196 450 21628
rect 380 17396 450 17828
rect -450 16860 -380 17292
rect -450 13060 -380 13492
rect -284 16860 -214 17292
rect -284 13060 -214 13492
rect -118 16860 -48 17292
rect -118 13060 -48 13492
rect 48 16860 118 17292
rect 48 13060 118 13492
rect 214 16860 284 17292
rect 214 13060 284 13492
rect 380 16860 450 17292
rect 380 13060 450 13492
rect -450 12524 -380 12956
rect -450 8724 -380 9156
rect -284 12524 -214 12956
rect -284 8724 -214 9156
rect -118 12524 -48 12956
rect -118 8724 -48 9156
rect 48 12524 118 12956
rect 48 8724 118 9156
rect 214 12524 284 12956
rect 214 8724 284 9156
rect 380 12524 450 12956
rect 380 8724 450 9156
rect -450 8188 -380 8620
rect -450 4388 -380 4820
rect -284 8188 -214 8620
rect -284 4388 -214 4820
rect -118 8188 -48 8620
rect -118 4388 -48 4820
rect 48 8188 118 8620
rect 48 4388 118 4820
rect 214 8188 284 8620
rect 214 4388 284 4820
rect 380 8188 450 8620
rect 380 4388 450 4820
rect -450 3852 -380 4284
rect -450 52 -380 484
rect -284 3852 -214 4284
rect -284 52 -214 484
rect -118 3852 -48 4284
rect -118 52 -48 484
rect 48 3852 118 4284
rect 48 52 118 484
rect 214 3852 284 4284
rect 214 52 284 484
rect 380 3852 450 4284
rect 380 52 450 484
rect -450 -484 -380 -52
rect -450 -4284 -380 -3852
rect -284 -484 -214 -52
rect -284 -4284 -214 -3852
rect -118 -484 -48 -52
rect -118 -4284 -48 -3852
rect 48 -484 118 -52
rect 48 -4284 118 -3852
rect 214 -484 284 -52
rect 214 -4284 284 -3852
rect 380 -484 450 -52
rect 380 -4284 450 -3852
rect -450 -4820 -380 -4388
rect -450 -8620 -380 -8188
rect -284 -4820 -214 -4388
rect -284 -8620 -214 -8188
rect -118 -4820 -48 -4388
rect -118 -8620 -48 -8188
rect 48 -4820 118 -4388
rect 48 -8620 118 -8188
rect 214 -4820 284 -4388
rect 214 -8620 284 -8188
rect 380 -4820 450 -4388
rect 380 -8620 450 -8188
rect -450 -9156 -380 -8724
rect -450 -12956 -380 -12524
rect -284 -9156 -214 -8724
rect -284 -12956 -214 -12524
rect -118 -9156 -48 -8724
rect -118 -12956 -48 -12524
rect 48 -9156 118 -8724
rect 48 -12956 118 -12524
rect 214 -9156 284 -8724
rect 214 -12956 284 -12524
rect 380 -9156 450 -8724
rect 380 -12956 450 -12524
rect -450 -13492 -380 -13060
rect -450 -17292 -380 -16860
rect -284 -13492 -214 -13060
rect -284 -17292 -214 -16860
rect -118 -13492 -48 -13060
rect -118 -17292 -48 -16860
rect 48 -13492 118 -13060
rect 48 -17292 118 -16860
rect 214 -13492 284 -13060
rect 214 -17292 284 -16860
rect 380 -13492 450 -13060
rect 380 -17292 450 -16860
rect -450 -17828 -380 -17396
rect -450 -21628 -380 -21196
rect -284 -17828 -214 -17396
rect -284 -21628 -214 -21196
rect -118 -17828 -48 -17396
rect -118 -21628 -48 -21196
rect 48 -17828 118 -17396
rect 48 -21628 118 -21196
rect 214 -17828 284 -17396
rect 214 -21628 284 -21196
rect 380 -17828 450 -17396
rect 380 -21628 450 -21196
rect -450 -22164 -380 -21732
rect -450 -25964 -380 -25532
rect -284 -22164 -214 -21732
rect -284 -25964 -214 -25532
rect -118 -22164 -48 -21732
rect -118 -25964 -48 -25532
rect 48 -22164 118 -21732
rect 48 -25964 118 -25532
rect 214 -22164 284 -21732
rect 214 -25964 284 -25532
rect 380 -22164 450 -21732
rect 380 -25964 450 -25532
<< ppolyres >>
rect -450 22164 -380 25532
rect -284 22164 -214 25532
rect -118 22164 -48 25532
rect 48 22164 118 25532
rect 214 22164 284 25532
rect 380 22164 450 25532
rect -450 17828 -380 21196
rect -284 17828 -214 21196
rect -118 17828 -48 21196
rect 48 17828 118 21196
rect 214 17828 284 21196
rect 380 17828 450 21196
rect -450 13492 -380 16860
rect -284 13492 -214 16860
rect -118 13492 -48 16860
rect 48 13492 118 16860
rect 214 13492 284 16860
rect 380 13492 450 16860
rect -450 9156 -380 12524
rect -284 9156 -214 12524
rect -118 9156 -48 12524
rect 48 9156 118 12524
rect 214 9156 284 12524
rect 380 9156 450 12524
rect -450 4820 -380 8188
rect -284 4820 -214 8188
rect -118 4820 -48 8188
rect 48 4820 118 8188
rect 214 4820 284 8188
rect 380 4820 450 8188
rect -450 484 -380 3852
rect -284 484 -214 3852
rect -118 484 -48 3852
rect 48 484 118 3852
rect 214 484 284 3852
rect 380 484 450 3852
rect -450 -3852 -380 -484
rect -284 -3852 -214 -484
rect -118 -3852 -48 -484
rect 48 -3852 118 -484
rect 214 -3852 284 -484
rect 380 -3852 450 -484
rect -450 -8188 -380 -4820
rect -284 -8188 -214 -4820
rect -118 -8188 -48 -4820
rect 48 -8188 118 -4820
rect 214 -8188 284 -4820
rect 380 -8188 450 -4820
rect -450 -12524 -380 -9156
rect -284 -12524 -214 -9156
rect -118 -12524 -48 -9156
rect 48 -12524 118 -9156
rect 214 -12524 284 -9156
rect 380 -12524 450 -9156
rect -450 -16860 -380 -13492
rect -284 -16860 -214 -13492
rect -118 -16860 -48 -13492
rect 48 -16860 118 -13492
rect 214 -16860 284 -13492
rect 380 -16860 450 -13492
rect -450 -21196 -380 -17828
rect -284 -21196 -214 -17828
rect -118 -21196 -48 -17828
rect 48 -21196 118 -17828
rect 214 -21196 284 -17828
rect 380 -21196 450 -17828
rect -450 -25532 -380 -22164
rect -284 -25532 -214 -22164
rect -118 -25532 -48 -22164
rect 48 -25532 118 -22164
rect 214 -25532 284 -22164
rect 380 -25532 450 -22164
<< locali >>
rect -580 26060 -484 26094
rect 484 26060 580 26094
rect -580 25998 -546 26060
rect 546 25998 580 26060
rect -580 -26060 -546 -25998
rect 546 -26060 580 -25998
rect -580 -26094 -484 -26060
rect 484 -26094 580 -26060
<< viali >>
rect -434 25549 -396 25946
rect -268 25549 -230 25946
rect -102 25549 -64 25946
rect 64 25549 102 25946
rect 230 25549 268 25946
rect 396 25549 434 25946
rect -434 21750 -396 22147
rect -268 21750 -230 22147
rect -102 21750 -64 22147
rect 64 21750 102 22147
rect 230 21750 268 22147
rect 396 21750 434 22147
rect -434 21213 -396 21610
rect -268 21213 -230 21610
rect -102 21213 -64 21610
rect 64 21213 102 21610
rect 230 21213 268 21610
rect 396 21213 434 21610
rect -434 17414 -396 17811
rect -268 17414 -230 17811
rect -102 17414 -64 17811
rect 64 17414 102 17811
rect 230 17414 268 17811
rect 396 17414 434 17811
rect -434 16877 -396 17274
rect -268 16877 -230 17274
rect -102 16877 -64 17274
rect 64 16877 102 17274
rect 230 16877 268 17274
rect 396 16877 434 17274
rect -434 13078 -396 13475
rect -268 13078 -230 13475
rect -102 13078 -64 13475
rect 64 13078 102 13475
rect 230 13078 268 13475
rect 396 13078 434 13475
rect -434 12541 -396 12938
rect -268 12541 -230 12938
rect -102 12541 -64 12938
rect 64 12541 102 12938
rect 230 12541 268 12938
rect 396 12541 434 12938
rect -434 8742 -396 9139
rect -268 8742 -230 9139
rect -102 8742 -64 9139
rect 64 8742 102 9139
rect 230 8742 268 9139
rect 396 8742 434 9139
rect -434 8205 -396 8602
rect -268 8205 -230 8602
rect -102 8205 -64 8602
rect 64 8205 102 8602
rect 230 8205 268 8602
rect 396 8205 434 8602
rect -434 4406 -396 4803
rect -268 4406 -230 4803
rect -102 4406 -64 4803
rect 64 4406 102 4803
rect 230 4406 268 4803
rect 396 4406 434 4803
rect -434 3869 -396 4266
rect -268 3869 -230 4266
rect -102 3869 -64 4266
rect 64 3869 102 4266
rect 230 3869 268 4266
rect 396 3869 434 4266
rect -434 70 -396 467
rect -268 70 -230 467
rect -102 70 -64 467
rect 64 70 102 467
rect 230 70 268 467
rect 396 70 434 467
rect -434 -467 -396 -70
rect -268 -467 -230 -70
rect -102 -467 -64 -70
rect 64 -467 102 -70
rect 230 -467 268 -70
rect 396 -467 434 -70
rect -434 -4266 -396 -3869
rect -268 -4266 -230 -3869
rect -102 -4266 -64 -3869
rect 64 -4266 102 -3869
rect 230 -4266 268 -3869
rect 396 -4266 434 -3869
rect -434 -4803 -396 -4406
rect -268 -4803 -230 -4406
rect -102 -4803 -64 -4406
rect 64 -4803 102 -4406
rect 230 -4803 268 -4406
rect 396 -4803 434 -4406
rect -434 -8602 -396 -8205
rect -268 -8602 -230 -8205
rect -102 -8602 -64 -8205
rect 64 -8602 102 -8205
rect 230 -8602 268 -8205
rect 396 -8602 434 -8205
rect -434 -9139 -396 -8742
rect -268 -9139 -230 -8742
rect -102 -9139 -64 -8742
rect 64 -9139 102 -8742
rect 230 -9139 268 -8742
rect 396 -9139 434 -8742
rect -434 -12938 -396 -12541
rect -268 -12938 -230 -12541
rect -102 -12938 -64 -12541
rect 64 -12938 102 -12541
rect 230 -12938 268 -12541
rect 396 -12938 434 -12541
rect -434 -13475 -396 -13078
rect -268 -13475 -230 -13078
rect -102 -13475 -64 -13078
rect 64 -13475 102 -13078
rect 230 -13475 268 -13078
rect 396 -13475 434 -13078
rect -434 -17274 -396 -16877
rect -268 -17274 -230 -16877
rect -102 -17274 -64 -16877
rect 64 -17274 102 -16877
rect 230 -17274 268 -16877
rect 396 -17274 434 -16877
rect -434 -17811 -396 -17414
rect -268 -17811 -230 -17414
rect -102 -17811 -64 -17414
rect 64 -17811 102 -17414
rect 230 -17811 268 -17414
rect 396 -17811 434 -17414
rect -434 -21610 -396 -21213
rect -268 -21610 -230 -21213
rect -102 -21610 -64 -21213
rect 64 -21610 102 -21213
rect 230 -21610 268 -21213
rect 396 -21610 434 -21213
rect -434 -22147 -396 -21750
rect -268 -22147 -230 -21750
rect -102 -22147 -64 -21750
rect 64 -22147 102 -21750
rect 230 -22147 268 -21750
rect 396 -22147 434 -21750
rect -434 -25946 -396 -25549
rect -268 -25946 -230 -25549
rect -102 -25946 -64 -25549
rect 64 -25946 102 -25549
rect 230 -25946 268 -25549
rect 396 -25946 434 -25549
<< metal1 >>
rect -440 25946 -390 25958
rect -440 25549 -434 25946
rect -396 25549 -390 25946
rect -440 25537 -390 25549
rect -274 25946 -224 25958
rect -274 25549 -268 25946
rect -230 25549 -224 25946
rect -274 25537 -224 25549
rect -108 25946 -58 25958
rect -108 25549 -102 25946
rect -64 25549 -58 25946
rect -108 25537 -58 25549
rect 58 25946 108 25958
rect 58 25549 64 25946
rect 102 25549 108 25946
rect 58 25537 108 25549
rect 224 25946 274 25958
rect 224 25549 230 25946
rect 268 25549 274 25946
rect 224 25537 274 25549
rect 390 25946 440 25958
rect 390 25549 396 25946
rect 434 25549 440 25946
rect 390 25537 440 25549
rect -440 22147 -390 22159
rect -440 21750 -434 22147
rect -396 21750 -390 22147
rect -440 21738 -390 21750
rect -274 22147 -224 22159
rect -274 21750 -268 22147
rect -230 21750 -224 22147
rect -274 21738 -224 21750
rect -108 22147 -58 22159
rect -108 21750 -102 22147
rect -64 21750 -58 22147
rect -108 21738 -58 21750
rect 58 22147 108 22159
rect 58 21750 64 22147
rect 102 21750 108 22147
rect 58 21738 108 21750
rect 224 22147 274 22159
rect 224 21750 230 22147
rect 268 21750 274 22147
rect 224 21738 274 21750
rect 390 22147 440 22159
rect 390 21750 396 22147
rect 434 21750 440 22147
rect 390 21738 440 21750
rect -440 21610 -390 21622
rect -440 21213 -434 21610
rect -396 21213 -390 21610
rect -440 21201 -390 21213
rect -274 21610 -224 21622
rect -274 21213 -268 21610
rect -230 21213 -224 21610
rect -274 21201 -224 21213
rect -108 21610 -58 21622
rect -108 21213 -102 21610
rect -64 21213 -58 21610
rect -108 21201 -58 21213
rect 58 21610 108 21622
rect 58 21213 64 21610
rect 102 21213 108 21610
rect 58 21201 108 21213
rect 224 21610 274 21622
rect 224 21213 230 21610
rect 268 21213 274 21610
rect 224 21201 274 21213
rect 390 21610 440 21622
rect 390 21213 396 21610
rect 434 21213 440 21610
rect 390 21201 440 21213
rect -440 17811 -390 17823
rect -440 17414 -434 17811
rect -396 17414 -390 17811
rect -440 17402 -390 17414
rect -274 17811 -224 17823
rect -274 17414 -268 17811
rect -230 17414 -224 17811
rect -274 17402 -224 17414
rect -108 17811 -58 17823
rect -108 17414 -102 17811
rect -64 17414 -58 17811
rect -108 17402 -58 17414
rect 58 17811 108 17823
rect 58 17414 64 17811
rect 102 17414 108 17811
rect 58 17402 108 17414
rect 224 17811 274 17823
rect 224 17414 230 17811
rect 268 17414 274 17811
rect 224 17402 274 17414
rect 390 17811 440 17823
rect 390 17414 396 17811
rect 434 17414 440 17811
rect 390 17402 440 17414
rect -440 17274 -390 17286
rect -440 16877 -434 17274
rect -396 16877 -390 17274
rect -440 16865 -390 16877
rect -274 17274 -224 17286
rect -274 16877 -268 17274
rect -230 16877 -224 17274
rect -274 16865 -224 16877
rect -108 17274 -58 17286
rect -108 16877 -102 17274
rect -64 16877 -58 17274
rect -108 16865 -58 16877
rect 58 17274 108 17286
rect 58 16877 64 17274
rect 102 16877 108 17274
rect 58 16865 108 16877
rect 224 17274 274 17286
rect 224 16877 230 17274
rect 268 16877 274 17274
rect 224 16865 274 16877
rect 390 17274 440 17286
rect 390 16877 396 17274
rect 434 16877 440 17274
rect 390 16865 440 16877
rect -440 13475 -390 13487
rect -440 13078 -434 13475
rect -396 13078 -390 13475
rect -440 13066 -390 13078
rect -274 13475 -224 13487
rect -274 13078 -268 13475
rect -230 13078 -224 13475
rect -274 13066 -224 13078
rect -108 13475 -58 13487
rect -108 13078 -102 13475
rect -64 13078 -58 13475
rect -108 13066 -58 13078
rect 58 13475 108 13487
rect 58 13078 64 13475
rect 102 13078 108 13475
rect 58 13066 108 13078
rect 224 13475 274 13487
rect 224 13078 230 13475
rect 268 13078 274 13475
rect 224 13066 274 13078
rect 390 13475 440 13487
rect 390 13078 396 13475
rect 434 13078 440 13475
rect 390 13066 440 13078
rect -440 12938 -390 12950
rect -440 12541 -434 12938
rect -396 12541 -390 12938
rect -440 12529 -390 12541
rect -274 12938 -224 12950
rect -274 12541 -268 12938
rect -230 12541 -224 12938
rect -274 12529 -224 12541
rect -108 12938 -58 12950
rect -108 12541 -102 12938
rect -64 12541 -58 12938
rect -108 12529 -58 12541
rect 58 12938 108 12950
rect 58 12541 64 12938
rect 102 12541 108 12938
rect 58 12529 108 12541
rect 224 12938 274 12950
rect 224 12541 230 12938
rect 268 12541 274 12938
rect 224 12529 274 12541
rect 390 12938 440 12950
rect 390 12541 396 12938
rect 434 12541 440 12938
rect 390 12529 440 12541
rect -440 9139 -390 9151
rect -440 8742 -434 9139
rect -396 8742 -390 9139
rect -440 8730 -390 8742
rect -274 9139 -224 9151
rect -274 8742 -268 9139
rect -230 8742 -224 9139
rect -274 8730 -224 8742
rect -108 9139 -58 9151
rect -108 8742 -102 9139
rect -64 8742 -58 9139
rect -108 8730 -58 8742
rect 58 9139 108 9151
rect 58 8742 64 9139
rect 102 8742 108 9139
rect 58 8730 108 8742
rect 224 9139 274 9151
rect 224 8742 230 9139
rect 268 8742 274 9139
rect 224 8730 274 8742
rect 390 9139 440 9151
rect 390 8742 396 9139
rect 434 8742 440 9139
rect 390 8730 440 8742
rect -440 8602 -390 8614
rect -440 8205 -434 8602
rect -396 8205 -390 8602
rect -440 8193 -390 8205
rect -274 8602 -224 8614
rect -274 8205 -268 8602
rect -230 8205 -224 8602
rect -274 8193 -224 8205
rect -108 8602 -58 8614
rect -108 8205 -102 8602
rect -64 8205 -58 8602
rect -108 8193 -58 8205
rect 58 8602 108 8614
rect 58 8205 64 8602
rect 102 8205 108 8602
rect 58 8193 108 8205
rect 224 8602 274 8614
rect 224 8205 230 8602
rect 268 8205 274 8602
rect 224 8193 274 8205
rect 390 8602 440 8614
rect 390 8205 396 8602
rect 434 8205 440 8602
rect 390 8193 440 8205
rect -440 4803 -390 4815
rect -440 4406 -434 4803
rect -396 4406 -390 4803
rect -440 4394 -390 4406
rect -274 4803 -224 4815
rect -274 4406 -268 4803
rect -230 4406 -224 4803
rect -274 4394 -224 4406
rect -108 4803 -58 4815
rect -108 4406 -102 4803
rect -64 4406 -58 4803
rect -108 4394 -58 4406
rect 58 4803 108 4815
rect 58 4406 64 4803
rect 102 4406 108 4803
rect 58 4394 108 4406
rect 224 4803 274 4815
rect 224 4406 230 4803
rect 268 4406 274 4803
rect 224 4394 274 4406
rect 390 4803 440 4815
rect 390 4406 396 4803
rect 434 4406 440 4803
rect 390 4394 440 4406
rect -440 4266 -390 4278
rect -440 3869 -434 4266
rect -396 3869 -390 4266
rect -440 3857 -390 3869
rect -274 4266 -224 4278
rect -274 3869 -268 4266
rect -230 3869 -224 4266
rect -274 3857 -224 3869
rect -108 4266 -58 4278
rect -108 3869 -102 4266
rect -64 3869 -58 4266
rect -108 3857 -58 3869
rect 58 4266 108 4278
rect 58 3869 64 4266
rect 102 3869 108 4266
rect 58 3857 108 3869
rect 224 4266 274 4278
rect 224 3869 230 4266
rect 268 3869 274 4266
rect 224 3857 274 3869
rect 390 4266 440 4278
rect 390 3869 396 4266
rect 434 3869 440 4266
rect 390 3857 440 3869
rect -440 467 -390 479
rect -440 70 -434 467
rect -396 70 -390 467
rect -440 58 -390 70
rect -274 467 -224 479
rect -274 70 -268 467
rect -230 70 -224 467
rect -274 58 -224 70
rect -108 467 -58 479
rect -108 70 -102 467
rect -64 70 -58 467
rect -108 58 -58 70
rect 58 467 108 479
rect 58 70 64 467
rect 102 70 108 467
rect 58 58 108 70
rect 224 467 274 479
rect 224 70 230 467
rect 268 70 274 467
rect 224 58 274 70
rect 390 467 440 479
rect 390 70 396 467
rect 434 70 440 467
rect 390 58 440 70
rect -440 -70 -390 -58
rect -440 -467 -434 -70
rect -396 -467 -390 -70
rect -440 -479 -390 -467
rect -274 -70 -224 -58
rect -274 -467 -268 -70
rect -230 -467 -224 -70
rect -274 -479 -224 -467
rect -108 -70 -58 -58
rect -108 -467 -102 -70
rect -64 -467 -58 -70
rect -108 -479 -58 -467
rect 58 -70 108 -58
rect 58 -467 64 -70
rect 102 -467 108 -70
rect 58 -479 108 -467
rect 224 -70 274 -58
rect 224 -467 230 -70
rect 268 -467 274 -70
rect 224 -479 274 -467
rect 390 -70 440 -58
rect 390 -467 396 -70
rect 434 -467 440 -70
rect 390 -479 440 -467
rect -440 -3869 -390 -3857
rect -440 -4266 -434 -3869
rect -396 -4266 -390 -3869
rect -440 -4278 -390 -4266
rect -274 -3869 -224 -3857
rect -274 -4266 -268 -3869
rect -230 -4266 -224 -3869
rect -274 -4278 -224 -4266
rect -108 -3869 -58 -3857
rect -108 -4266 -102 -3869
rect -64 -4266 -58 -3869
rect -108 -4278 -58 -4266
rect 58 -3869 108 -3857
rect 58 -4266 64 -3869
rect 102 -4266 108 -3869
rect 58 -4278 108 -4266
rect 224 -3869 274 -3857
rect 224 -4266 230 -3869
rect 268 -4266 274 -3869
rect 224 -4278 274 -4266
rect 390 -3869 440 -3857
rect 390 -4266 396 -3869
rect 434 -4266 440 -3869
rect 390 -4278 440 -4266
rect -440 -4406 -390 -4394
rect -440 -4803 -434 -4406
rect -396 -4803 -390 -4406
rect -440 -4815 -390 -4803
rect -274 -4406 -224 -4394
rect -274 -4803 -268 -4406
rect -230 -4803 -224 -4406
rect -274 -4815 -224 -4803
rect -108 -4406 -58 -4394
rect -108 -4803 -102 -4406
rect -64 -4803 -58 -4406
rect -108 -4815 -58 -4803
rect 58 -4406 108 -4394
rect 58 -4803 64 -4406
rect 102 -4803 108 -4406
rect 58 -4815 108 -4803
rect 224 -4406 274 -4394
rect 224 -4803 230 -4406
rect 268 -4803 274 -4406
rect 224 -4815 274 -4803
rect 390 -4406 440 -4394
rect 390 -4803 396 -4406
rect 434 -4803 440 -4406
rect 390 -4815 440 -4803
rect -440 -8205 -390 -8193
rect -440 -8602 -434 -8205
rect -396 -8602 -390 -8205
rect -440 -8614 -390 -8602
rect -274 -8205 -224 -8193
rect -274 -8602 -268 -8205
rect -230 -8602 -224 -8205
rect -274 -8614 -224 -8602
rect -108 -8205 -58 -8193
rect -108 -8602 -102 -8205
rect -64 -8602 -58 -8205
rect -108 -8614 -58 -8602
rect 58 -8205 108 -8193
rect 58 -8602 64 -8205
rect 102 -8602 108 -8205
rect 58 -8614 108 -8602
rect 224 -8205 274 -8193
rect 224 -8602 230 -8205
rect 268 -8602 274 -8205
rect 224 -8614 274 -8602
rect 390 -8205 440 -8193
rect 390 -8602 396 -8205
rect 434 -8602 440 -8205
rect 390 -8614 440 -8602
rect -440 -8742 -390 -8730
rect -440 -9139 -434 -8742
rect -396 -9139 -390 -8742
rect -440 -9151 -390 -9139
rect -274 -8742 -224 -8730
rect -274 -9139 -268 -8742
rect -230 -9139 -224 -8742
rect -274 -9151 -224 -9139
rect -108 -8742 -58 -8730
rect -108 -9139 -102 -8742
rect -64 -9139 -58 -8742
rect -108 -9151 -58 -9139
rect 58 -8742 108 -8730
rect 58 -9139 64 -8742
rect 102 -9139 108 -8742
rect 58 -9151 108 -9139
rect 224 -8742 274 -8730
rect 224 -9139 230 -8742
rect 268 -9139 274 -8742
rect 224 -9151 274 -9139
rect 390 -8742 440 -8730
rect 390 -9139 396 -8742
rect 434 -9139 440 -8742
rect 390 -9151 440 -9139
rect -440 -12541 -390 -12529
rect -440 -12938 -434 -12541
rect -396 -12938 -390 -12541
rect -440 -12950 -390 -12938
rect -274 -12541 -224 -12529
rect -274 -12938 -268 -12541
rect -230 -12938 -224 -12541
rect -274 -12950 -224 -12938
rect -108 -12541 -58 -12529
rect -108 -12938 -102 -12541
rect -64 -12938 -58 -12541
rect -108 -12950 -58 -12938
rect 58 -12541 108 -12529
rect 58 -12938 64 -12541
rect 102 -12938 108 -12541
rect 58 -12950 108 -12938
rect 224 -12541 274 -12529
rect 224 -12938 230 -12541
rect 268 -12938 274 -12541
rect 224 -12950 274 -12938
rect 390 -12541 440 -12529
rect 390 -12938 396 -12541
rect 434 -12938 440 -12541
rect 390 -12950 440 -12938
rect -440 -13078 -390 -13066
rect -440 -13475 -434 -13078
rect -396 -13475 -390 -13078
rect -440 -13487 -390 -13475
rect -274 -13078 -224 -13066
rect -274 -13475 -268 -13078
rect -230 -13475 -224 -13078
rect -274 -13487 -224 -13475
rect -108 -13078 -58 -13066
rect -108 -13475 -102 -13078
rect -64 -13475 -58 -13078
rect -108 -13487 -58 -13475
rect 58 -13078 108 -13066
rect 58 -13475 64 -13078
rect 102 -13475 108 -13078
rect 58 -13487 108 -13475
rect 224 -13078 274 -13066
rect 224 -13475 230 -13078
rect 268 -13475 274 -13078
rect 224 -13487 274 -13475
rect 390 -13078 440 -13066
rect 390 -13475 396 -13078
rect 434 -13475 440 -13078
rect 390 -13487 440 -13475
rect -440 -16877 -390 -16865
rect -440 -17274 -434 -16877
rect -396 -17274 -390 -16877
rect -440 -17286 -390 -17274
rect -274 -16877 -224 -16865
rect -274 -17274 -268 -16877
rect -230 -17274 -224 -16877
rect -274 -17286 -224 -17274
rect -108 -16877 -58 -16865
rect -108 -17274 -102 -16877
rect -64 -17274 -58 -16877
rect -108 -17286 -58 -17274
rect 58 -16877 108 -16865
rect 58 -17274 64 -16877
rect 102 -17274 108 -16877
rect 58 -17286 108 -17274
rect 224 -16877 274 -16865
rect 224 -17274 230 -16877
rect 268 -17274 274 -16877
rect 224 -17286 274 -17274
rect 390 -16877 440 -16865
rect 390 -17274 396 -16877
rect 434 -17274 440 -16877
rect 390 -17286 440 -17274
rect -440 -17414 -390 -17402
rect -440 -17811 -434 -17414
rect -396 -17811 -390 -17414
rect -440 -17823 -390 -17811
rect -274 -17414 -224 -17402
rect -274 -17811 -268 -17414
rect -230 -17811 -224 -17414
rect -274 -17823 -224 -17811
rect -108 -17414 -58 -17402
rect -108 -17811 -102 -17414
rect -64 -17811 -58 -17414
rect -108 -17823 -58 -17811
rect 58 -17414 108 -17402
rect 58 -17811 64 -17414
rect 102 -17811 108 -17414
rect 58 -17823 108 -17811
rect 224 -17414 274 -17402
rect 224 -17811 230 -17414
rect 268 -17811 274 -17414
rect 224 -17823 274 -17811
rect 390 -17414 440 -17402
rect 390 -17811 396 -17414
rect 434 -17811 440 -17414
rect 390 -17823 440 -17811
rect -440 -21213 -390 -21201
rect -440 -21610 -434 -21213
rect -396 -21610 -390 -21213
rect -440 -21622 -390 -21610
rect -274 -21213 -224 -21201
rect -274 -21610 -268 -21213
rect -230 -21610 -224 -21213
rect -274 -21622 -224 -21610
rect -108 -21213 -58 -21201
rect -108 -21610 -102 -21213
rect -64 -21610 -58 -21213
rect -108 -21622 -58 -21610
rect 58 -21213 108 -21201
rect 58 -21610 64 -21213
rect 102 -21610 108 -21213
rect 58 -21622 108 -21610
rect 224 -21213 274 -21201
rect 224 -21610 230 -21213
rect 268 -21610 274 -21213
rect 224 -21622 274 -21610
rect 390 -21213 440 -21201
rect 390 -21610 396 -21213
rect 434 -21610 440 -21213
rect 390 -21622 440 -21610
rect -440 -21750 -390 -21738
rect -440 -22147 -434 -21750
rect -396 -22147 -390 -21750
rect -440 -22159 -390 -22147
rect -274 -21750 -224 -21738
rect -274 -22147 -268 -21750
rect -230 -22147 -224 -21750
rect -274 -22159 -224 -22147
rect -108 -21750 -58 -21738
rect -108 -22147 -102 -21750
rect -64 -22147 -58 -21750
rect -108 -22159 -58 -22147
rect 58 -21750 108 -21738
rect 58 -22147 64 -21750
rect 102 -22147 108 -21750
rect 58 -22159 108 -22147
rect 224 -21750 274 -21738
rect 224 -22147 230 -21750
rect 268 -22147 274 -21750
rect 224 -22159 274 -22147
rect 390 -21750 440 -21738
rect 390 -22147 396 -21750
rect 434 -22147 440 -21750
rect 390 -22159 440 -22147
rect -440 -25549 -390 -25537
rect -440 -25946 -434 -25549
rect -396 -25946 -390 -25549
rect -440 -25958 -390 -25946
rect -274 -25549 -224 -25537
rect -274 -25946 -268 -25549
rect -230 -25946 -224 -25549
rect -274 -25958 -224 -25946
rect -108 -25549 -58 -25537
rect -108 -25946 -102 -25549
rect -64 -25946 -58 -25549
rect -108 -25958 -58 -25946
rect 58 -25549 108 -25537
rect 58 -25946 64 -25549
rect 102 -25946 108 -25549
rect 58 -25958 108 -25946
rect 224 -25549 274 -25537
rect 224 -25946 230 -25549
rect 268 -25946 274 -25549
rect 224 -25958 274 -25946
rect 390 -25549 440 -25537
rect 390 -25946 396 -25549
rect 434 -25946 440 -25549
rect 390 -25958 440 -25946
<< properties >>
string FIXED_BBOX -563 -26077 563 26077
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.350 l 17 m 12 nx 6 wmin 0.350 lmin 0.50 rho 319.8 val 16.646k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
