magic
tech sky130A
magscale 1 2
timestamp 1717511437
<< checkpaint >>
rect -575 -1578 4337 2888
<< error_p >>
rect 12785 13275 12820 13309
rect 12786 13256 12820 13275
rect 12687 13126 12694 13144
rect 12616 12995 12674 13001
rect 12616 12961 12628 12995
rect 12616 12955 12674 12961
rect 12616 12675 12674 12681
rect 12616 12641 12628 12675
rect 12616 12635 12674 12641
rect 12616 12567 12674 12573
rect 12616 12544 12628 12567
rect 12616 12527 12674 12544
rect 12588 12499 12687 12516
rect 12616 12247 12674 12253
rect 12616 12213 12628 12247
rect 12616 12207 12674 12213
rect 12805 11899 12820 13256
rect 12839 13222 12874 13256
rect 12839 11899 12873 13222
rect 12985 13154 13043 13160
rect 12985 13120 12997 13154
rect 12985 13114 13043 13120
rect 13723 13048 13781 13054
rect 13723 13014 13735 13048
rect 13723 13008 13781 13014
rect 12985 12942 13043 12948
rect 12985 12908 12997 12942
rect 12985 12902 13043 12908
rect 12985 12834 13043 12840
rect 13723 12836 13781 12842
rect 12985 12800 12997 12834
rect 13723 12802 13735 12836
rect 12985 12794 13043 12800
rect 13723 12796 13781 12802
rect 13723 12728 13781 12734
rect 13723 12694 13735 12728
rect 13723 12688 13781 12694
rect 12985 12622 13043 12628
rect 12985 12588 12997 12622
rect 12985 12582 13043 12588
rect 13155 12563 13189 12581
rect 13577 12563 13611 12581
rect 13155 12527 13225 12563
rect 12985 12514 13043 12520
rect 12985 12480 12997 12514
rect 13172 12493 13243 12527
rect 12985 12474 13043 12480
rect 12985 12302 13043 12308
rect 12985 12268 12997 12302
rect 12985 12262 13043 12268
rect 12985 12194 13043 12200
rect 12985 12160 12997 12194
rect 12985 12154 13043 12160
rect 12985 11982 13043 11988
rect 12985 11948 12997 11982
rect 12985 11942 13043 11948
rect 12839 11865 12854 11899
rect 13172 11846 13242 12493
rect 13354 12425 13412 12431
rect 13354 12391 13366 12425
rect 13354 12385 13412 12391
rect 13354 12231 13412 12237
rect 13354 12197 13366 12231
rect 13354 12191 13412 12197
rect 13354 12123 13412 12129
rect 13354 12089 13366 12123
rect 13354 12083 13412 12089
rect 13354 11929 13412 11935
rect 13354 11895 13366 11929
rect 13354 11889 13412 11895
rect 13172 11810 13225 11846
rect 13541 11793 13611 12563
rect 13723 12516 13781 12522
rect 13723 12482 13735 12516
rect 13723 12476 13781 12482
rect 13893 12457 13927 12475
rect 13893 12421 13963 12457
rect 13723 12408 13781 12414
rect 13723 12374 13735 12408
rect 13910 12387 13981 12421
rect 13723 12368 13781 12374
rect 13723 12196 13781 12202
rect 13723 12162 13735 12196
rect 13723 12156 13781 12162
rect 13723 12088 13781 12094
rect 13723 12054 13735 12088
rect 13723 12048 13781 12054
rect 13723 11876 13781 11882
rect 13723 11842 13735 11876
rect 13723 11836 13781 11842
rect 13541 11757 13594 11793
rect 13910 11740 13980 12387
rect 14092 12319 14150 12325
rect 14092 12285 14104 12319
rect 14092 12279 14150 12285
rect 14092 12125 14150 12131
rect 14092 12091 14104 12125
rect 14092 12085 14150 12091
rect 14092 12017 14150 12023
rect 14092 11983 14104 12017
rect 14092 11977 14150 11983
rect 14092 11823 14150 11829
rect 14092 11789 14104 11823
rect 14092 11783 14150 11789
rect 13910 11704 13963 11740
rect 18382 2712 18417 2746
rect 18383 2693 18417 2712
rect 18217 2184 18287 2186
rect 18402 1554 18417 2693
rect 18436 2659 18471 2693
rect 18436 1554 18470 2659
rect 18566 2131 18636 2133
rect 18436 1520 18451 1554
rect 18751 1501 18766 2693
rect 18785 1501 18819 2747
rect 18931 2684 18989 2690
rect 18931 2650 18943 2684
rect 18931 2644 18989 2650
rect 18931 2490 18989 2496
rect 18931 2456 18943 2490
rect 18931 2450 18989 2456
rect 18931 2382 18989 2388
rect 18931 2348 18943 2382
rect 18931 2342 18989 2348
rect 19101 2201 19135 2219
rect 18931 2188 18989 2194
rect 18931 2154 18943 2188
rect 19101 2165 19171 2201
rect 18931 2148 18989 2154
rect 19118 2131 19189 2165
rect 19469 2131 19504 2165
rect 18931 2080 18989 2086
rect 18931 2046 18943 2080
rect 18931 2040 18989 2046
rect 18931 1886 18989 1892
rect 18931 1852 18943 1886
rect 18931 1846 18989 1852
rect 18931 1778 18989 1784
rect 18931 1744 18943 1778
rect 18931 1738 18989 1744
rect 18931 1584 18989 1590
rect 18931 1550 18943 1584
rect 18931 1544 18989 1550
rect 18785 1467 18800 1501
rect 19118 1448 19188 2131
rect 19470 2112 19504 2131
rect 19300 2063 19358 2069
rect 19300 2029 19312 2063
rect 19300 2023 19358 2029
rect 19300 1851 19358 1857
rect 19300 1817 19312 1851
rect 19300 1811 19358 1817
rect 19300 1743 19358 1749
rect 19300 1709 19312 1743
rect 19300 1703 19358 1709
rect 19300 1531 19358 1537
rect 19300 1497 19312 1531
rect 19300 1491 19358 1497
rect 19118 1412 19171 1448
rect 19489 1395 19504 2112
rect 19523 2078 19558 2112
rect 19523 1395 19557 2078
rect 19839 2059 19873 2077
rect 19839 2023 19909 2059
rect 19669 2010 19727 2016
rect 19669 1976 19681 2010
rect 19856 1989 19927 2023
rect 20207 1989 20242 2023
rect 19669 1970 19727 1976
rect 19669 1798 19727 1804
rect 19669 1764 19681 1798
rect 19669 1758 19727 1764
rect 19669 1690 19727 1696
rect 19669 1656 19681 1690
rect 19669 1650 19727 1656
rect 19669 1478 19727 1484
rect 19669 1444 19681 1478
rect 19669 1438 19727 1444
rect 19523 1361 19538 1395
rect 19856 1342 19926 1989
rect 20208 1970 20242 1989
rect 20038 1921 20096 1927
rect 20038 1887 20050 1921
rect 20038 1881 20096 1887
rect 20038 1727 20096 1733
rect 20038 1693 20050 1727
rect 20038 1687 20096 1693
rect 20038 1619 20096 1625
rect 20038 1585 20050 1619
rect 20038 1579 20096 1585
rect 20038 1425 20096 1431
rect 20038 1391 20050 1425
rect 20038 1385 20096 1391
rect 19856 1306 19909 1342
rect 20227 1289 20242 1970
rect 20261 1936 20296 1970
rect 20261 1289 20295 1936
rect 20407 1868 20465 1874
rect 20407 1834 20419 1868
rect 20407 1828 20465 1834
rect 20407 1674 20465 1680
rect 20407 1640 20419 1674
rect 20407 1634 20465 1640
rect 20407 1566 20465 1572
rect 20407 1532 20419 1566
rect 20407 1526 20465 1532
rect 20407 1372 20465 1378
rect 20407 1338 20419 1372
rect 20407 1332 20465 1338
rect 20261 1255 20276 1289
rect 20596 1236 20611 1970
rect 20630 1236 20664 2024
rect 20760 1813 20830 1815
rect 20630 1202 20645 1236
rect 20945 1183 20960 2375
rect 20979 1183 21013 2429
rect 21125 2366 21183 2372
rect 21125 2332 21137 2366
rect 21125 2326 21183 2332
rect 21125 2172 21183 2178
rect 21125 2138 21137 2172
rect 21125 2132 21183 2138
rect 21125 2064 21183 2070
rect 21125 2030 21137 2064
rect 21125 2024 21183 2030
rect 21125 1870 21183 1876
rect 21125 1836 21137 1870
rect 21125 1830 21183 1836
rect 21125 1762 21183 1768
rect 21125 1728 21137 1762
rect 21125 1722 21183 1728
rect 21125 1568 21183 1574
rect 21125 1534 21137 1568
rect 21125 1528 21183 1534
rect 21125 1460 21183 1466
rect 21125 1426 21137 1460
rect 21125 1420 21183 1426
rect 21125 1266 21183 1272
rect 21125 1232 21137 1266
rect 21125 1226 21183 1232
rect 20979 1149 20994 1183
rect 28493 968 28528 1002
rect 28494 949 28528 968
rect 28513 436 28528 949
rect 28547 915 28582 949
rect 30832 915 30867 949
rect 33225 932 33259 950
rect 28547 436 28581 915
rect 30833 896 30867 915
rect 28547 402 28562 436
rect 30852 383 30867 896
rect 30886 862 30921 896
rect 30886 383 30920 862
rect 30886 349 30901 383
rect 33189 330 33259 932
rect 33189 294 33242 330
<< error_s >>
rect 298 1209 333 1234
rect -17 1200 333 1209
rect -17 1181 17 1200
rect 299 1181 333 1200
rect -17 1155 738 1181
rect -8 -159 738 1155
rect 1366 26 1368 1209
rect 25777 1917 25823 1934
rect 25749 1889 25851 1906
rect 25749 1706 25851 1727
rect 25777 1678 25823 1699
rect 25749 1306 25851 1309
rect 25777 1278 25823 1281
rect 26155 1038 26189 1056
rect 26155 1002 26225 1038
rect 26172 968 26243 1002
rect 26172 489 26242 968
rect 24455 434 24490 468
rect 26172 453 26225 489
rect 24456 415 24490 434
rect 24286 366 24344 372
rect 24286 332 24298 366
rect 24286 326 24344 332
rect 24286 172 24344 178
rect 24286 138 24298 172
rect 24286 132 24344 138
rect 24475 36 24490 415
rect 24509 381 24544 415
rect 24824 381 24859 415
rect 24509 36 24543 381
rect 24825 362 24859 381
rect 24655 313 24713 319
rect 24655 279 24667 313
rect 24655 273 24713 279
rect 24655 119 24713 125
rect 24655 85 24667 119
rect 24655 79 24713 85
rect 24509 2 24524 36
rect 24844 -17 24859 362
rect 24878 328 24913 362
rect 25193 328 25228 362
rect 24878 -17 24912 328
rect 25194 309 25228 328
rect 25024 260 25082 266
rect 25024 226 25036 260
rect 25024 220 25082 226
rect 25024 66 25082 72
rect 25024 32 25036 66
rect 25024 26 25082 32
rect 24878 -51 24893 -17
rect 25213 -70 25228 309
rect 25247 275 25282 309
rect 25247 -70 25281 275
rect 25393 207 25451 213
rect 25393 173 25405 207
rect 25393 167 25451 173
rect 25393 13 25451 19
rect 25393 -21 25405 13
rect 25393 -27 25451 -21
rect 25247 -104 25262 -70
rect -8 -167 299 -159
rect 318 -176 333 -159
rect 352 -176 386 -159
rect 352 -210 367 -176
use op5  x1
timestamp 1717511434
transform 1 0 12487 0 1 13516
box -53 -12422 8878 1335
use Resistor492k_1  x2
timestamp 1717511435
transform 1 0 23704 0 1 1441
box 0 -1600 200 200
use Resistor492k_1  x3
timestamp 1717511435
transform 1 0 23904 0 1 1441
box 0 -1600 200 200
use Resistor50k_1  x4
timestamp 1717511435
transform 1 0 24151 0 1 453
box -47 -612 1482 200
use Startup  x5
timestamp 1717511437
transform 1 0 25686 0 1 2106
box -53 -1865 7934 2699
use sky130_fd_pr__pfet_01v8_M47T9Z  XM1
timestamp 0
transform 1 0 158 0 1 529
box -211 -741 211 741
use sky130_fd_pr__pfet_01v8_M47T9Z  XM2
timestamp 0
transform 1 0 527 0 1 476
box -211 -741 211 741
use sky130_fd_pr__pfet_01v8_6H4VWJ  XM15
timestamp 0
transform 1 0 1881 0 1 655
box -1196 -973 1196 973
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  XQ1 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1716538025
transform 1 0 0 0 1 -159
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  XQ2
array 0 7 1288 0 0 1288
timestamp 1716538025
transform 1 0 1340 0 1 0
box 0 0 1340 1340
<< end >>
