magic
tech sky130A
magscale 1 2
timestamp 1717383984
<< nwell >>
rect -1723 -164 1723 198
<< pmos >>
rect -1629 -64 -29 136
rect 29 -64 1629 136
<< pdiff >>
rect -1687 124 -1629 136
rect -1687 -52 -1675 124
rect -1641 -52 -1629 124
rect -1687 -64 -1629 -52
rect -29 124 29 136
rect -29 -52 -17 124
rect 17 -52 29 124
rect -29 -64 29 -52
rect 1629 124 1687 136
rect 1629 -52 1641 124
rect 1675 -52 1687 124
rect 1629 -64 1687 -52
<< pdiffc >>
rect -1675 -52 -1641 124
rect -17 -52 17 124
rect 1641 -52 1675 124
<< poly >>
rect -1629 136 -29 162
rect 29 136 1629 162
rect -1629 -111 -29 -64
rect -1629 -145 -1613 -111
rect -45 -145 -29 -111
rect -1629 -161 -29 -145
rect 29 -111 1629 -64
rect 29 -145 45 -111
rect 1613 -145 1629 -111
rect 29 -161 1629 -145
<< polycont >>
rect -1613 -145 -45 -111
rect 45 -145 1613 -111
<< locali >>
rect -1675 124 -1641 140
rect -1675 -68 -1641 -52
rect -17 124 17 140
rect -17 -68 17 -52
rect 1641 124 1675 140
rect 1641 -68 1675 -52
rect -1629 -145 -1613 -111
rect -45 -145 -29 -111
rect 29 -145 45 -111
rect 1613 -145 1629 -111
<< viali >>
rect -1675 -52 -1641 124
rect -17 -52 17 124
rect 1641 -52 1675 124
rect -1613 -145 -45 -111
rect 45 -145 1613 -111
<< metal1 >>
rect -1681 124 -1635 136
rect -1681 -52 -1675 124
rect -1641 -52 -1635 124
rect -1681 -64 -1635 -52
rect -23 124 23 136
rect -23 -52 -17 124
rect 17 -52 23 124
rect -23 -64 23 -52
rect 1635 124 1681 136
rect 1635 -52 1641 124
rect 1675 -52 1681 124
rect 1635 -64 1681 -52
rect -1625 -111 -33 -105
rect -1625 -145 -1613 -111
rect -45 -145 -33 -111
rect -1625 -151 -33 -145
rect 33 -111 1625 -105
rect 33 -145 45 -111
rect 1613 -145 1625 -111
rect 33 -151 1625 -145
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 8 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
