magic
tech sky130A
magscale 1 2
timestamp 1720116957
<< psubdiff >>
rect -594 846 -532 880
rect 5166 846 5228 880
rect -594 805 -560 846
rect 5194 805 5228 846
rect -594 -78 -560 -37
rect 5194 -78 5228 -37
rect -594 -112 -532 -78
rect 5166 -112 5228 -78
<< psubdiffcont >>
rect -532 846 5166 880
rect -594 -37 -560 805
rect 5194 -37 5228 805
rect -532 -112 5166 -78
<< poly >>
rect -462 430 -370 446
rect -462 396 -446 430
rect -412 396 -370 430
rect -462 380 -370 396
rect 5004 430 5096 446
rect 5004 396 5046 430
rect 5080 396 5096 430
rect 5004 380 5096 396
rect -462 288 -370 304
rect -462 254 -446 288
rect -412 254 -370 288
rect -462 238 -370 254
rect 5004 288 5096 304
rect 5004 254 5046 288
rect 5080 254 5096 288
rect 5004 238 5096 254
<< polycont >>
rect -446 396 -412 430
rect 5046 396 5080 430
rect -446 254 -412 288
rect 5046 254 5080 288
<< locali >>
rect -446 430 -412 470
rect -446 380 -412 396
rect 5046 430 5080 470
rect 5046 380 5080 396
rect -446 288 -412 304
rect -446 214 -412 254
rect 5046 288 5080 304
rect 5046 214 5080 254
<< viali >>
rect -594 846 -532 880
rect -532 846 5166 880
rect 5166 846 5228 880
rect -594 805 -560 846
rect -594 -37 -560 805
rect 5194 805 5228 846
rect -446 396 -412 430
rect 5046 396 5080 430
rect -446 254 -412 288
rect 5046 254 5080 288
rect -594 -78 -560 -37
rect 5194 -37 5228 805
rect 5194 -78 5228 -37
rect -594 -112 -532 -78
rect -532 -112 5166 -78
rect 5166 -112 5228 -78
<< metal1 >>
rect -600 886 -554 892
rect 5188 886 5234 892
rect -606 880 5240 886
rect -606 840 -594 880
rect -600 -72 -594 840
rect -606 -112 -594 -72
rect -560 840 5194 846
rect -560 -72 -554 840
rect -526 766 5160 812
rect -526 2 -480 766
rect -452 636 -305 648
rect -452 480 -367 636
rect -315 480 -305 636
rect 2294 630 2340 766
rect 4939 636 5086 648
rect -452 468 -305 480
rect 4939 480 4949 636
rect 5001 480 5086 636
rect 4939 468 5086 480
rect -452 430 -406 468
rect -452 396 -446 430
rect -412 396 -406 430
rect -452 384 -406 396
rect 1600 390 2188 436
rect 2142 365 2188 390
rect 2994 387 3004 439
rect 4288 387 4298 439
rect 5040 430 5086 468
rect 5040 396 5046 430
rect 5080 396 5086 430
rect 5040 384 5086 396
rect 2142 319 2492 365
rect -452 288 -406 300
rect -452 254 -446 288
rect -412 254 -406 288
rect -452 216 -406 254
rect 336 245 346 297
rect 1630 245 1640 297
rect 2446 294 2492 319
rect 2446 248 3022 294
rect 5040 288 5086 300
rect 5040 254 5046 288
rect 5080 254 5086 288
rect 5040 216 5086 254
rect -452 204 -305 216
rect -452 48 -367 204
rect -315 48 -305 204
rect 4939 204 5086 216
rect -452 36 -305 48
rect 2294 2 2340 72
rect 4939 48 4949 204
rect 5001 48 5086 204
rect 4939 36 5086 48
rect 5114 2 5160 766
rect -526 -44 5160 2
rect 5188 -72 5194 840
rect -560 -78 5194 -72
rect 5228 840 5240 880
rect 5228 -72 5234 840
rect 5228 -112 5240 -72
rect -606 -118 5240 -112
rect -600 -124 -554 -118
rect 5188 -124 5234 -118
<< via1 >>
rect -367 480 -315 636
rect 4949 480 5001 636
rect 3004 387 4288 439
rect 346 245 1630 297
rect -367 48 -315 204
rect 4949 48 5001 204
<< metal2 >>
rect -369 636 -313 646
rect -369 470 -313 480
rect 4947 636 5003 646
rect 4947 470 5003 480
rect 2446 439 4288 449
rect 2446 387 3004 439
rect 2446 378 4288 387
rect 2116 377 4288 378
rect 2116 307 2518 377
rect 346 306 2518 307
rect 346 297 2188 306
rect 1630 245 2188 297
rect 346 235 2188 245
rect -369 204 -313 214
rect -369 38 -313 48
rect 4947 204 5003 214
rect 4947 38 5003 48
<< via2 >>
rect -369 480 -367 636
rect -367 480 -315 636
rect -315 480 -313 636
rect 4947 480 4949 636
rect 4949 480 5001 636
rect 5001 480 5003 636
rect -369 48 -367 204
rect -367 48 -315 204
rect -315 48 -313 204
rect 4947 48 4949 204
rect 4949 48 5001 204
rect 5001 48 5003 204
<< metal3 >>
rect -379 636 -303 641
rect 4937 636 5013 641
rect -383 480 -373 636
rect -309 480 -299 636
rect 4937 480 4947 636
rect 5003 480 5013 636
rect -379 475 -303 480
rect 4937 475 5013 480
rect 4945 372 5005 475
rect -371 312 5005 372
rect -371 209 -311 312
rect -379 204 -303 209
rect 4937 204 5013 209
rect -379 48 -369 204
rect -313 48 -303 204
rect 4933 48 4943 204
rect 5007 48 5017 204
rect -379 43 -303 48
rect 4937 43 5013 48
<< via3 >>
rect -373 480 -369 636
rect -369 480 -313 636
rect -313 480 -309 636
rect 4943 48 4947 204
rect 4947 48 5003 204
rect 5003 48 5007 204
<< metal4 >>
rect -374 636 -308 637
rect -374 480 -373 636
rect -309 480 -308 636
rect -374 479 -308 480
rect -371 372 -311 479
rect -371 312 5005 372
rect 4945 205 5005 312
rect 4942 204 5008 205
rect 4942 48 4943 204
rect 5007 48 5008 204
rect 4942 47 5008 48
use sky130_fd_pr__nfet_01v8_2A7GYR  sky130_fd_pr__nfet_01v8_2A7GYR_0
timestamp 1720116957
transform 1 0 5019 0 1 558
box -73 -116 73 116
use sky130_fd_pr__nfet_01v8_2A7GYR  sky130_fd_pr__nfet_01v8_2A7GYR_1
timestamp 1720116957
transform 1 0 -385 0 1 558
box -73 -116 73 116
use sky130_fd_pr__nfet_01v8_2A7GYR  sky130_fd_pr__nfet_01v8_2A7GYR_2
timestamp 1720116957
transform 1 0 5019 0 1 126
box -73 -116 73 116
use sky130_fd_pr__nfet_01v8_2A7GYR  sky130_fd_pr__nfet_01v8_2A7GYR_4
timestamp 1720116957
transform 1 0 -385 0 1 126
box -73 -116 73 116
use sky130_fd_pr__nfet_01v8_7RJ44K  sky130_fd_pr__nfet_01v8_7RJ44K_0
timestamp 1720116957
transform 1 0 2317 0 1 157
box -2687 -147 2687 147
use sky130_fd_pr__nfet_01v8_G26DVX  sky130_fd_pr__nfet_01v8_G26DVX_0
timestamp 1720116957
transform 1 0 2317 0 -1 558
box -2687 -178 2687 178
<< labels >>
flabel metal1 5231 853 5231 853 0 FreeSans 160 0 0 0 AVSS
port 0 nsew
flabel metal1 2316 -10 2316 -10 0 FreeSans 160 0 0 0 S
port 1 nsew
flabel metal2 2613 401 2613 401 0 FreeSans 160 0 0 0 PLUS
port 2 nsew
flabel metal1 2556 285 2556 285 0 FreeSans 160 0 0 0 MINUS
port 3 nsew
flabel metal3 4973 406 4973 406 0 FreeSans 160 0 0 0 D3
port 4 nsew
flabel metal4 4984 293 4984 293 0 FreeSans 160 0 0 0 D4
port 5 nsew
<< end >>
