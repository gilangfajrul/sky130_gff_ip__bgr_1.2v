magic
tech sky130A
magscale 1 2
timestamp 1720267898
<< nwell >>
rect -176 -494 4422 430
<< nsubdiff >>
rect -140 360 -80 394
rect 4326 360 4386 394
rect -140 334 -106 360
rect 4352 334 4386 360
rect -140 -424 -106 -398
rect 4352 -424 4386 -398
rect -140 -458 -80 -424
rect 4326 -458 4386 -424
<< nsubdiffcont >>
rect -80 360 4326 394
rect -140 -398 -106 334
rect 4352 -398 4386 334
rect -80 -458 4326 -424
<< poly >>
rect 6 75 36 98
rect -56 59 36 75
rect -56 25 -40 59
rect -6 25 36 59
rect -56 9 36 25
rect 4210 74 4240 126
rect 4210 58 4302 74
rect 4210 24 4252 58
rect 4286 24 4302 58
rect 4210 8 4302 24
rect -56 -89 36 -73
rect -56 -123 -40 -89
rect -6 -123 36 -89
rect -56 -139 36 -123
rect 6 -144 36 -139
rect 4210 -89 4302 -73
rect 4210 -123 4252 -89
rect 4286 -123 4302 -89
rect 4210 -139 4302 -123
rect 4210 -152 4240 -139
<< polycont >>
rect -40 25 -6 59
rect 4252 24 4286 58
rect -40 -123 -6 -89
rect 4252 -123 4286 -89
<< locali >>
rect -40 59 -6 111
rect -40 9 -6 25
rect 4252 58 4286 114
rect 4252 8 4286 24
rect -40 -89 -6 -73
rect -40 -175 -6 -123
rect 4252 -89 4286 -73
rect 4252 -173 4286 -123
<< viali >>
rect -140 360 -80 394
rect -80 360 4326 394
rect 4326 360 4386 394
rect -140 334 -106 360
rect -140 -398 -106 334
rect 4352 334 4386 360
rect -40 25 -6 59
rect 4252 24 4286 58
rect -40 -123 -6 -89
rect 4252 -123 4286 -89
rect -140 -424 -106 -398
rect 4352 -398 4386 334
rect 4352 -424 4386 -398
rect -140 -458 -80 -424
rect -80 -458 4326 -424
rect 4326 -458 4386 -424
<< metal1 >>
rect -146 400 -100 406
rect 4346 400 4392 406
rect -152 394 4398 400
rect -152 354 -140 394
rect -146 -418 -140 354
rect -152 -458 -140 -418
rect -106 354 4352 360
rect -106 -418 -100 354
rect -24 108 79 300
rect -46 107 79 108
rect -46 106 88 107
rect 2087 106 2097 282
rect 2149 106 2159 282
rect 4179 124 4282 300
rect 4179 106 4292 124
rect -46 59 0 106
rect -46 25 -40 59
rect -6 25 0 59
rect -46 13 0 25
rect 42 59 88 106
rect 4158 105 4292 106
rect 42 19 620 59
rect 1594 19 2669 65
rect 88 13 620 19
rect 4158 -9 4204 105
rect 4246 58 4292 105
rect 4246 24 4252 58
rect 4286 24 4292 58
rect 4246 12 4292 24
rect 1552 -55 4204 -9
rect -46 -89 0 -77
rect -46 -123 -40 -89
rect -6 -123 0 -89
rect -46 -170 0 -123
rect 1552 -129 1598 -55
rect 2100 -129 4204 -83
rect -46 -176 60 -170
rect -43 -370 60 -176
rect 2100 -182 2146 -129
rect 4158 -170 4204 -129
rect 4246 -89 4292 -77
rect 4246 -123 4252 -89
rect 4286 -123 4292 -89
rect 4246 -170 4292 -123
rect 4158 -179 4292 -170
rect 2087 -358 2097 -182
rect 2149 -358 2159 -182
rect 2100 -418 2146 -358
rect 4158 -370 4261 -179
rect 4158 -418 4204 -370
rect 4346 -418 4352 354
rect -106 -424 4352 -418
rect 4386 354 4398 394
rect 4386 -418 4392 354
rect 4386 -458 4398 -418
rect -152 -464 4398 -458
rect -146 -470 -100 -464
rect 4346 -470 4392 -464
<< via1 >>
rect 2097 106 2149 282
rect 2097 -358 2149 -182
<< metal2 >>
rect 2097 282 2149 292
rect 2097 -182 2149 106
rect 2097 -368 2149 -358
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_0
timestamp 1717765832
transform 1 0 4225 0 1 206
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_1
timestamp 1717765832
transform 1 0 4225 0 1 -270
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_2
timestamp 1717765832
transform 1 0 21 0 1 206
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_4
timestamp 1717765832
transform 1 0 21 0 1 -270
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_8RMJP2  sky130_fd_pr__pfet_01v8_8RMJP2_0
timestamp 1717765832
transform 1 0 2123 0 1 -234
box -2123 -198 2123 164
use sky130_fd_pr__pfet_01v8_CVRJBD  sky130_fd_pr__pfet_01v8_CVRJBD_1
timestamp 1717765832
transform 1 0 2123 0 1 170
box -2123 -164 2123 198
<< labels >>
flabel metal1 62 30 62 30 0 FreeSans 1600 0 0 0 D3
port 1 nsew
flabel metal1 4184 55 4184 55 0 FreeSans 1600 0 0 0 D2
port 2 nsew
flabel metal1 17 -267 17 -267 0 FreeSans 1600 0 0 0 D4
port 3 nsew
flabel metal1 2119 -408 2119 -408 0 FreeSans 1600 0 0 0 VDDE
port 4 nsew
<< end >>
