.param i_tail = 2.00e-06
.param lrz = 3.72e+01
.param mrz = 1.00e+00
.param lrs = 3.73e-01
.param mrs = 1.00e+00
.param mc = 4.00e+00
.param wc = 3.09e-01
.param w0 = 3.34
.param l0 = 0.60
.param nf0 = 1.00
.param w1 = 4.85
.param l1 = 0.60
.param nf1 = 1.00
.param w2 = 0.52
.param l2 = 0.60
.param nf2 = 1.00
.param w3 = 2.32
.param l3 = 0.80
.param nf3 = 1.00
.param w4 = 0.03
.param l4 = 0.60
.param nf4 = 1.00
