magic
tech sky130A
magscale 1 2
timestamp 1717262354
<< nwell >>
rect -4181 -164 4181 198
<< pmos >>
rect -4087 -64 -2087 136
rect -2029 -64 -29 136
rect 29 -64 2029 136
rect 2087 -64 4087 136
<< pdiff >>
rect -4145 124 -4087 136
rect -4145 -52 -4133 124
rect -4099 -52 -4087 124
rect -4145 -64 -4087 -52
rect -2087 124 -2029 136
rect -2087 -52 -2075 124
rect -2041 -52 -2029 124
rect -2087 -64 -2029 -52
rect -29 124 29 136
rect -29 -52 -17 124
rect 17 -52 29 124
rect -29 -64 29 -52
rect 2029 124 2087 136
rect 2029 -52 2041 124
rect 2075 -52 2087 124
rect 2029 -64 2087 -52
rect 4087 124 4145 136
rect 4087 -52 4099 124
rect 4133 -52 4145 124
rect 4087 -64 4145 -52
<< pdiffc >>
rect -4133 -52 -4099 124
rect -2075 -52 -2041 124
rect -17 -52 17 124
rect 2041 -52 2075 124
rect 4099 -52 4133 124
<< poly >>
rect -4087 136 -2087 162
rect -2029 136 -29 162
rect 29 136 2029 162
rect 2087 136 4087 162
rect -4087 -111 -2087 -64
rect -4087 -128 -3579 -111
rect -3595 -145 -3579 -128
rect -2595 -128 -2087 -111
rect -2029 -111 -29 -64
rect -2029 -128 -1521 -111
rect -2595 -145 -2579 -128
rect -3595 -161 -2579 -145
rect -1537 -145 -1521 -128
rect -537 -128 -29 -111
rect 29 -111 2029 -64
rect 29 -128 537 -111
rect -537 -145 -521 -128
rect -1537 -161 -521 -145
rect 521 -145 537 -128
rect 1521 -128 2029 -111
rect 2087 -111 4087 -64
rect 2087 -128 2595 -111
rect 1521 -145 1537 -128
rect 521 -161 1537 -145
rect 2579 -145 2595 -128
rect 3579 -128 4087 -111
rect 3579 -145 3595 -128
rect 2579 -161 3595 -145
<< polycont >>
rect -3579 -145 -2595 -111
rect -1521 -145 -537 -111
rect 537 -145 1521 -111
rect 2595 -145 3579 -111
<< locali >>
rect -4133 124 -4099 140
rect -4133 -68 -4099 -52
rect -2075 124 -2041 140
rect -2075 -68 -2041 -52
rect -17 124 17 140
rect -17 -68 17 -52
rect 2041 124 2075 140
rect 2041 -68 2075 -52
rect 4099 124 4133 140
rect 4099 -68 4133 -52
rect -3595 -145 -3579 -111
rect -2595 -145 -2579 -111
rect -1537 -145 -1521 -111
rect -537 -145 -521 -111
rect 521 -145 537 -111
rect 1521 -145 1537 -111
rect 2579 -145 2595 -111
rect 3579 -145 3595 -111
<< viali >>
rect -4133 -52 -4099 124
rect -2075 -52 -2041 124
rect -17 -52 17 124
rect 2041 -52 2075 124
rect 4099 -52 4133 124
rect -3579 -145 -2595 -111
rect -1521 -145 -537 -111
rect 537 -145 1521 -111
rect 2595 -145 3579 -111
<< metal1 >>
rect -4139 124 -4093 136
rect -4139 -52 -4133 124
rect -4099 -52 -4093 124
rect -4139 -64 -4093 -52
rect -2081 124 -2035 136
rect -2081 -52 -2075 124
rect -2041 -52 -2035 124
rect -2081 -64 -2035 -52
rect -23 124 23 136
rect -23 -52 -17 124
rect 17 -52 23 124
rect -23 -64 23 -52
rect 2035 124 2081 136
rect 2035 -52 2041 124
rect 2075 -52 2081 124
rect 2035 -64 2081 -52
rect 4093 124 4139 136
rect 4093 -52 4099 124
rect 4133 -52 4139 124
rect 4093 -64 4139 -52
rect -3591 -111 -2583 -105
rect -3591 -145 -3579 -111
rect -2595 -145 -2583 -111
rect -3591 -151 -2583 -145
rect -1533 -111 -525 -105
rect -1533 -145 -1521 -111
rect -537 -145 -525 -111
rect -1533 -151 -525 -145
rect 525 -111 1533 -105
rect 525 -145 537 -111
rect 1521 -145 1533 -111
rect 525 -151 1533 -145
rect 2583 -111 3591 -105
rect 2583 -145 2595 -111
rect 3579 -145 3591 -111
rect 2583 -151 3591 -145
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 10 m 1 nf 4 diffcov 100 polycov 50 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
