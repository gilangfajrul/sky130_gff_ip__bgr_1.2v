magic
tech sky130A
timestamp 1716188352
<< nwell >>
rect -1176 -81 1176 81
<< pmos >>
rect -1129 -50 -629 50
rect -543 -50 -43 50
rect 43 -50 543 50
rect 629 -50 1129 50
<< pdiff >>
rect -1158 44 -1129 50
rect -1158 -44 -1152 44
rect -1135 -44 -1129 44
rect -1158 -50 -1129 -44
rect -629 44 -600 50
rect -629 -44 -623 44
rect -606 -44 -600 44
rect -629 -50 -600 -44
rect -572 44 -543 50
rect -572 -44 -566 44
rect -549 -44 -543 44
rect -572 -50 -543 -44
rect -43 44 -14 50
rect -43 -44 -37 44
rect -20 -44 -14 44
rect -43 -50 -14 -44
rect 14 44 43 50
rect 14 -44 20 44
rect 37 -44 43 44
rect 14 -50 43 -44
rect 543 44 572 50
rect 543 -44 549 44
rect 566 -44 572 44
rect 543 -50 572 -44
rect 600 44 629 50
rect 600 -44 606 44
rect 623 -44 629 44
rect 600 -50 629 -44
rect 1129 44 1158 50
rect 1129 -44 1135 44
rect 1152 -44 1158 44
rect 1129 -50 1158 -44
<< pdiffc >>
rect -1152 -44 -1135 44
rect -623 -44 -606 44
rect -566 -44 -549 44
rect -37 -44 -20 44
rect 20 -44 37 44
rect 549 -44 566 44
rect 606 -44 623 44
rect 1135 -44 1152 44
<< poly >>
rect -1129 50 -629 63
rect -543 50 -43 63
rect 43 50 543 63
rect 629 50 1129 63
rect -1129 -63 -629 -50
rect -543 -63 -43 -50
rect 43 -63 543 -50
rect 629 -63 1129 -50
<< locali >>
rect -1152 44 -1135 52
rect -1152 -52 -1135 -44
rect -623 44 -606 52
rect -623 -52 -606 -44
rect -566 44 -549 52
rect -566 -52 -549 -44
rect -37 44 -20 52
rect -37 -52 -20 -44
rect 20 44 37 52
rect 20 -52 37 -44
rect 549 44 566 52
rect 549 -52 566 -44
rect 606 44 623 52
rect 606 -52 623 -44
rect 1135 44 1152 52
rect 1135 -52 1152 -44
<< viali >>
rect -1152 -44 -1135 44
rect -623 -44 -606 44
rect -566 -44 -549 44
rect -37 -44 -20 44
rect 20 -44 37 44
rect 549 -44 566 44
rect 606 -44 623 44
rect 1135 -44 1152 44
<< metal1 >>
rect -1155 44 -1132 50
rect -1155 -44 -1152 44
rect -1135 -44 -1132 44
rect -1155 -50 -1132 -44
rect -626 44 -603 50
rect -626 -44 -623 44
rect -606 -44 -603 44
rect -626 -50 -603 -44
rect -569 44 -546 50
rect -569 -44 -566 44
rect -549 -44 -546 44
rect -569 -50 -546 -44
rect -40 44 -17 50
rect -40 -44 -37 44
rect -20 -44 -17 44
rect -40 -50 -17 -44
rect 17 44 40 50
rect 17 -44 20 44
rect 37 -44 40 44
rect 17 -50 40 -44
rect 546 44 569 50
rect 546 -44 549 44
rect 566 -44 569 44
rect 546 -50 569 -44
rect 603 44 626 50
rect 603 -44 606 44
rect 623 -44 626 44
rect 603 -50 626 -44
rect 1132 44 1155 50
rect 1132 -44 1135 44
rect 1152 -44 1155 44
rect 1132 -50 1155 -44
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 5 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
