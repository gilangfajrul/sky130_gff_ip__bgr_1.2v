magic
tech sky130A
magscale 1 2
timestamp 1717076529
<< nmos >>
rect -2000 -69 2000 131
<< ndiff >>
rect -2058 119 -2000 131
rect -2058 -57 -2046 119
rect -2012 -57 -2000 119
rect -2058 -69 -2000 -57
rect 2000 119 2058 131
rect 2000 -57 2012 119
rect 2046 -57 2058 119
rect 2000 -69 2058 -57
<< ndiffc >>
rect -2046 -57 -2012 119
rect 2012 -57 2046 119
<< poly >>
rect -2000 131 2000 157
rect -2000 -107 2000 -69
rect -2000 -124 -992 -107
rect -1008 -141 -992 -124
rect 992 -124 2000 -107
rect 992 -141 1008 -124
rect -1008 -157 1008 -141
<< polycont >>
rect -992 -141 992 -107
<< locali >>
rect -2046 119 -2012 135
rect -2046 -73 -2012 -57
rect 2012 119 2046 135
rect 2012 -73 2046 -57
rect -1008 -141 -992 -107
rect 992 -141 1008 -107
<< viali >>
rect -2046 -57 -2012 119
rect 2012 -57 2046 119
rect -992 -141 992 -107
<< metal1 >>
rect -2052 119 -2006 131
rect -2052 -57 -2046 119
rect -2012 -57 -2006 119
rect -2052 -69 -2006 -57
rect 2006 119 2052 131
rect 2006 -57 2012 119
rect 2046 -57 2052 119
rect 2006 -69 2052 -57
rect -1004 -107 1004 -101
rect -1004 -141 -992 -107
rect 992 -141 1004 -107
rect -1004 -147 1004 -141
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 20 m 1 nf 1 diffcov 100 polycov 50 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
