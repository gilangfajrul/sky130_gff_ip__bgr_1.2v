magic
tech sky130A
magscale 1 2
timestamp 1716133296
<< pwell >>
rect -4283 -937 4283 937
<< nmos >>
rect -4087 527 -2087 727
rect -2029 527 -29 727
rect 29 527 2029 727
rect 2087 527 4087 727
rect -4087 109 -2087 309
rect -2029 109 -29 309
rect 29 109 2029 309
rect 2087 109 4087 309
rect -4087 -309 -2087 -109
rect -2029 -309 -29 -109
rect 29 -309 2029 -109
rect 2087 -309 4087 -109
rect -4087 -727 -2087 -527
rect -2029 -727 -29 -527
rect 29 -727 2029 -527
rect 2087 -727 4087 -527
<< ndiff >>
rect -4145 715 -4087 727
rect -4145 539 -4133 715
rect -4099 539 -4087 715
rect -4145 527 -4087 539
rect -2087 715 -2029 727
rect -2087 539 -2075 715
rect -2041 539 -2029 715
rect -2087 527 -2029 539
rect -29 715 29 727
rect -29 539 -17 715
rect 17 539 29 715
rect -29 527 29 539
rect 2029 715 2087 727
rect 2029 539 2041 715
rect 2075 539 2087 715
rect 2029 527 2087 539
rect 4087 715 4145 727
rect 4087 539 4099 715
rect 4133 539 4145 715
rect 4087 527 4145 539
rect -4145 297 -4087 309
rect -4145 121 -4133 297
rect -4099 121 -4087 297
rect -4145 109 -4087 121
rect -2087 297 -2029 309
rect -2087 121 -2075 297
rect -2041 121 -2029 297
rect -2087 109 -2029 121
rect -29 297 29 309
rect -29 121 -17 297
rect 17 121 29 297
rect -29 109 29 121
rect 2029 297 2087 309
rect 2029 121 2041 297
rect 2075 121 2087 297
rect 2029 109 2087 121
rect 4087 297 4145 309
rect 4087 121 4099 297
rect 4133 121 4145 297
rect 4087 109 4145 121
rect -4145 -121 -4087 -109
rect -4145 -297 -4133 -121
rect -4099 -297 -4087 -121
rect -4145 -309 -4087 -297
rect -2087 -121 -2029 -109
rect -2087 -297 -2075 -121
rect -2041 -297 -2029 -121
rect -2087 -309 -2029 -297
rect -29 -121 29 -109
rect -29 -297 -17 -121
rect 17 -297 29 -121
rect -29 -309 29 -297
rect 2029 -121 2087 -109
rect 2029 -297 2041 -121
rect 2075 -297 2087 -121
rect 2029 -309 2087 -297
rect 4087 -121 4145 -109
rect 4087 -297 4099 -121
rect 4133 -297 4145 -121
rect 4087 -309 4145 -297
rect -4145 -539 -4087 -527
rect -4145 -715 -4133 -539
rect -4099 -715 -4087 -539
rect -4145 -727 -4087 -715
rect -2087 -539 -2029 -527
rect -2087 -715 -2075 -539
rect -2041 -715 -2029 -539
rect -2087 -727 -2029 -715
rect -29 -539 29 -527
rect -29 -715 -17 -539
rect 17 -715 29 -539
rect -29 -727 29 -715
rect 2029 -539 2087 -527
rect 2029 -715 2041 -539
rect 2075 -715 2087 -539
rect 2029 -727 2087 -715
rect 4087 -539 4145 -527
rect 4087 -715 4099 -539
rect 4133 -715 4145 -539
rect 4087 -727 4145 -715
<< ndiffc >>
rect -4133 539 -4099 715
rect -2075 539 -2041 715
rect -17 539 17 715
rect 2041 539 2075 715
rect 4099 539 4133 715
rect -4133 121 -4099 297
rect -2075 121 -2041 297
rect -17 121 17 297
rect 2041 121 2075 297
rect 4099 121 4133 297
rect -4133 -297 -4099 -121
rect -2075 -297 -2041 -121
rect -17 -297 17 -121
rect 2041 -297 2075 -121
rect 4099 -297 4133 -121
rect -4133 -715 -4099 -539
rect -2075 -715 -2041 -539
rect -17 -715 17 -539
rect 2041 -715 2075 -539
rect 4099 -715 4133 -539
<< psubdiff >>
rect -4247 867 -4151 901
rect 4151 867 4247 901
rect -4247 805 -4213 867
rect 4213 805 4247 867
rect -4247 -867 -4213 -805
rect 4213 -867 4247 -805
rect -4247 -901 -4151 -867
rect 4151 -901 4247 -867
<< psubdiffcont >>
rect -4151 867 4151 901
rect -4247 -805 -4213 805
rect 4213 -805 4247 805
rect -4151 -901 4151 -867
<< poly >>
rect -4087 799 -2087 815
rect -4087 765 -4071 799
rect -2103 765 -2087 799
rect -4087 727 -2087 765
rect -2029 799 -29 815
rect -2029 765 -2013 799
rect -45 765 -29 799
rect -2029 727 -29 765
rect 29 799 2029 815
rect 29 765 45 799
rect 2013 765 2029 799
rect 29 727 2029 765
rect 2087 799 4087 815
rect 2087 765 2103 799
rect 4071 765 4087 799
rect 2087 727 4087 765
rect -4087 489 -2087 527
rect -4087 455 -4071 489
rect -2103 455 -2087 489
rect -4087 439 -2087 455
rect -2029 489 -29 527
rect -2029 455 -2013 489
rect -45 455 -29 489
rect -2029 439 -29 455
rect 29 489 2029 527
rect 29 455 45 489
rect 2013 455 2029 489
rect 29 439 2029 455
rect 2087 489 4087 527
rect 2087 455 2103 489
rect 4071 455 4087 489
rect 2087 439 4087 455
rect -4087 381 -2087 397
rect -4087 347 -4071 381
rect -2103 347 -2087 381
rect -4087 309 -2087 347
rect -2029 381 -29 397
rect -2029 347 -2013 381
rect -45 347 -29 381
rect -2029 309 -29 347
rect 29 381 2029 397
rect 29 347 45 381
rect 2013 347 2029 381
rect 29 309 2029 347
rect 2087 381 4087 397
rect 2087 347 2103 381
rect 4071 347 4087 381
rect 2087 309 4087 347
rect -4087 71 -2087 109
rect -4087 37 -4071 71
rect -2103 37 -2087 71
rect -4087 21 -2087 37
rect -2029 71 -29 109
rect -2029 37 -2013 71
rect -45 37 -29 71
rect -2029 21 -29 37
rect 29 71 2029 109
rect 29 37 45 71
rect 2013 37 2029 71
rect 29 21 2029 37
rect 2087 71 4087 109
rect 2087 37 2103 71
rect 4071 37 4087 71
rect 2087 21 4087 37
rect -4087 -37 -2087 -21
rect -4087 -71 -4071 -37
rect -2103 -71 -2087 -37
rect -4087 -109 -2087 -71
rect -2029 -37 -29 -21
rect -2029 -71 -2013 -37
rect -45 -71 -29 -37
rect -2029 -109 -29 -71
rect 29 -37 2029 -21
rect 29 -71 45 -37
rect 2013 -71 2029 -37
rect 29 -109 2029 -71
rect 2087 -37 4087 -21
rect 2087 -71 2103 -37
rect 4071 -71 4087 -37
rect 2087 -109 4087 -71
rect -4087 -347 -2087 -309
rect -4087 -381 -4071 -347
rect -2103 -381 -2087 -347
rect -4087 -397 -2087 -381
rect -2029 -347 -29 -309
rect -2029 -381 -2013 -347
rect -45 -381 -29 -347
rect -2029 -397 -29 -381
rect 29 -347 2029 -309
rect 29 -381 45 -347
rect 2013 -381 2029 -347
rect 29 -397 2029 -381
rect 2087 -347 4087 -309
rect 2087 -381 2103 -347
rect 4071 -381 4087 -347
rect 2087 -397 4087 -381
rect -4087 -455 -2087 -439
rect -4087 -489 -4071 -455
rect -2103 -489 -2087 -455
rect -4087 -527 -2087 -489
rect -2029 -455 -29 -439
rect -2029 -489 -2013 -455
rect -45 -489 -29 -455
rect -2029 -527 -29 -489
rect 29 -455 2029 -439
rect 29 -489 45 -455
rect 2013 -489 2029 -455
rect 29 -527 2029 -489
rect 2087 -455 4087 -439
rect 2087 -489 2103 -455
rect 4071 -489 4087 -455
rect 2087 -527 4087 -489
rect -4087 -765 -2087 -727
rect -4087 -799 -4071 -765
rect -2103 -799 -2087 -765
rect -4087 -815 -2087 -799
rect -2029 -765 -29 -727
rect -2029 -799 -2013 -765
rect -45 -799 -29 -765
rect -2029 -815 -29 -799
rect 29 -765 2029 -727
rect 29 -799 45 -765
rect 2013 -799 2029 -765
rect 29 -815 2029 -799
rect 2087 -765 4087 -727
rect 2087 -799 2103 -765
rect 4071 -799 4087 -765
rect 2087 -815 4087 -799
<< polycont >>
rect -4071 765 -2103 799
rect -2013 765 -45 799
rect 45 765 2013 799
rect 2103 765 4071 799
rect -4071 455 -2103 489
rect -2013 455 -45 489
rect 45 455 2013 489
rect 2103 455 4071 489
rect -4071 347 -2103 381
rect -2013 347 -45 381
rect 45 347 2013 381
rect 2103 347 4071 381
rect -4071 37 -2103 71
rect -2013 37 -45 71
rect 45 37 2013 71
rect 2103 37 4071 71
rect -4071 -71 -2103 -37
rect -2013 -71 -45 -37
rect 45 -71 2013 -37
rect 2103 -71 4071 -37
rect -4071 -381 -2103 -347
rect -2013 -381 -45 -347
rect 45 -381 2013 -347
rect 2103 -381 4071 -347
rect -4071 -489 -2103 -455
rect -2013 -489 -45 -455
rect 45 -489 2013 -455
rect 2103 -489 4071 -455
rect -4071 -799 -2103 -765
rect -2013 -799 -45 -765
rect 45 -799 2013 -765
rect 2103 -799 4071 -765
<< locali >>
rect -4247 867 -4151 901
rect 4151 867 4247 901
rect -4247 805 -4213 867
rect 4213 805 4247 867
rect -4087 765 -4071 799
rect -2103 765 -2087 799
rect -2029 765 -2013 799
rect -45 765 -29 799
rect 29 765 45 799
rect 2013 765 2029 799
rect 2087 765 2103 799
rect 4071 765 4087 799
rect -4133 715 -4099 731
rect -4133 523 -4099 539
rect -2075 715 -2041 731
rect -2075 523 -2041 539
rect -17 715 17 731
rect -17 523 17 539
rect 2041 715 2075 731
rect 2041 523 2075 539
rect 4099 715 4133 731
rect 4099 523 4133 539
rect -4087 455 -4071 489
rect -2103 455 -2087 489
rect -2029 455 -2013 489
rect -45 455 -29 489
rect 29 455 45 489
rect 2013 455 2029 489
rect 2087 455 2103 489
rect 4071 455 4087 489
rect -4087 347 -4071 381
rect -2103 347 -2087 381
rect -2029 347 -2013 381
rect -45 347 -29 381
rect 29 347 45 381
rect 2013 347 2029 381
rect 2087 347 2103 381
rect 4071 347 4087 381
rect -4133 297 -4099 313
rect -4133 105 -4099 121
rect -2075 297 -2041 313
rect -2075 105 -2041 121
rect -17 297 17 313
rect -17 105 17 121
rect 2041 297 2075 313
rect 2041 105 2075 121
rect 4099 297 4133 313
rect 4099 105 4133 121
rect -4087 37 -4071 71
rect -2103 37 -2087 71
rect -2029 37 -2013 71
rect -45 37 -29 71
rect 29 37 45 71
rect 2013 37 2029 71
rect 2087 37 2103 71
rect 4071 37 4087 71
rect -4087 -71 -4071 -37
rect -2103 -71 -2087 -37
rect -2029 -71 -2013 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 2013 -71 2029 -37
rect 2087 -71 2103 -37
rect 4071 -71 4087 -37
rect -4133 -121 -4099 -105
rect -4133 -313 -4099 -297
rect -2075 -121 -2041 -105
rect -2075 -313 -2041 -297
rect -17 -121 17 -105
rect -17 -313 17 -297
rect 2041 -121 2075 -105
rect 2041 -313 2075 -297
rect 4099 -121 4133 -105
rect 4099 -313 4133 -297
rect -4087 -381 -4071 -347
rect -2103 -381 -2087 -347
rect -2029 -381 -2013 -347
rect -45 -381 -29 -347
rect 29 -381 45 -347
rect 2013 -381 2029 -347
rect 2087 -381 2103 -347
rect 4071 -381 4087 -347
rect -4087 -489 -4071 -455
rect -2103 -489 -2087 -455
rect -2029 -489 -2013 -455
rect -45 -489 -29 -455
rect 29 -489 45 -455
rect 2013 -489 2029 -455
rect 2087 -489 2103 -455
rect 4071 -489 4087 -455
rect -4133 -539 -4099 -523
rect -4133 -731 -4099 -715
rect -2075 -539 -2041 -523
rect -2075 -731 -2041 -715
rect -17 -539 17 -523
rect -17 -731 17 -715
rect 2041 -539 2075 -523
rect 2041 -731 2075 -715
rect 4099 -539 4133 -523
rect 4099 -731 4133 -715
rect -4087 -799 -4071 -765
rect -2103 -799 -2087 -765
rect -2029 -799 -2013 -765
rect -45 -799 -29 -765
rect 29 -799 45 -765
rect 2013 -799 2029 -765
rect 2087 -799 2103 -765
rect 4071 -799 4087 -765
rect -4247 -867 -4213 -805
rect 4213 -867 4247 -805
rect -4247 -901 -4151 -867
rect 4151 -901 4247 -867
<< viali >>
rect -4071 765 -2103 799
rect -2013 765 -45 799
rect 45 765 2013 799
rect 2103 765 4071 799
rect -4133 539 -4099 715
rect -2075 539 -2041 715
rect -17 539 17 715
rect 2041 539 2075 715
rect 4099 539 4133 715
rect -4071 455 -2103 489
rect -2013 455 -45 489
rect 45 455 2013 489
rect 2103 455 4071 489
rect -4071 347 -2103 381
rect -2013 347 -45 381
rect 45 347 2013 381
rect 2103 347 4071 381
rect -4133 121 -4099 297
rect -2075 121 -2041 297
rect -17 121 17 297
rect 2041 121 2075 297
rect 4099 121 4133 297
rect -4071 37 -2103 71
rect -2013 37 -45 71
rect 45 37 2013 71
rect 2103 37 4071 71
rect -4071 -71 -2103 -37
rect -2013 -71 -45 -37
rect 45 -71 2013 -37
rect 2103 -71 4071 -37
rect -4133 -297 -4099 -121
rect -2075 -297 -2041 -121
rect -17 -297 17 -121
rect 2041 -297 2075 -121
rect 4099 -297 4133 -121
rect -4071 -381 -2103 -347
rect -2013 -381 -45 -347
rect 45 -381 2013 -347
rect 2103 -381 4071 -347
rect -4071 -489 -2103 -455
rect -2013 -489 -45 -455
rect 45 -489 2013 -455
rect 2103 -489 4071 -455
rect -4133 -715 -4099 -539
rect -2075 -715 -2041 -539
rect -17 -715 17 -539
rect 2041 -715 2075 -539
rect 4099 -715 4133 -539
rect -4071 -799 -2103 -765
rect -2013 -799 -45 -765
rect 45 -799 2013 -765
rect 2103 -799 4071 -765
<< metal1 >>
rect -4083 799 -2091 805
rect -4083 765 -4071 799
rect -2103 765 -2091 799
rect -4083 759 -2091 765
rect -2025 799 -33 805
rect -2025 765 -2013 799
rect -45 765 -33 799
rect -2025 759 -33 765
rect 33 799 2025 805
rect 33 765 45 799
rect 2013 765 2025 799
rect 33 759 2025 765
rect 2091 799 4083 805
rect 2091 765 2103 799
rect 4071 765 4083 799
rect 2091 759 4083 765
rect -4139 715 -4093 727
rect -4139 539 -4133 715
rect -4099 539 -4093 715
rect -4139 527 -4093 539
rect -2081 715 -2035 727
rect -2081 539 -2075 715
rect -2041 539 -2035 715
rect -2081 527 -2035 539
rect -23 715 23 727
rect -23 539 -17 715
rect 17 539 23 715
rect -23 527 23 539
rect 2035 715 2081 727
rect 2035 539 2041 715
rect 2075 539 2081 715
rect 2035 527 2081 539
rect 4093 715 4139 727
rect 4093 539 4099 715
rect 4133 539 4139 715
rect 4093 527 4139 539
rect -4083 489 -2091 495
rect -4083 455 -4071 489
rect -2103 455 -2091 489
rect -4083 449 -2091 455
rect -2025 489 -33 495
rect -2025 455 -2013 489
rect -45 455 -33 489
rect -2025 449 -33 455
rect 33 489 2025 495
rect 33 455 45 489
rect 2013 455 2025 489
rect 33 449 2025 455
rect 2091 489 4083 495
rect 2091 455 2103 489
rect 4071 455 4083 489
rect 2091 449 4083 455
rect -4083 381 -2091 387
rect -4083 347 -4071 381
rect -2103 347 -2091 381
rect -4083 341 -2091 347
rect -2025 381 -33 387
rect -2025 347 -2013 381
rect -45 347 -33 381
rect -2025 341 -33 347
rect 33 381 2025 387
rect 33 347 45 381
rect 2013 347 2025 381
rect 33 341 2025 347
rect 2091 381 4083 387
rect 2091 347 2103 381
rect 4071 347 4083 381
rect 2091 341 4083 347
rect -4139 297 -4093 309
rect -4139 121 -4133 297
rect -4099 121 -4093 297
rect -4139 109 -4093 121
rect -2081 297 -2035 309
rect -2081 121 -2075 297
rect -2041 121 -2035 297
rect -2081 109 -2035 121
rect -23 297 23 309
rect -23 121 -17 297
rect 17 121 23 297
rect -23 109 23 121
rect 2035 297 2081 309
rect 2035 121 2041 297
rect 2075 121 2081 297
rect 2035 109 2081 121
rect 4093 297 4139 309
rect 4093 121 4099 297
rect 4133 121 4139 297
rect 4093 109 4139 121
rect -4083 71 -2091 77
rect -4083 37 -4071 71
rect -2103 37 -2091 71
rect -4083 31 -2091 37
rect -2025 71 -33 77
rect -2025 37 -2013 71
rect -45 37 -33 71
rect -2025 31 -33 37
rect 33 71 2025 77
rect 33 37 45 71
rect 2013 37 2025 71
rect 33 31 2025 37
rect 2091 71 4083 77
rect 2091 37 2103 71
rect 4071 37 4083 71
rect 2091 31 4083 37
rect -4083 -37 -2091 -31
rect -4083 -71 -4071 -37
rect -2103 -71 -2091 -37
rect -4083 -77 -2091 -71
rect -2025 -37 -33 -31
rect -2025 -71 -2013 -37
rect -45 -71 -33 -37
rect -2025 -77 -33 -71
rect 33 -37 2025 -31
rect 33 -71 45 -37
rect 2013 -71 2025 -37
rect 33 -77 2025 -71
rect 2091 -37 4083 -31
rect 2091 -71 2103 -37
rect 4071 -71 4083 -37
rect 2091 -77 4083 -71
rect -4139 -121 -4093 -109
rect -4139 -297 -4133 -121
rect -4099 -297 -4093 -121
rect -4139 -309 -4093 -297
rect -2081 -121 -2035 -109
rect -2081 -297 -2075 -121
rect -2041 -297 -2035 -121
rect -2081 -309 -2035 -297
rect -23 -121 23 -109
rect -23 -297 -17 -121
rect 17 -297 23 -121
rect -23 -309 23 -297
rect 2035 -121 2081 -109
rect 2035 -297 2041 -121
rect 2075 -297 2081 -121
rect 2035 -309 2081 -297
rect 4093 -121 4139 -109
rect 4093 -297 4099 -121
rect 4133 -297 4139 -121
rect 4093 -309 4139 -297
rect -4083 -347 -2091 -341
rect -4083 -381 -4071 -347
rect -2103 -381 -2091 -347
rect -4083 -387 -2091 -381
rect -2025 -347 -33 -341
rect -2025 -381 -2013 -347
rect -45 -381 -33 -347
rect -2025 -387 -33 -381
rect 33 -347 2025 -341
rect 33 -381 45 -347
rect 2013 -381 2025 -347
rect 33 -387 2025 -381
rect 2091 -347 4083 -341
rect 2091 -381 2103 -347
rect 4071 -381 4083 -347
rect 2091 -387 4083 -381
rect -4083 -455 -2091 -449
rect -4083 -489 -4071 -455
rect -2103 -489 -2091 -455
rect -4083 -495 -2091 -489
rect -2025 -455 -33 -449
rect -2025 -489 -2013 -455
rect -45 -489 -33 -455
rect -2025 -495 -33 -489
rect 33 -455 2025 -449
rect 33 -489 45 -455
rect 2013 -489 2025 -455
rect 33 -495 2025 -489
rect 2091 -455 4083 -449
rect 2091 -489 2103 -455
rect 4071 -489 4083 -455
rect 2091 -495 4083 -489
rect -4139 -539 -4093 -527
rect -4139 -715 -4133 -539
rect -4099 -715 -4093 -539
rect -4139 -727 -4093 -715
rect -2081 -539 -2035 -527
rect -2081 -715 -2075 -539
rect -2041 -715 -2035 -539
rect -2081 -727 -2035 -715
rect -23 -539 23 -527
rect -23 -715 -17 -539
rect 17 -715 23 -539
rect -23 -727 23 -715
rect 2035 -539 2081 -527
rect 2035 -715 2041 -539
rect 2075 -715 2081 -539
rect 2035 -727 2081 -715
rect 4093 -539 4139 -527
rect 4093 -715 4099 -539
rect 4133 -715 4139 -539
rect 4093 -727 4139 -715
rect -4083 -765 -2091 -759
rect -4083 -799 -4071 -765
rect -2103 -799 -2091 -765
rect -4083 -805 -2091 -799
rect -2025 -765 -33 -759
rect -2025 -799 -2013 -765
rect -45 -799 -33 -765
rect -2025 -805 -33 -799
rect 33 -765 2025 -759
rect 33 -799 45 -765
rect 2013 -799 2025 -765
rect 33 -805 2025 -799
rect 2091 -765 4083 -759
rect 2091 -799 2103 -765
rect 4071 -799 4083 -765
rect 2091 -805 4083 -799
<< properties >>
string FIXED_BBOX -4230 -884 4230 884
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 10 m 4 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
