magic
tech sky130A
magscale 1 2
timestamp 1717771017
<< nwell >>
rect -523 -198 523 164
<< pmos >>
rect -429 -136 -29 64
rect 29 -136 429 64
<< pdiff >>
rect -487 52 -429 64
rect -487 -124 -475 52
rect -441 -124 -429 52
rect -487 -136 -429 -124
rect -29 52 29 64
rect -29 -124 -17 52
rect 17 -124 29 52
rect -29 -136 29 -124
rect 429 52 487 64
rect 429 -124 441 52
rect 475 -124 487 52
rect 429 -136 487 -124
<< pdiffc >>
rect -475 -124 -441 52
rect -17 -124 17 52
rect 441 -124 475 52
<< poly >>
rect -337 145 -121 161
rect -337 128 -321 145
rect -429 111 -321 128
rect -137 128 -121 145
rect 121 145 337 161
rect 121 128 137 145
rect -137 111 -29 128
rect -429 64 -29 111
rect 29 111 137 128
rect 321 128 337 145
rect 321 111 429 128
rect 29 64 429 111
rect -429 -162 -29 -136
rect 29 -162 429 -136
<< polycont >>
rect -321 111 -137 145
rect 137 111 321 145
<< locali >>
rect -337 111 -321 145
rect -137 111 -121 145
rect 121 111 137 145
rect 321 111 337 145
rect -475 52 -441 68
rect -475 -140 -441 -124
rect -17 52 17 68
rect -17 -140 17 -124
rect 441 52 475 68
rect 441 -140 475 -124
<< viali >>
rect -321 111 -137 145
rect 137 111 321 145
rect -475 -124 -441 52
rect -17 -124 17 52
rect 441 -124 475 52
<< metal1 >>
rect -333 145 -125 151
rect -333 111 -321 145
rect -137 111 -125 145
rect -333 105 -125 111
rect 125 145 333 151
rect 125 111 137 145
rect 321 111 333 145
rect 125 105 333 111
rect -481 52 -435 64
rect -481 -124 -475 52
rect -441 -124 -435 52
rect -481 -136 -435 -124
rect -23 52 23 64
rect -23 -124 -17 52
rect 17 -124 23 52
rect -23 -136 23 -124
rect 435 52 481 64
rect 435 -124 441 52
rect 475 -124 481 52
rect 435 -136 481 -124
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 2 m 1 nf 2 diffcov 100 polycov 50 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
