magic
tech sky130A
magscale 1 2
timestamp 1717930986
<< nwell >>
rect -225 -1450 4471 516
<< nsubdiff >>
rect -189 446 -129 480
rect 4375 446 4435 480
rect -189 420 -155 446
rect 4401 420 4435 446
rect -189 -1380 -155 -1354
rect 4401 -1380 4435 -1354
rect -189 -1414 -129 -1380
rect 4375 -1414 4435 -1380
<< nsubdiffcont >>
rect -129 446 4375 480
rect -189 -1354 -155 420
rect 4401 -1354 4435 420
rect -129 -1414 4375 -1380
<< poly >>
rect -56 381 36 397
rect -56 347 -40 381
rect -6 347 36 381
rect -56 331 36 347
rect 6 300 36 331
rect 4210 381 4302 397
rect 4210 347 4252 381
rect 4286 347 4302 381
rect 4210 331 4302 347
rect 4210 326 4240 331
rect 6 -434 36 -332
rect -56 -450 36 -434
rect -56 -484 -40 -450
rect -6 -484 36 -450
rect -56 -500 36 -484
rect 6 -602 36 -500
rect 4210 -434 4240 -350
rect 4210 -450 4302 -434
rect 4210 -484 4252 -450
rect 4286 -484 4302 -450
rect 4210 -500 4302 -484
rect 4210 -583 4240 -500
rect 6 -1265 36 -1234
rect -56 -1281 36 -1265
rect -56 -1315 -40 -1281
rect -6 -1315 36 -1281
rect -56 -1331 36 -1315
rect 4210 -1265 4240 -1234
rect 4210 -1281 4302 -1265
rect 4210 -1315 4252 -1281
rect 4286 -1315 4302 -1281
rect 4210 -1331 4302 -1315
<< polycont >>
rect -40 347 -6 381
rect 4252 347 4286 381
rect -40 -484 -6 -450
rect 4252 -484 4286 -450
rect -40 -1315 -6 -1281
rect 4252 -1315 4286 -1281
<< locali >>
rect -189 446 -129 480
rect 4375 446 4435 480
rect -189 420 -155 446
rect 4401 420 4435 446
rect -40 381 -6 397
rect -40 300 -6 347
rect 4252 381 4286 397
rect 4252 298 4286 347
rect -40 -450 -6 -434
rect -40 -500 -6 -484
rect 4252 -450 4286 -434
rect 4252 -500 4286 -484
rect -40 -1281 -6 -1234
rect -40 -1331 -6 -1315
rect 4252 -1281 4286 -1234
rect 4252 -1331 4286 -1315
rect -189 -1380 -155 -1354
rect 4401 -1380 4435 -1354
rect -189 -1414 -129 -1380
rect 4375 -1414 4435 -1380
<< viali >>
rect 2106 446 2140 480
rect -189 347 -155 381
rect -40 347 -6 381
rect 4252 347 4286 381
rect 4401 347 4435 381
rect -189 -484 -155 -450
rect -40 -484 -6 -450
rect 4252 -484 4286 -450
rect 4401 -484 4435 -450
rect -189 -1315 -155 -1281
rect -40 -1315 -6 -1281
rect 4252 -1315 4286 -1281
rect 4401 -1315 4435 -1281
rect 2106 -1414 2140 -1380
<< metal1 >>
rect 2100 480 2146 492
rect 2100 446 2106 480
rect 2140 446 2146 480
rect -195 381 0 393
rect -195 347 -189 381
rect -155 347 -40 381
rect -6 347 0 381
rect -195 335 0 347
rect -46 300 0 335
rect 2100 288 2146 446
rect 4246 381 4441 393
rect 4246 347 4252 381
rect 4286 347 4401 381
rect 4435 347 4441 381
rect 4246 335 4441 347
rect 4246 295 4292 335
rect 2087 112 2097 288
rect 2149 112 2159 288
rect 4145 112 4155 288
rect 4207 112 4217 288
rect -150 10 -140 62
rect -88 59 -78 62
rect 42 59 88 108
rect 4324 59 4334 62
rect -88 13 4334 59
rect -88 10 -78 13
rect 4324 10 4334 13
rect 4386 10 4396 62
rect 29 -320 39 -144
rect 91 -320 101 -144
rect 2087 -320 2097 -144
rect 2149 -320 2159 -144
rect -46 -438 0 -325
rect -195 -450 0 -438
rect 590 -444 1598 -411
rect 2648 -444 3656 -412
rect 4158 -444 4204 -322
rect -195 -484 -189 -450
rect -155 -484 -40 -450
rect -6 -484 0 -450
rect -195 -496 0 -484
rect -46 -603 0 -496
rect 42 -490 4204 -444
rect 4246 -438 4292 -324
rect 4246 -450 4441 -438
rect 4246 -484 4252 -450
rect 4286 -484 4401 -450
rect 4435 -484 4441 -450
rect 42 -611 88 -490
rect 590 -518 1598 -490
rect 2648 -519 3656 -490
rect 4246 -496 4441 -484
rect 4246 -605 4292 -496
rect 2087 -790 2097 -614
rect 2149 -790 2159 -614
rect 4145 -790 4155 -614
rect 4207 -790 4217 -614
rect -150 -996 -140 -944
rect -88 -947 -78 -944
rect 4324 -947 4334 -944
rect -88 -993 740 -947
rect 1575 -993 2671 -947
rect 3624 -993 4334 -947
rect -88 -996 -78 -993
rect 4158 -1041 4204 -993
rect 4324 -996 4334 -993
rect 4386 -996 4396 -944
rect 29 -1222 39 -1046
rect 91 -1222 101 -1046
rect 2087 -1222 2097 -1046
rect 2149 -1222 2159 -1046
rect -46 -1269 0 -1234
rect -195 -1281 0 -1269
rect -195 -1315 -189 -1281
rect -155 -1315 -40 -1281
rect -6 -1315 0 -1281
rect -195 -1327 0 -1315
rect 2100 -1380 2146 -1222
rect 4246 -1269 4292 -1234
rect 4246 -1281 4441 -1269
rect 4246 -1315 4252 -1281
rect 4286 -1315 4401 -1281
rect 4435 -1315 4441 -1281
rect 4246 -1327 4441 -1315
rect 2100 -1414 2106 -1380
rect 2140 -1414 2146 -1380
rect 2100 -1426 2146 -1414
<< via1 >>
rect 2097 112 2149 288
rect 4155 112 4207 288
rect -140 10 -88 62
rect 4334 10 4386 62
rect 39 -320 91 -144
rect 2097 -320 2149 -144
rect 2097 -790 2149 -614
rect 4155 -790 4207 -614
rect -140 -996 -88 -944
rect 4334 -996 4386 -944
rect 39 -1222 91 -1046
rect 2097 -1222 2149 -1046
<< metal2 >>
rect 2097 288 2149 298
rect 2095 112 2097 152
rect -140 62 -88 72
rect -140 -944 -88 10
rect 2095 -134 2149 112
rect 4153 288 4209 298
rect 4153 102 4209 112
rect 4334 62 4386 72
rect 39 -144 91 -134
rect 39 -441 91 -320
rect 2095 -144 2151 -134
rect 2095 -330 2151 -320
rect 39 -493 4207 -441
rect 2095 -614 2151 -604
rect 2095 -800 2151 -790
rect 4155 -614 4207 -493
rect 4155 -800 4207 -790
rect -140 -1006 -88 -996
rect 37 -1046 93 -1036
rect 37 -1232 93 -1222
rect 2097 -1046 2151 -800
rect 4334 -944 4386 10
rect 4334 -1006 4386 -996
rect 2149 -1064 2151 -1046
rect 2097 -1232 2149 -1222
<< via2 >>
rect 4153 112 4155 288
rect 4155 112 4207 288
rect 4207 112 4209 288
rect 2095 -320 2097 -144
rect 2097 -320 2149 -144
rect 2149 -320 2151 -144
rect 2095 -790 2097 -614
rect 2097 -790 2149 -614
rect 2149 -790 2151 -614
rect 37 -1222 39 -1046
rect 39 -1222 91 -1046
rect 91 -1222 93 -1046
<< metal3 >>
rect 4143 288 4219 293
rect 4143 112 4153 288
rect 4209 112 4219 288
rect 4143 107 4219 112
rect 4151 26 4211 107
rect 4151 -34 4386 26
rect 2085 -144 2161 -139
rect 2081 -320 2091 -144
rect 2155 -320 2165 -144
rect 2085 -325 2161 -320
rect 4326 -437 4386 -34
rect -140 -497 4386 -437
rect -140 -900 -80 -497
rect 2085 -614 2161 -609
rect 2081 -790 2091 -614
rect 2155 -790 2165 -614
rect 2085 -795 2161 -790
rect -140 -960 95 -900
rect 35 -1041 95 -960
rect 27 -1046 103 -1041
rect 27 -1222 37 -1046
rect 93 -1222 103 -1046
rect 27 -1227 103 -1222
<< via3 >>
rect 2091 -320 2095 -144
rect 2095 -320 2151 -144
rect 2151 -320 2155 -144
rect 2091 -790 2095 -614
rect 2095 -790 2151 -614
rect 2151 -790 2155 -614
<< metal4 >>
rect 2090 -144 2156 -143
rect 2090 -320 2091 -144
rect 2155 -320 2156 -144
rect 2090 -321 2156 -320
rect 2091 -613 2155 -321
rect 2090 -614 2156 -613
rect 2090 -790 2091 -614
rect 2155 -790 2156 -614
rect 2090 -791 2156 -790
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_0
timestamp 1717765832
transform 1 0 21 0 1 -702
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_1
timestamp 1717765832
transform 1 0 4225 0 1 -1134
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_2
timestamp 1717765832
transform 1 0 4225 0 1 -702
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_3
timestamp 1717765832
transform 1 0 4225 0 1 -232
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_4
timestamp 1717765832
transform 1 0 4225 0 1 200
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_5
timestamp 1717765832
transform 1 0 21 0 1 200
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_6
timestamp 1717765832
transform 1 0 21 0 1 -232
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_7
timestamp 1717765832
transform 1 0 21 0 1 -1134
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_8RMJP2  sky130_fd_pr__pfet_01v8_8RMJP2_0
timestamp 1717765832
transform 1 0 2123 0 1 -1098
box -2123 -198 2123 164
use sky130_fd_pr__pfet_01v8_8RMJP2  sky130_fd_pr__pfet_01v8_8RMJP2_1
timestamp 1717765832
transform 1 0 2123 0 1 -666
box -2123 -198 2123 164
use sky130_fd_pr__pfet_01v8_CVRJBD  sky130_fd_pr__pfet_01v8_CVRJBD_0
timestamp 1717765832
transform 1 0 2123 0 1 -268
box -2123 -164 2123 198
use sky130_fd_pr__pfet_01v8_CVRJBD  sky130_fd_pr__pfet_01v8_CVRJBD_1
timestamp 1717765832
transform 1 0 2123 0 1 164
box -2123 -164 2123 198
<< labels >>
flabel metal1 2119 423 2119 423 1 FreeSans 160 0 0 0 vdde
port 0 n
flabel metal3 4176 73 4176 73 1 FreeSans 160 0 0 0 D3
port 1 n
flabel metal1 4048 25 4048 25 1 FreeSans 160 0 0 0 D4
port 3 n
flabel metal1 4190 -425 4190 -425 1 FreeSans 160 0 0 0 D9
port 4 n
flabel metal2 4182 -560 4182 -560 1 FreeSans 160 0 0 0 D8
port 5 n
<< end >>
