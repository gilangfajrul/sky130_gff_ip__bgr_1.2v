magic
tech sky130A
magscale 1 2
timestamp 1717596886
<< metal1 >>
rect -14 14 14 71
rect -14 -71 14 -14
<< rmetal1 >>
rect -14 -14 14 14
<< properties >>
string gencell sky130_fd_pr__res_generic_m1
string library sky130
string parameters w 0.140 l 0.140 m 1 nx 1 wmin 0.14 lmin 0.14 rho 0.125 val 125.0m dummy 0 dw 0.0 term 0.0 roverlap 0
<< end >>
