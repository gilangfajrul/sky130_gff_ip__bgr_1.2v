magic
tech sky130A
magscale 1 2
timestamp 1717511400
<< checkpaint >>
rect 15711 1523 18653 1576
rect 15711 1470 19022 1523
rect 15711 1417 19391 1470
rect 15711 -1982 19760 1417
rect 16080 -2035 19760 -1982
rect 16449 -2088 19760 -2035
rect 16818 -2141 19760 -2088
<< error_s >>
rect -287 492 -275 526
rect -253 458 -241 492
rect -204 458 -58 492
rect -4 458 3971 492
rect -343 -163 -315 458
rect -309 -95 -275 458
rect -192 428 -158 458
rect -104 428 -70 458
rect 8 428 42 458
rect -204 424 -58 428
rect -4 424 3833 428
rect -204 422 3833 424
rect -192 418 -158 422
rect -104 418 -70 422
rect 8 418 42 422
rect -185 394 76 396
rect -189 384 -36 390
rect -26 384 76 390
rect -247 266 -221 318
rect -247 118 -201 266
rect -226 114 -201 118
rect -192 227 -167 232
rect 3811 228 3869 318
rect -192 118 -158 227
rect -115 216 -70 227
rect -3 216 42 227
rect -104 118 -70 216
rect 8 118 42 216
rect 3823 130 3857 228
rect -192 114 -146 118
rect -207 80 -146 114
rect -116 80 -58 118
rect -189 46 -58 80
rect -189 30 -146 46
rect -116 30 -58 46
rect -73 28 -58 30
rect -4 80 54 118
rect 3795 80 3833 118
rect -4 46 3833 80
rect -4 30 54 46
rect -4 28 11 30
rect 54 2 3853 30
rect 3937 2 3971 458
rect 8236 439 8248 473
rect 8336 440 8364 493
rect 3937 0 3948 2
rect 3956 0 3971 2
rect -192 -28 -139 -11
rect -192 -45 0 -28
rect -173 -61 0 -45
rect -189 -62 3811 -61
rect -269 -95 -167 -78
rect 3789 -95 3891 -78
rect 3937 -95 3971 0
rect 3990 422 4112 439
rect 4166 422 8310 439
rect 8336 422 8482 440
rect 3990 416 4054 422
rect 4224 416 8224 422
rect 3990 407 4065 416
rect 4213 407 8235 416
rect 3990 405 8235 407
rect 8275 405 8310 422
rect 8348 418 8382 420
rect 8436 418 8470 420
rect 3990 -95 4024 405
rect 8276 386 8310 405
rect 8553 386 8587 1485
rect 4100 265 4150 304
rect 8276 266 8278 282
rect 8295 266 8310 386
rect 4092 254 4150 265
rect 4092 253 4134 254
rect 4092 239 4138 253
rect 4070 216 4100 232
rect 4066 40 4100 216
rect 4104 77 4138 239
rect 8150 228 8208 265
rect 4167 216 4212 227
rect 4104 61 4134 77
rect 4178 65 4212 216
rect 8162 77 8196 228
rect 4070 27 4100 40
rect 4166 28 8172 65
rect 4166 18 8134 27
rect 8242 24 8270 232
rect 4166 2 4250 18
rect 5182 -7 7266 18
rect 5216 -23 7232 -10
rect 4224 -27 8192 -23
rect 5216 -47 7232 -27
rect 5216 -50 8174 -47
rect 5216 -60 7232 -50
rect 4166 -75 8134 -61
rect 4166 -78 8146 -75
rect 4166 -81 8134 -78
rect 5194 -82 7254 -81
rect 8276 -95 8310 266
rect 8329 384 12553 386
rect 8329 352 8364 384
rect 8425 352 12553 384
rect 12614 352 12649 386
rect 8329 228 8363 352
rect 8489 250 8504 266
rect 8505 250 8520 266
rect 8493 244 8504 250
rect 8455 228 8470 232
rect 8329 28 8364 228
rect 8455 216 8482 228
rect 8436 200 8470 216
rect 8474 212 8482 216
rect 8436 40 8477 200
rect 8443 29 8477 40
rect 8329 -95 8363 28
rect 8431 27 8439 28
rect 8443 27 8483 29
rect 8489 27 8528 47
rect 8431 12 8528 27
rect 8455 -11 8470 8
rect 8489 1 8528 12
rect 8436 -14 8470 -11
rect 8455 -61 8470 -14
rect 8476 -16 8528 1
rect 8489 -48 8528 -16
rect 8553 -48 8587 352
rect 12615 333 12649 352
rect 8489 -60 8587 -48
rect 8489 -61 8528 -60
rect 8553 -76 8587 -60
rect 8553 -87 8564 -76
rect 8576 -87 8587 -76
rect 8553 -95 8587 -87
rect -309 -96 8587 -95
rect -309 -100 -201 -96
rect -200 -100 8587 -96
rect -309 -112 8587 -100
rect -309 -129 -261 -112
rect -249 -129 8587 -112
rect 3937 -378 3971 -129
rect 3956 -474 3971 -378
rect 3990 -474 4024 -129
rect 4104 -153 4138 -149
rect 8162 -153 8196 -149
rect 4092 -154 4150 -153
rect 8150 -154 8208 -153
rect 4104 -163 4138 -154
rect 8162 -163 8196 -154
rect 8276 -431 8310 -129
rect 3990 -508 4005 -474
rect 8295 -527 8310 -431
rect 8329 -527 8363 -129
rect 8489 -163 8621 -134
rect 8329 -561 8344 -527
rect 12634 -580 12649 333
rect 12668 299 12703 333
rect 16953 299 16988 333
rect 12668 -580 12702 299
rect 16954 280 16988 299
rect 12668 -614 12683 -580
rect 16973 -633 16988 280
rect 17007 246 17042 280
rect 17322 246 17357 280
rect 17007 -633 17041 246
rect 17323 227 17357 246
rect 17153 178 17211 184
rect 17153 144 17165 178
rect 17153 138 17211 144
rect 17153 -132 17211 -126
rect 17153 -166 17165 -132
rect 17153 -172 17211 -166
rect 17153 -240 17211 -234
rect 17153 -274 17165 -240
rect 17153 -280 17211 -274
rect 17153 -550 17211 -544
rect 17153 -584 17165 -550
rect 17153 -590 17211 -584
rect 17007 -667 17022 -633
rect 17342 -686 17357 227
rect 17376 193 17411 227
rect 17691 193 17726 227
rect 17376 -686 17410 193
rect 17692 174 17726 193
rect 17522 125 17580 131
rect 17522 91 17534 125
rect 17522 85 17580 91
rect 17522 -185 17580 -179
rect 17522 -219 17534 -185
rect 17522 -225 17580 -219
rect 17522 -293 17580 -287
rect 17522 -327 17534 -293
rect 17522 -333 17580 -327
rect 17522 -603 17580 -597
rect 17522 -637 17534 -603
rect 17522 -643 17580 -637
rect 17376 -720 17391 -686
rect 17711 -739 17726 174
rect 17745 140 17780 174
rect 17745 -739 17779 140
rect 17891 72 17949 78
rect 17891 38 17903 72
rect 17891 32 17949 38
rect 17891 -238 17949 -232
rect 17891 -272 17903 -238
rect 17891 -278 17949 -272
rect 17891 -346 17949 -340
rect 17891 -380 17903 -346
rect 17891 -386 17949 -380
rect 17891 -656 17949 -650
rect 17891 -690 17903 -656
rect 17891 -696 17949 -690
rect 17745 -773 17760 -739
<< psubdiff >>
rect -309 1533 -249 1567
rect 8527 1533 8587 1567
rect -309 1485 -275 1533
rect 8553 1485 8587 1533
rect -309 -95 -275 -69
rect 8553 -95 8587 -69
rect -309 -129 -249 -95
rect 8527 -129 8587 -95
<< psubdiffcont >>
rect -249 1533 8527 1567
rect -309 -69 -275 1485
rect 8553 -69 8587 1485
rect -249 -129 8527 -95
<< poly >>
rect -208 1483 -116 1499
rect -208 1449 -192 1483
rect -158 1449 -116 1483
rect -208 1433 -116 1449
rect 8394 1187 8424 1210
rect 54 1042 8224 1184
rect 8394 1171 8486 1187
rect 8394 1137 8436 1171
rect 8470 1137 8486 1171
rect 8394 1121 8486 1137
rect -146 793 -116 816
rect -208 777 -116 793
rect 8394 793 8424 816
rect -208 743 -192 777
rect -158 743 -116 777
rect -208 695 -116 743
rect -208 661 -192 695
rect -158 661 -116 695
rect -208 645 -116 661
rect 54 648 8224 790
rect 8394 777 8486 793
rect 8394 743 8436 777
rect 8470 743 8486 777
rect 8394 695 8486 743
rect 8394 661 8436 695
rect 8470 661 8486 695
rect -146 622 -116 645
rect 8394 645 8486 661
rect 8394 622 8424 645
rect 54 254 8224 396
rect -146 5 -116 28
rect -208 -11 -116 5
rect -208 -45 -192 -11
rect -158 -45 -116 -11
rect -208 -61 -116 -45
rect 8394 5 8424 28
rect 8394 -11 8486 5
rect 8394 -45 8436 -11
rect 8470 -45 8486 -11
rect 8394 -61 8486 -45
<< polycont >>
rect -192 1449 -158 1483
rect 8436 1137 8470 1171
rect -192 743 -158 777
rect -192 661 -158 695
rect 8436 743 8470 777
rect 8436 661 8470 695
rect -192 -45 -158 -11
rect 8436 -45 8470 -11
<< locali >>
rect -309 1533 -249 1567
rect 8527 1533 8587 1567
rect -309 1485 -275 1533
rect -192 1483 -158 1499
rect -192 1410 -158 1449
rect 8553 1485 8587 1533
rect 8436 1171 8470 1210
rect 8436 1121 8470 1137
rect -192 777 -158 816
rect -192 695 -158 743
rect -192 622 -158 661
rect 8436 777 8470 816
rect 8436 695 8470 743
rect 8436 622 8470 661
rect -192 -11 -158 28
rect -192 -61 -158 -45
rect 8436 -11 8470 28
rect 8436 -61 8470 -45
rect -309 -95 -275 -69
rect 8553 -95 8587 -69
rect -309 -129 -249 -95
rect 8527 -129 8587 -95
<< viali >>
rect 4066 1533 4100 1567
rect -309 1449 -275 1483
rect -192 1449 -158 1483
rect 8436 1137 8470 1171
rect 8553 1137 8587 1171
rect -309 702 -275 736
rect -192 743 -158 777
rect -192 661 -158 695
rect 8436 743 8470 777
rect 8436 661 8470 695
rect 8553 702 8587 736
rect -309 -45 -275 -11
rect -192 -45 -158 -11
rect 8436 -45 8470 -11
rect 8553 -45 8587 -11
rect 4178 -129 4212 -95
<< metal1 >>
rect 4060 1567 4106 1579
rect 4060 1533 4066 1567
rect 4100 1533 4106 1567
rect -315 1483 -152 1495
rect -315 1449 -309 1483
rect -275 1449 -192 1483
rect -158 1449 -152 1483
rect -315 1437 -152 1449
rect -198 1408 -152 1437
rect 8 1442 1089 1488
rect 8 1410 42 1442
rect -110 1210 48 1410
rect 4060 1405 4106 1533
rect 8230 1398 8388 1410
rect 4060 1016 4106 1227
rect 4153 1222 4163 1398
rect 4227 1222 4237 1398
rect 8230 1222 8283 1398
rect 8335 1222 8388 1398
rect 8230 1210 8388 1222
rect 8430 1183 8476 1210
rect 8430 1171 8593 1183
rect 8430 1137 8436 1171
rect 8470 1137 8553 1171
rect 8587 1137 8593 1171
rect 8430 1125 8593 1137
rect -110 1004 48 1016
rect -110 828 -57 1004
rect -5 828 48 1004
rect -110 816 48 828
rect -198 777 -152 816
rect -198 748 -192 777
rect -315 743 -192 748
rect -158 743 -152 777
rect -315 736 -152 743
rect -315 702 -309 736
rect -275 702 -152 736
rect -315 695 -152 702
rect -315 690 -192 695
rect -198 661 -192 690
rect -158 661 -152 695
rect -198 622 -152 661
rect -110 610 48 622
rect -110 434 -57 610
rect -5 434 48 610
rect -110 422 48 434
rect 4060 450 4217 1016
rect 8230 1004 8388 1016
rect 8230 828 8283 1004
rect 8335 828 8388 1004
rect 8230 820 8388 828
rect 8230 816 8387 820
rect 8430 777 8476 816
rect 8430 743 8436 777
rect 8470 748 8476 777
rect 8470 743 8593 748
rect 8430 736 8593 743
rect 8430 702 8553 736
rect 8587 702 8593 736
rect 8430 695 8593 702
rect 8430 661 8436 695
rect 8470 690 8593 695
rect 8470 661 8476 690
rect 8430 622 8476 661
rect 8230 610 8388 622
rect 4060 422 4218 450
rect 8230 434 8283 610
rect 8335 434 8388 610
rect 8230 422 8388 434
rect -110 216 48 228
rect 4172 216 4218 422
rect -110 40 -57 216
rect -5 40 48 216
rect 4041 40 4051 216
rect 4115 40 4125 216
rect -110 28 48 40
rect -198 1 -152 28
rect -315 -11 -152 1
rect -315 -45 -309 -11
rect -275 -45 -192 -11
rect -158 -45 -152 -11
rect -315 -57 -152 -45
rect 4172 -95 4218 40
rect 8230 28 8388 228
rect 8236 -4 8270 28
rect 7161 -50 8270 -4
rect 8430 1 8476 28
rect 8430 -11 8593 1
rect 8430 -45 8436 -11
rect 8470 -45 8553 -11
rect 8587 -45 8593 -11
rect 8430 -57 8593 -45
rect 4172 -129 4178 -95
rect 4212 -129 4218 -95
rect 4172 -141 4218 -129
<< via1 >>
rect 4163 1222 4227 1398
rect 8283 1222 8335 1398
rect -57 828 -5 1004
rect -57 434 -5 610
rect 8283 828 8335 1004
rect 8283 434 8335 610
rect -57 40 -5 216
rect 4051 40 4115 216
<< metal2 >>
rect 4163 1398 4227 1408
rect 4163 1212 4227 1222
rect 8283 1398 8335 1408
rect 8283 1139 8335 1222
rect -270 1087 8548 1139
rect -270 351 -218 1087
rect -57 1004 -5 1014
rect -57 745 -5 828
rect 8281 1004 8337 1014
rect 8281 818 8337 828
rect -57 693 8335 745
rect -59 610 -3 620
rect -59 424 -3 434
rect 8283 610 8335 693
rect 8283 424 8335 434
rect 8496 351 8548 1087
rect -270 299 8548 351
rect -57 216 -5 299
rect -57 30 -5 40
rect 4051 216 4115 226
rect 4051 30 4115 40
<< via2 >>
rect 4163 1222 4227 1398
rect 8281 828 8283 1004
rect 8283 828 8335 1004
rect 8335 828 8337 1004
rect -59 434 -57 610
rect -57 434 -5 610
rect -5 434 -3 610
rect 4051 40 4115 216
<< metal3 >>
rect 4153 1398 4237 1403
rect 4153 1222 4163 1398
rect 4227 1222 4237 1398
rect 4153 1217 4237 1222
rect 8271 1004 8347 1009
rect 8271 828 8281 1004
rect 8337 828 8347 1004
rect 8271 823 8347 828
rect 8279 749 8339 823
rect -61 689 8339 749
rect -61 615 -1 689
rect -69 610 7 615
rect -69 434 -59 610
rect -3 434 7 610
rect -69 429 7 434
rect 4041 216 4125 221
rect 4041 40 4051 216
rect 4115 40 4125 216
rect 4041 35 4125 40
<< via3 >>
rect 4163 1222 4227 1398
rect 4051 40 4115 216
<< metal4 >>
rect 4106 1398 4228 1399
rect 4106 1222 4163 1398
rect 4227 1222 4228 1398
rect 4106 1221 4228 1222
rect 4106 217 4172 1221
rect 4050 216 4172 217
rect 4050 40 4051 216
rect 4115 40 4172 216
rect 4050 39 4172 40
use sky130_fd_pr__nfet_01v8_3KF9AC  sky130_fd_pr__nfet_01v8_3KF9AC_0
timestamp 1717076529
transform 1 0 2054 0 1 1341
box -2058 -157 2058 157
use sky130_fd_pr__nfet_01v8_3YKU97  sky130_fd_pr__nfet_01v8_3YKU97_0
timestamp 1717076529
transform 1 0 6224 0 1 97
box -2058 -157 2058 157
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_0
timestamp 1717432527
transform 1 0 -131 0 1 916
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_1
timestamp 1717432527
transform 1 0 -131 0 1 1308
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_2
timestamp 1717432527
transform 1 0 -131 0 1 522
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_3
timestamp 1717432527
transform 1 0 -131 0 1 128
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_4
timestamp 1717432527
transform 1 0 8409 0 1 128
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_5
timestamp 1717432527
transform 1 0 8409 0 1 522
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_6
timestamp 1717432527
transform 1 0 8409 0 1 916
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_7
timestamp 1717432527
transform 1 0 8409 0 1 1310
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_BSRS8Q  sky130_fd_pr__nfet_01v8_BSRS8Q_0
timestamp 1717249617
transform 1 0 6224 0 1 1310
box -2058 -126 2058 126
use sky130_fd_pr__nfet_01v8_P5G96Q  sky130_fd_pr__nfet_01v8_P5G96Q_1
timestamp 1716212328
transform 1 0 2054 0 1 128
box -2058 -126 2058 126
use sky130_fd_pr__nfet_01v8_P5G96Q  sky130_fd_pr__nfet_01v8_P5G96Q_4
timestamp 1716212328
transform 1 0 6224 0 1 522
box -2058 -126 2058 126
use sky130_fd_pr__nfet_01v8_P5G96Q  sky130_fd_pr__nfet_01v8_P5G96Q_5
timestamp 1716212328
transform 1 0 2054 0 1 522
box -2058 -126 2058 126
use sky130_fd_pr__nfet_01v8_P5G96Q  sky130_fd_pr__nfet_01v8_P5G96Q_6
timestamp 1716212328
transform 1 0 6224 0 1 916
box -2058 -126 2058 126
use sky130_fd_pr__nfet_01v8_P5G96Q  sky130_fd_pr__nfet_01v8_P5G96Q_7
timestamp 1716212328
transform 1 0 2054 0 1 916
box -2058 -126 2058 126
use sky130_fd_pr__nfet_01v8_BBNS5X  XM1
timestamp 0
transform 1 0 17182 0 1 -203
box -211 -519 211 519
use sky130_fd_pr__nfet_01v8_BBNS5X  XM2
timestamp 0
transform 1 0 17551 0 1 -256
box -211 -519 211 519
use sky130_fd_pr__nfet_01v8_BBNS5X  XM3
timestamp 0
transform 1 0 17920 0 1 -309
box -211 -519 211 519
use sky130_fd_pr__nfet_01v8_BBNS5X  XM4
timestamp 0
transform 1 0 18289 0 1 -362
box -211 -519 211 519
use sky130_fd_pr__nfet_01v8_L2333Z  XM5
timestamp 0
transform 1 0 14828 0 1 -150
box -2196 -519 2196 519
use sky130_fd_pr__nfet_01v8_L2333Z  XM6
timestamp 0
transform 1 0 6150 0 1 -44
box -2196 -519 2196 519
use sky130_fd_pr__nfet_01v8_L2333Z  XM7
timestamp 0
transform 1 0 10489 0 1 -97
box -2196 -519 2196 519
use sky130_fd_pr__nfet_01v8_L2333Z  XM8
timestamp 0
transform 1 0 1811 0 1 9
box -2196 -519 2196 519
<< labels >>
flabel metal1 8516 -20 8516 -20 0 FreeSans 160 0 0 0 GND
port 4 nsew
flabel metal1 8310 134 8310 134 0 FreeSans 160 0 0 0 D2
port 3 nsew
flabel metal2 8302 652 8302 652 0 FreeSans 160 0 0 0 D3
port 2 nsew
flabel metal3 8310 784 8310 784 0 FreeSans 160 0 0 0 D4
port 1 nsew
flabel metal2 8306 1160 8306 1160 0 FreeSans 160 0 0 0 D1
port 0 nsew
flabel metal4 4136 80 4136 80 0 FreeSans 160 0 0 0 S2
port 5 nsew
<< end >>
