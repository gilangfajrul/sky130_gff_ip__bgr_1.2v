magic
tech sky130A
magscale 1 2
timestamp 1716392850
<< nwell >>
rect 1588 980 1648 986
rect 1542 978 1648 980
rect 1542 934 3160 978
rect 3112 899 3160 934
rect 34 848 168 898
rect 34 812 82 848
rect 34 810 202 812
rect 68 768 202 810
rect 34 480 82 726
rect 1542 516 1588 732
rect 1610 682 1680 732
rect 3112 730 3168 899
rect 6120 848 6238 898
rect 4648 732 4696 808
rect 6014 768 6230 812
rect 3044 684 3260 730
rect 4602 725 4696 732
rect 1612 566 1658 682
rect 3112 650 3168 684
rect 4602 682 4704 725
rect 3112 598 3239 650
rect 1608 516 1678 566
rect 3112 564 3168 598
rect 4648 566 4704 682
rect 3042 518 3258 564
rect 34 436 176 480
rect 34 400 82 436
rect 34 350 154 400
rect 3112 349 3168 518
rect 4596 516 4704 566
rect 4648 515 4704 516
rect 4648 436 4696 515
rect 6132 436 6226 480
rect 6124 350 6236 400
rect 3112 304 3140 349
<< viali >>
rect -17 1020 17 1058
rect 6267 1020 6301 1058
rect -17 190 17 228
rect 6267 190 6301 228
<< metal1 >>
rect -23 1064 23 1070
rect 6261 1064 6307 1070
rect -23 1058 135 1064
rect -23 1020 -17 1058
rect 17 1020 135 1058
rect -23 1014 135 1020
rect 1526 1014 1668 1064
rect 3063 1014 3205 1064
rect 4600 1014 4742 1064
rect 6134 1058 6307 1064
rect 6134 1020 6267 1058
rect 6301 1020 6307 1058
rect 6134 1014 6307 1020
rect -23 1008 23 1014
rect 6261 1008 6307 1014
rect 1546 934 4736 978
rect 46 848 174 898
rect 1548 848 1594 934
rect 46 812 94 848
rect 1666 847 1676 899
rect 1728 847 1738 899
rect 3010 847 3020 899
rect 3072 847 3082 899
rect 46 768 1634 812
rect 46 480 94 768
rect 130 681 140 733
rect 192 681 202 733
rect 1474 681 1484 733
rect 1536 681 1546 733
rect 1586 732 1634 768
rect 1586 682 1686 732
rect 3118 730 3166 934
rect 3202 847 3212 899
rect 3264 847 3274 899
rect 4546 847 4556 899
rect 4608 847 4618 899
rect 4690 848 4736 934
rect 6120 848 6238 898
rect 6190 812 6238 848
rect 4654 768 6238 812
rect 4654 732 4702 768
rect 3050 684 3266 730
rect 130 515 140 567
rect 192 515 202 567
rect 1474 515 1484 567
rect 1536 515 1546 567
rect 1586 566 1634 682
rect 1586 516 1684 566
rect 3118 564 3166 684
rect 4608 682 4702 732
rect 4654 566 4702 682
rect 4738 681 4748 733
rect 4800 681 4810 733
rect 6082 681 6092 733
rect 6144 681 6154 733
rect 3048 518 3264 564
rect 1586 480 1634 516
rect 46 436 1634 480
rect 46 400 94 436
rect 46 350 160 400
rect 1548 314 1594 400
rect 1666 349 1676 401
rect 1728 349 1738 401
rect 3010 349 3020 401
rect 3072 349 3082 401
rect 3118 314 3166 518
rect 4602 516 4702 566
rect 4654 480 4702 516
rect 4738 515 4748 567
rect 4800 515 4810 567
rect 6082 515 6092 567
rect 6144 515 6154 567
rect 6190 480 6238 768
rect 4654 436 6238 480
rect 3202 349 3212 401
rect 3264 349 3274 401
rect 4546 349 4556 401
rect 4608 349 4618 401
rect 6190 400 6238 436
rect 4690 314 4736 400
rect 6124 350 6238 400
rect 1548 270 4736 314
rect -23 234 23 240
rect 6261 234 6307 240
rect -23 228 143 234
rect -23 190 -17 228
rect 17 190 143 228
rect -23 184 143 190
rect 1532 184 1674 234
rect 3062 184 3204 234
rect 4604 184 4746 234
rect 6136 228 6307 234
rect 6136 190 6267 228
rect 6301 190 6307 228
rect 6136 184 6307 190
rect -23 178 23 184
rect 6261 178 6307 184
<< via1 >>
rect 1676 847 1728 899
rect 3020 847 3072 899
rect 140 681 192 733
rect 1484 681 1536 733
rect 3212 847 3264 899
rect 4556 847 4608 899
rect 140 515 192 567
rect 1484 515 1536 567
rect 4748 681 4800 733
rect 6092 681 6144 733
rect 1676 349 1728 401
rect 3020 349 3072 401
rect 4748 515 4800 567
rect 6092 515 6144 567
rect 3212 349 3264 401
rect 4556 349 4608 401
<< metal2 >>
rect 42 937 6242 989
rect 42 733 94 937
rect 1676 899 1728 909
rect 1676 837 1728 847
rect 3020 899 3072 909
rect 3212 899 3264 909
rect 3072 847 3212 899
rect 3020 837 3072 847
rect 140 733 192 743
rect 42 681 140 733
rect 42 567 94 681
rect 140 671 192 681
rect 1484 733 1536 743
rect 1536 681 1632 733
rect 1484 671 1536 681
rect 1580 650 1632 681
rect 3116 650 3168 847
rect 3212 837 3264 847
rect 4556 899 4608 909
rect 4652 899 4704 937
rect 4608 847 4704 899
rect 4556 837 4608 847
rect 4748 733 4800 743
rect 6092 733 6144 743
rect 6190 733 6242 937
rect 4652 681 4748 733
rect 4800 681 4862 733
rect 6144 681 6242 733
rect 4652 650 4704 681
rect 4748 671 4800 681
rect 6092 671 6144 681
rect 1580 598 4704 650
rect 140 567 192 577
rect 42 515 140 567
rect 42 311 94 515
rect 140 505 192 515
rect 1484 567 1536 577
rect 1580 567 1632 598
rect 1536 515 1632 567
rect 1484 505 1536 515
rect 1676 401 1728 411
rect 1676 339 1728 349
rect 3020 401 3072 411
rect 3116 401 3168 598
rect 4652 567 4704 598
rect 4748 567 4800 577
rect 4652 515 4748 567
rect 4748 505 4800 515
rect 6092 567 6144 577
rect 6190 567 6242 681
rect 6144 515 6242 567
rect 6092 505 6144 515
rect 3212 401 3264 411
rect 3072 349 3212 401
rect 3020 339 3072 349
rect 3212 339 3264 349
rect 4556 401 4608 411
rect 4608 349 4704 401
rect 4556 339 4608 349
rect 4652 311 4704 349
rect 6190 311 6242 515
rect 42 259 6242 311
use sky130_fd_pr__res_high_po_0p35_3P95YJ  sky130_fd_pr__res_high_po_0p35_3P95YJ_0
timestamp 1716392830
transform 0 1 3142 -1 0 624
box -677 -3195 677 3195
<< end >>
