magic
tech sky130A
timestamp 1717263778
<< nwell >>
rect -1090 -81 1090 81
<< pmos >>
rect -1043 -50 -43 50
rect 43 -50 1043 50
<< pdiff >>
rect -1072 44 -1043 50
rect -1072 -44 -1066 44
rect -1049 -44 -1043 44
rect -1072 -50 -1043 -44
rect -43 44 -14 50
rect -43 -44 -37 44
rect -20 -44 -14 44
rect -43 -50 -14 -44
rect 14 44 43 50
rect 14 -44 20 44
rect 37 -44 43 44
rect 14 -50 43 -44
rect 1043 44 1072 50
rect 1043 -44 1049 44
rect 1066 -44 1072 44
rect 1043 -50 1072 -44
<< pdiffc >>
rect -1066 -44 -1049 44
rect -37 -44 -20 44
rect 20 -44 37 44
rect 1049 -44 1066 44
<< poly >>
rect -1043 50 -43 63
rect 43 50 1043 63
rect -1043 -63 -43 -50
rect 43 -63 1043 -50
<< locali >>
rect -1066 44 -1049 52
rect -1066 -52 -1049 -44
rect -37 44 -20 52
rect -37 -52 -20 -44
rect 20 44 37 52
rect 20 -52 37 -44
rect 1049 44 1066 52
rect 1049 -52 1066 -44
<< viali >>
rect -1066 -44 -1049 44
rect -37 -44 -20 44
rect 20 -44 37 44
rect 1049 -44 1066 44
<< metal1 >>
rect -1069 44 -1046 50
rect -1069 -44 -1066 44
rect -1049 -44 -1046 44
rect -1069 -50 -1046 -44
rect -40 44 -17 50
rect -40 -44 -37 44
rect -20 -44 -17 44
rect -40 -50 -17 -44
rect 17 44 40 50
rect 17 -44 20 44
rect 37 -44 40 44
rect 17 -50 40 -44
rect 1046 44 1069 50
rect 1046 -44 1049 44
rect 1066 -44 1069 44
rect 1046 -50 1069 -44
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 10 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
