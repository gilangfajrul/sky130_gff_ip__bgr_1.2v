magic
tech sky130A
magscale 1 2
timestamp 1716351939
<< xpolycontact >>
rect -284 1596 -214 2028
rect -284 1092 -214 1524
rect -118 1596 -48 2028
rect -118 1092 -48 1524
rect 48 1596 118 2028
rect 48 1092 118 1524
rect 214 1596 284 2028
rect 214 1092 284 1524
rect -284 556 -214 988
rect -284 52 -214 484
rect -118 556 -48 988
rect -118 52 -48 484
rect 48 556 118 988
rect 48 52 118 484
rect 214 556 284 988
rect 214 52 284 484
rect -284 -484 -214 -52
rect -284 -988 -214 -556
rect -118 -484 -48 -52
rect -118 -988 -48 -556
rect 48 -484 118 -52
rect 48 -988 118 -556
rect 214 -484 284 -52
rect 214 -988 284 -556
rect -284 -1524 -214 -1092
rect -284 -2028 -214 -1596
rect -118 -1524 -48 -1092
rect -118 -2028 -48 -1596
rect 48 -1524 118 -1092
rect 48 -2028 118 -1596
rect 214 -1524 284 -1092
rect 214 -2028 284 -1596
<< ppolyres >>
rect -284 1524 -214 1596
rect -118 1524 -48 1596
rect 48 1524 118 1596
rect 214 1524 284 1596
rect -284 484 -214 556
rect -118 484 -48 556
rect 48 484 118 556
rect 214 484 284 556
rect -284 -556 -214 -484
rect -118 -556 -48 -484
rect 48 -556 118 -484
rect 214 -556 284 -484
rect -284 -1596 -214 -1524
rect -118 -1596 -48 -1524
rect 48 -1596 118 -1524
rect 214 -1596 284 -1524
<< viali >>
rect -268 1613 -230 2010
rect -102 1613 -64 2010
rect 64 1613 102 2010
rect 230 1613 268 2010
rect -268 1110 -230 1507
rect -102 1110 -64 1507
rect 64 1110 102 1507
rect 230 1110 268 1507
rect -268 573 -230 970
rect -102 573 -64 970
rect 64 573 102 970
rect 230 573 268 970
rect -268 70 -230 467
rect -102 70 -64 467
rect 64 70 102 467
rect 230 70 268 467
rect -268 -467 -230 -70
rect -102 -467 -64 -70
rect 64 -467 102 -70
rect 230 -467 268 -70
rect -268 -970 -230 -573
rect -102 -970 -64 -573
rect 64 -970 102 -573
rect 230 -970 268 -573
rect -268 -1507 -230 -1110
rect -102 -1507 -64 -1110
rect 64 -1507 102 -1110
rect 230 -1507 268 -1110
rect -268 -2010 -230 -1613
rect -102 -2010 -64 -1613
rect 64 -2010 102 -1613
rect 230 -2010 268 -1613
<< metal1 >>
rect -274 2010 -224 2022
rect -274 1613 -268 2010
rect -230 1613 -224 2010
rect -274 1601 -224 1613
rect -108 2010 -58 2022
rect -108 1613 -102 2010
rect -64 1613 -58 2010
rect -108 1601 -58 1613
rect 58 2010 108 2022
rect 58 1613 64 2010
rect 102 1613 108 2010
rect 58 1601 108 1613
rect 224 2010 274 2022
rect 224 1613 230 2010
rect 268 1613 274 2010
rect 224 1601 274 1613
rect -274 1507 -224 1519
rect -274 1110 -268 1507
rect -230 1110 -224 1507
rect -274 1098 -224 1110
rect -108 1507 -58 1519
rect -108 1110 -102 1507
rect -64 1110 -58 1507
rect -108 1098 -58 1110
rect 58 1507 108 1519
rect 58 1110 64 1507
rect 102 1110 108 1507
rect 58 1098 108 1110
rect 224 1507 274 1519
rect 224 1110 230 1507
rect 268 1110 274 1507
rect 224 1098 274 1110
rect -274 970 -224 982
rect -274 573 -268 970
rect -230 573 -224 970
rect -274 561 -224 573
rect -108 970 -58 982
rect -108 573 -102 970
rect -64 573 -58 970
rect -108 561 -58 573
rect 58 970 108 982
rect 58 573 64 970
rect 102 573 108 970
rect 58 561 108 573
rect 224 970 274 982
rect 224 573 230 970
rect 268 573 274 970
rect 224 561 274 573
rect -274 467 -224 479
rect -274 70 -268 467
rect -230 70 -224 467
rect -274 58 -224 70
rect -108 467 -58 479
rect -108 70 -102 467
rect -64 70 -58 467
rect -108 58 -58 70
rect 58 467 108 479
rect 58 70 64 467
rect 102 70 108 467
rect 58 58 108 70
rect 224 467 274 479
rect 224 70 230 467
rect 268 70 274 467
rect 224 58 274 70
rect -274 -70 -224 -58
rect -274 -467 -268 -70
rect -230 -467 -224 -70
rect -274 -479 -224 -467
rect -108 -70 -58 -58
rect -108 -467 -102 -70
rect -64 -467 -58 -70
rect -108 -479 -58 -467
rect 58 -70 108 -58
rect 58 -467 64 -70
rect 102 -467 108 -70
rect 58 -479 108 -467
rect 224 -70 274 -58
rect 224 -467 230 -70
rect 268 -467 274 -70
rect 224 -479 274 -467
rect -274 -573 -224 -561
rect -274 -970 -268 -573
rect -230 -970 -224 -573
rect -274 -982 -224 -970
rect -108 -573 -58 -561
rect -108 -970 -102 -573
rect -64 -970 -58 -573
rect -108 -982 -58 -970
rect 58 -573 108 -561
rect 58 -970 64 -573
rect 102 -970 108 -573
rect 58 -982 108 -970
rect 224 -573 274 -561
rect 224 -970 230 -573
rect 268 -970 274 -573
rect 224 -982 274 -970
rect -274 -1110 -224 -1098
rect -274 -1507 -268 -1110
rect -230 -1507 -224 -1110
rect -274 -1519 -224 -1507
rect -108 -1110 -58 -1098
rect -108 -1507 -102 -1110
rect -64 -1507 -58 -1110
rect -108 -1519 -58 -1507
rect 58 -1110 108 -1098
rect 58 -1507 64 -1110
rect 102 -1507 108 -1110
rect 58 -1519 108 -1507
rect 224 -1110 274 -1098
rect 224 -1507 230 -1110
rect 268 -1507 274 -1110
rect 224 -1519 274 -1507
rect -274 -1613 -224 -1601
rect -274 -2010 -268 -1613
rect -230 -2010 -224 -1613
rect -274 -2022 -224 -2010
rect -108 -1613 -58 -1601
rect -108 -2010 -102 -1613
rect -64 -2010 -58 -1613
rect -108 -2022 -58 -2010
rect 58 -1613 108 -1601
rect 58 -2010 64 -1613
rect 102 -2010 108 -1613
rect 58 -2022 108 -2010
rect 224 -1613 274 -1601
rect 224 -2010 230 -1613
rect 268 -2010 274 -1613
rect 224 -2022 274 -2010
<< properties >>
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.350 l 0.52 m 4 nx 4 wmin 0.350 lmin 0.50 rho 319.8 val 1.588k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
