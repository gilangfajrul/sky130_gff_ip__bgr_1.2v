magic
tech sky130A
magscale 1 2
timestamp 1717755416
<< pwell >>
rect -699 -13122 699 13122
<< psubdiff >>
rect -663 13052 -567 13086
rect 567 13052 663 13086
rect -663 12990 -629 13052
rect 629 12990 663 13052
rect -663 -13052 -629 -12990
rect 629 -13052 663 -12990
rect -663 -13086 -567 -13052
rect 567 -13086 663 -13052
<< psubdiffcont >>
rect -567 13052 567 13086
rect -663 -12990 -629 12990
rect 629 -12990 663 12990
rect -567 -13086 567 -13052
<< xpolycontact >>
rect -533 12524 -463 12956
rect -533 8724 -463 9156
rect -367 12524 -297 12956
rect -367 8724 -297 9156
rect -201 12524 -131 12956
rect -201 8724 -131 9156
rect -35 12524 35 12956
rect -35 8724 35 9156
rect 131 12524 201 12956
rect 131 8724 201 9156
rect 297 12524 367 12956
rect 297 8724 367 9156
rect 463 12524 533 12956
rect 463 8724 533 9156
rect -533 8188 -463 8620
rect -533 4388 -463 4820
rect -367 8188 -297 8620
rect -367 4388 -297 4820
rect -201 8188 -131 8620
rect -201 4388 -131 4820
rect -35 8188 35 8620
rect -35 4388 35 4820
rect 131 8188 201 8620
rect 131 4388 201 4820
rect 297 8188 367 8620
rect 297 4388 367 4820
rect 463 8188 533 8620
rect 463 4388 533 4820
rect -533 3852 -463 4284
rect -533 52 -463 484
rect -367 3852 -297 4284
rect -367 52 -297 484
rect -201 3852 -131 4284
rect -201 52 -131 484
rect -35 3852 35 4284
rect -35 52 35 484
rect 131 3852 201 4284
rect 131 52 201 484
rect 297 3852 367 4284
rect 297 52 367 484
rect 463 3852 533 4284
rect 463 52 533 484
rect -533 -484 -463 -52
rect -533 -4284 -463 -3852
rect -367 -484 -297 -52
rect -367 -4284 -297 -3852
rect -201 -484 -131 -52
rect -201 -4284 -131 -3852
rect -35 -484 35 -52
rect -35 -4284 35 -3852
rect 131 -484 201 -52
rect 131 -4284 201 -3852
rect 297 -484 367 -52
rect 297 -4284 367 -3852
rect 463 -484 533 -52
rect 463 -4284 533 -3852
rect -533 -4820 -463 -4388
rect -533 -8620 -463 -8188
rect -367 -4820 -297 -4388
rect -367 -8620 -297 -8188
rect -201 -4820 -131 -4388
rect -201 -8620 -131 -8188
rect -35 -4820 35 -4388
rect -35 -8620 35 -8188
rect 131 -4820 201 -4388
rect 131 -8620 201 -8188
rect 297 -4820 367 -4388
rect 297 -8620 367 -8188
rect 463 -4820 533 -4388
rect 463 -8620 533 -8188
rect -533 -9156 -463 -8724
rect -533 -12956 -463 -12524
rect -367 -9156 -297 -8724
rect -367 -12956 -297 -12524
rect -201 -9156 -131 -8724
rect -201 -12956 -131 -12524
rect -35 -9156 35 -8724
rect -35 -12956 35 -12524
rect 131 -9156 201 -8724
rect 131 -12956 201 -12524
rect 297 -9156 367 -8724
rect 297 -12956 367 -12524
rect 463 -9156 533 -8724
rect 463 -12956 533 -12524
<< ppolyres >>
rect -533 9156 -463 12524
rect -367 9156 -297 12524
rect -201 9156 -131 12524
rect -35 9156 35 12524
rect 131 9156 201 12524
rect 297 9156 367 12524
rect 463 9156 533 12524
rect -533 4820 -463 8188
rect -367 4820 -297 8188
rect -201 4820 -131 8188
rect -35 4820 35 8188
rect 131 4820 201 8188
rect 297 4820 367 8188
rect 463 4820 533 8188
rect -533 484 -463 3852
rect -367 484 -297 3852
rect -201 484 -131 3852
rect -35 484 35 3852
rect 131 484 201 3852
rect 297 484 367 3852
rect 463 484 533 3852
rect -533 -3852 -463 -484
rect -367 -3852 -297 -484
rect -201 -3852 -131 -484
rect -35 -3852 35 -484
rect 131 -3852 201 -484
rect 297 -3852 367 -484
rect 463 -3852 533 -484
rect -533 -8188 -463 -4820
rect -367 -8188 -297 -4820
rect -201 -8188 -131 -4820
rect -35 -8188 35 -4820
rect 131 -8188 201 -4820
rect 297 -8188 367 -4820
rect 463 -8188 533 -4820
rect -533 -12524 -463 -9156
rect -367 -12524 -297 -9156
rect -201 -12524 -131 -9156
rect -35 -12524 35 -9156
rect 131 -12524 201 -9156
rect 297 -12524 367 -9156
rect 463 -12524 533 -9156
<< locali >>
rect -663 13052 -567 13086
rect 567 13052 663 13086
rect -663 12990 -629 13052
rect 629 12990 663 13052
rect -663 -13052 -629 -12990
rect 629 -13052 663 -12990
rect -663 -13086 -567 -13052
rect 567 -13086 663 -13052
<< viali >>
rect -517 12541 -479 12938
rect -351 12541 -313 12938
rect -185 12541 -147 12938
rect -19 12541 19 12938
rect 147 12541 185 12938
rect 313 12541 351 12938
rect 479 12541 517 12938
rect -517 8742 -479 9139
rect -351 8742 -313 9139
rect -185 8742 -147 9139
rect -19 8742 19 9139
rect 147 8742 185 9139
rect 313 8742 351 9139
rect 479 8742 517 9139
rect -517 8205 -479 8602
rect -351 8205 -313 8602
rect -185 8205 -147 8602
rect -19 8205 19 8602
rect 147 8205 185 8602
rect 313 8205 351 8602
rect 479 8205 517 8602
rect -517 4406 -479 4803
rect -351 4406 -313 4803
rect -185 4406 -147 4803
rect -19 4406 19 4803
rect 147 4406 185 4803
rect 313 4406 351 4803
rect 479 4406 517 4803
rect -517 3869 -479 4266
rect -351 3869 -313 4266
rect -185 3869 -147 4266
rect -19 3869 19 4266
rect 147 3869 185 4266
rect 313 3869 351 4266
rect 479 3869 517 4266
rect -517 70 -479 467
rect -351 70 -313 467
rect -185 70 -147 467
rect -19 70 19 467
rect 147 70 185 467
rect 313 70 351 467
rect 479 70 517 467
rect -517 -467 -479 -70
rect -351 -467 -313 -70
rect -185 -467 -147 -70
rect -19 -467 19 -70
rect 147 -467 185 -70
rect 313 -467 351 -70
rect 479 -467 517 -70
rect -517 -4266 -479 -3869
rect -351 -4266 -313 -3869
rect -185 -4266 -147 -3869
rect -19 -4266 19 -3869
rect 147 -4266 185 -3869
rect 313 -4266 351 -3869
rect 479 -4266 517 -3869
rect -517 -4803 -479 -4406
rect -351 -4803 -313 -4406
rect -185 -4803 -147 -4406
rect -19 -4803 19 -4406
rect 147 -4803 185 -4406
rect 313 -4803 351 -4406
rect 479 -4803 517 -4406
rect -517 -8602 -479 -8205
rect -351 -8602 -313 -8205
rect -185 -8602 -147 -8205
rect -19 -8602 19 -8205
rect 147 -8602 185 -8205
rect 313 -8602 351 -8205
rect 479 -8602 517 -8205
rect -517 -9139 -479 -8742
rect -351 -9139 -313 -8742
rect -185 -9139 -147 -8742
rect -19 -9139 19 -8742
rect 147 -9139 185 -8742
rect 313 -9139 351 -8742
rect 479 -9139 517 -8742
rect -517 -12938 -479 -12541
rect -351 -12938 -313 -12541
rect -185 -12938 -147 -12541
rect -19 -12938 19 -12541
rect 147 -12938 185 -12541
rect 313 -12938 351 -12541
rect 479 -12938 517 -12541
<< metal1 >>
rect -523 12938 -473 12950
rect -523 12541 -517 12938
rect -479 12541 -473 12938
rect -523 12529 -473 12541
rect -357 12938 -307 12950
rect -357 12541 -351 12938
rect -313 12541 -307 12938
rect -357 12529 -307 12541
rect -191 12938 -141 12950
rect -191 12541 -185 12938
rect -147 12541 -141 12938
rect -191 12529 -141 12541
rect -25 12938 25 12950
rect -25 12541 -19 12938
rect 19 12541 25 12938
rect -25 12529 25 12541
rect 141 12938 191 12950
rect 141 12541 147 12938
rect 185 12541 191 12938
rect 141 12529 191 12541
rect 307 12938 357 12950
rect 307 12541 313 12938
rect 351 12541 357 12938
rect 307 12529 357 12541
rect 473 12938 523 12950
rect 473 12541 479 12938
rect 517 12541 523 12938
rect 473 12529 523 12541
rect -523 9139 -473 9151
rect -523 8742 -517 9139
rect -479 8742 -473 9139
rect -523 8730 -473 8742
rect -357 9139 -307 9151
rect -357 8742 -351 9139
rect -313 8742 -307 9139
rect -357 8730 -307 8742
rect -191 9139 -141 9151
rect -191 8742 -185 9139
rect -147 8742 -141 9139
rect -191 8730 -141 8742
rect -25 9139 25 9151
rect -25 8742 -19 9139
rect 19 8742 25 9139
rect -25 8730 25 8742
rect 141 9139 191 9151
rect 141 8742 147 9139
rect 185 8742 191 9139
rect 141 8730 191 8742
rect 307 9139 357 9151
rect 307 8742 313 9139
rect 351 8742 357 9139
rect 307 8730 357 8742
rect 473 9139 523 9151
rect 473 8742 479 9139
rect 517 8742 523 9139
rect 473 8730 523 8742
rect -523 8602 -473 8614
rect -523 8205 -517 8602
rect -479 8205 -473 8602
rect -523 8193 -473 8205
rect -357 8602 -307 8614
rect -357 8205 -351 8602
rect -313 8205 -307 8602
rect -357 8193 -307 8205
rect -191 8602 -141 8614
rect -191 8205 -185 8602
rect -147 8205 -141 8602
rect -191 8193 -141 8205
rect -25 8602 25 8614
rect -25 8205 -19 8602
rect 19 8205 25 8602
rect -25 8193 25 8205
rect 141 8602 191 8614
rect 141 8205 147 8602
rect 185 8205 191 8602
rect 141 8193 191 8205
rect 307 8602 357 8614
rect 307 8205 313 8602
rect 351 8205 357 8602
rect 307 8193 357 8205
rect 473 8602 523 8614
rect 473 8205 479 8602
rect 517 8205 523 8602
rect 473 8193 523 8205
rect -523 4803 -473 4815
rect -523 4406 -517 4803
rect -479 4406 -473 4803
rect -523 4394 -473 4406
rect -357 4803 -307 4815
rect -357 4406 -351 4803
rect -313 4406 -307 4803
rect -357 4394 -307 4406
rect -191 4803 -141 4815
rect -191 4406 -185 4803
rect -147 4406 -141 4803
rect -191 4394 -141 4406
rect -25 4803 25 4815
rect -25 4406 -19 4803
rect 19 4406 25 4803
rect -25 4394 25 4406
rect 141 4803 191 4815
rect 141 4406 147 4803
rect 185 4406 191 4803
rect 141 4394 191 4406
rect 307 4803 357 4815
rect 307 4406 313 4803
rect 351 4406 357 4803
rect 307 4394 357 4406
rect 473 4803 523 4815
rect 473 4406 479 4803
rect 517 4406 523 4803
rect 473 4394 523 4406
rect -523 4266 -473 4278
rect -523 3869 -517 4266
rect -479 3869 -473 4266
rect -523 3857 -473 3869
rect -357 4266 -307 4278
rect -357 3869 -351 4266
rect -313 3869 -307 4266
rect -357 3857 -307 3869
rect -191 4266 -141 4278
rect -191 3869 -185 4266
rect -147 3869 -141 4266
rect -191 3857 -141 3869
rect -25 4266 25 4278
rect -25 3869 -19 4266
rect 19 3869 25 4266
rect -25 3857 25 3869
rect 141 4266 191 4278
rect 141 3869 147 4266
rect 185 3869 191 4266
rect 141 3857 191 3869
rect 307 4266 357 4278
rect 307 3869 313 4266
rect 351 3869 357 4266
rect 307 3857 357 3869
rect 473 4266 523 4278
rect 473 3869 479 4266
rect 517 3869 523 4266
rect 473 3857 523 3869
rect -523 467 -473 479
rect -523 70 -517 467
rect -479 70 -473 467
rect -523 58 -473 70
rect -357 467 -307 479
rect -357 70 -351 467
rect -313 70 -307 467
rect -357 58 -307 70
rect -191 467 -141 479
rect -191 70 -185 467
rect -147 70 -141 467
rect -191 58 -141 70
rect -25 467 25 479
rect -25 70 -19 467
rect 19 70 25 467
rect -25 58 25 70
rect 141 467 191 479
rect 141 70 147 467
rect 185 70 191 467
rect 141 58 191 70
rect 307 467 357 479
rect 307 70 313 467
rect 351 70 357 467
rect 307 58 357 70
rect 473 467 523 479
rect 473 70 479 467
rect 517 70 523 467
rect 473 58 523 70
rect -523 -70 -473 -58
rect -523 -467 -517 -70
rect -479 -467 -473 -70
rect -523 -479 -473 -467
rect -357 -70 -307 -58
rect -357 -467 -351 -70
rect -313 -467 -307 -70
rect -357 -479 -307 -467
rect -191 -70 -141 -58
rect -191 -467 -185 -70
rect -147 -467 -141 -70
rect -191 -479 -141 -467
rect -25 -70 25 -58
rect -25 -467 -19 -70
rect 19 -467 25 -70
rect -25 -479 25 -467
rect 141 -70 191 -58
rect 141 -467 147 -70
rect 185 -467 191 -70
rect 141 -479 191 -467
rect 307 -70 357 -58
rect 307 -467 313 -70
rect 351 -467 357 -70
rect 307 -479 357 -467
rect 473 -70 523 -58
rect 473 -467 479 -70
rect 517 -467 523 -70
rect 473 -479 523 -467
rect -523 -3869 -473 -3857
rect -523 -4266 -517 -3869
rect -479 -4266 -473 -3869
rect -523 -4278 -473 -4266
rect -357 -3869 -307 -3857
rect -357 -4266 -351 -3869
rect -313 -4266 -307 -3869
rect -357 -4278 -307 -4266
rect -191 -3869 -141 -3857
rect -191 -4266 -185 -3869
rect -147 -4266 -141 -3869
rect -191 -4278 -141 -4266
rect -25 -3869 25 -3857
rect -25 -4266 -19 -3869
rect 19 -4266 25 -3869
rect -25 -4278 25 -4266
rect 141 -3869 191 -3857
rect 141 -4266 147 -3869
rect 185 -4266 191 -3869
rect 141 -4278 191 -4266
rect 307 -3869 357 -3857
rect 307 -4266 313 -3869
rect 351 -4266 357 -3869
rect 307 -4278 357 -4266
rect 473 -3869 523 -3857
rect 473 -4266 479 -3869
rect 517 -4266 523 -3869
rect 473 -4278 523 -4266
rect -523 -4406 -473 -4394
rect -523 -4803 -517 -4406
rect -479 -4803 -473 -4406
rect -523 -4815 -473 -4803
rect -357 -4406 -307 -4394
rect -357 -4803 -351 -4406
rect -313 -4803 -307 -4406
rect -357 -4815 -307 -4803
rect -191 -4406 -141 -4394
rect -191 -4803 -185 -4406
rect -147 -4803 -141 -4406
rect -191 -4815 -141 -4803
rect -25 -4406 25 -4394
rect -25 -4803 -19 -4406
rect 19 -4803 25 -4406
rect -25 -4815 25 -4803
rect 141 -4406 191 -4394
rect 141 -4803 147 -4406
rect 185 -4803 191 -4406
rect 141 -4815 191 -4803
rect 307 -4406 357 -4394
rect 307 -4803 313 -4406
rect 351 -4803 357 -4406
rect 307 -4815 357 -4803
rect 473 -4406 523 -4394
rect 473 -4803 479 -4406
rect 517 -4803 523 -4406
rect 473 -4815 523 -4803
rect -523 -8205 -473 -8193
rect -523 -8602 -517 -8205
rect -479 -8602 -473 -8205
rect -523 -8614 -473 -8602
rect -357 -8205 -307 -8193
rect -357 -8602 -351 -8205
rect -313 -8602 -307 -8205
rect -357 -8614 -307 -8602
rect -191 -8205 -141 -8193
rect -191 -8602 -185 -8205
rect -147 -8602 -141 -8205
rect -191 -8614 -141 -8602
rect -25 -8205 25 -8193
rect -25 -8602 -19 -8205
rect 19 -8602 25 -8205
rect -25 -8614 25 -8602
rect 141 -8205 191 -8193
rect 141 -8602 147 -8205
rect 185 -8602 191 -8205
rect 141 -8614 191 -8602
rect 307 -8205 357 -8193
rect 307 -8602 313 -8205
rect 351 -8602 357 -8205
rect 307 -8614 357 -8602
rect 473 -8205 523 -8193
rect 473 -8602 479 -8205
rect 517 -8602 523 -8205
rect 473 -8614 523 -8602
rect -523 -8742 -473 -8730
rect -523 -9139 -517 -8742
rect -479 -9139 -473 -8742
rect -523 -9151 -473 -9139
rect -357 -8742 -307 -8730
rect -357 -9139 -351 -8742
rect -313 -9139 -307 -8742
rect -357 -9151 -307 -9139
rect -191 -8742 -141 -8730
rect -191 -9139 -185 -8742
rect -147 -9139 -141 -8742
rect -191 -9151 -141 -9139
rect -25 -8742 25 -8730
rect -25 -9139 -19 -8742
rect 19 -9139 25 -8742
rect -25 -9151 25 -9139
rect 141 -8742 191 -8730
rect 141 -9139 147 -8742
rect 185 -9139 191 -8742
rect 141 -9151 191 -9139
rect 307 -8742 357 -8730
rect 307 -9139 313 -8742
rect 351 -9139 357 -8742
rect 307 -9151 357 -9139
rect 473 -8742 523 -8730
rect 473 -9139 479 -8742
rect 517 -9139 523 -8742
rect 473 -9151 523 -9139
rect -523 -12541 -473 -12529
rect -523 -12938 -517 -12541
rect -479 -12938 -473 -12541
rect -523 -12950 -473 -12938
rect -357 -12541 -307 -12529
rect -357 -12938 -351 -12541
rect -313 -12938 -307 -12541
rect -357 -12950 -307 -12938
rect -191 -12541 -141 -12529
rect -191 -12938 -185 -12541
rect -147 -12938 -141 -12541
rect -191 -12950 -141 -12938
rect -25 -12541 25 -12529
rect -25 -12938 -19 -12541
rect 19 -12938 25 -12541
rect -25 -12950 25 -12938
rect 141 -12541 191 -12529
rect 141 -12938 147 -12541
rect 185 -12938 191 -12541
rect 141 -12950 191 -12938
rect 307 -12541 357 -12529
rect 307 -12938 313 -12541
rect 351 -12938 357 -12541
rect 307 -12950 357 -12938
rect 473 -12541 523 -12529
rect 473 -12938 479 -12541
rect 517 -12938 523 -12541
rect 473 -12950 523 -12938
<< properties >>
string FIXED_BBOX -646 -13069 646 13069
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.350 l 17 m 6 nx 7 wmin 0.350 lmin 0.50 rho 319.8 val 16.646k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
