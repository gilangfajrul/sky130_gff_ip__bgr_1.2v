magic
tech sky130A
magscale 1 2
timestamp 1762705629
<< nwell >>
rect -172 -89 4426 929
<< nsubdiff >>
rect -136 859 -76 893
rect 4330 859 4390 893
rect -136 833 -102 859
rect 4356 833 4390 859
rect -136 -19 -102 7
rect 4356 -19 4390 7
rect -136 -53 -76 -19
rect 4330 -53 4390 -19
<< nsubdiffcont >>
rect -76 859 4330 893
rect -136 7 -102 833
rect 4356 7 4390 833
rect -76 -53 4330 -19
<< poly >>
rect -26 819 40 835
rect -26 785 -10 819
rect 24 785 40 819
rect -26 769 40 785
rect 10 756 40 769
rect 4214 819 4280 835
rect 4214 785 4230 819
rect 4264 785 4280 819
rect 4214 769 4280 785
rect 4214 738 4244 769
rect 10 71 40 93
rect -26 55 40 71
rect -26 21 -10 55
rect 24 21 40 55
rect -26 5 40 21
rect 4214 71 4244 102
rect 4214 55 4280 71
rect 4214 21 4230 55
rect 4264 21 4280 55
rect 4214 5 4280 21
<< polycont >>
rect -10 785 24 819
rect 4230 785 4264 819
rect -10 21 24 55
rect 4230 21 4264 55
<< locali >>
rect -26 785 -10 819
rect 24 785 40 819
rect 4214 785 4230 819
rect 4264 785 4280 819
rect -26 21 -10 55
rect 24 21 40 55
rect 4214 21 4230 55
rect 4264 21 4280 55
<< viali >>
rect -136 859 -76 893
rect -76 859 4330 893
rect 4330 859 4390 893
rect -136 833 -102 859
rect -136 7 -102 833
rect 4356 833 4390 859
rect -10 785 24 819
rect 4230 785 4264 819
rect -10 21 24 55
rect 4230 21 4264 55
rect -136 -19 -102 7
rect 4356 7 4390 833
rect 4356 -19 4390 7
rect -136 -53 -76 -19
rect -76 -53 4330 -19
rect 4330 -53 4390 -19
<< metal1 >>
rect -142 899 -96 905
rect 4350 899 4396 905
rect -148 893 4402 899
rect -148 853 -136 893
rect -142 -13 -136 853
rect -148 -53 -136 -13
rect -102 853 4356 859
rect -102 -13 -96 853
rect -42 819 40 825
rect -42 785 -10 819
rect 24 785 40 819
rect -42 779 40 785
rect 2074 779 2172 825
rect 4214 819 4296 825
rect 4214 785 4230 819
rect 4264 785 4296 819
rect 4214 779 4296 785
rect -42 731 4 779
rect 4250 738 4296 779
rect -24 550 43 726
rect 95 550 105 726
rect 2091 550 2101 726
rect 2153 550 2163 726
rect 4149 550 4159 726
rect 4211 550 4268 726
rect 102 343 148 480
rect 2082 343 2172 497
rect 4106 343 4152 480
rect -42 114 43 290
rect 95 114 105 290
rect 2091 114 2101 290
rect 2153 114 2163 290
rect 4149 114 4159 290
rect 4211 114 4281 290
rect -42 61 4 114
rect 4250 61 4296 102
rect -42 55 40 61
rect -42 21 -10 55
rect 24 21 40 55
rect -42 15 40 21
rect 2084 15 2182 61
rect 4214 55 4296 61
rect 4214 21 4230 55
rect 4264 21 4296 55
rect 4214 15 4296 21
rect 4350 -13 4356 853
rect -102 -19 4356 -13
rect 4390 853 4402 893
rect 4390 -13 4396 853
rect 4390 -53 4402 -13
rect -148 -59 2101 -53
rect -142 -65 -96 -59
rect 2095 -81 2101 -59
rect 2153 -59 4402 -53
rect 2153 -81 2159 -59
rect 4350 -65 4396 -59
<< via1 >>
rect 43 550 95 726
rect 2101 550 2153 726
rect 4159 550 4211 726
rect 43 114 95 290
rect 2101 114 2153 290
rect 4159 114 4211 290
rect 2101 -53 2153 -29
rect 2101 -81 2153 -53
<< metal2 >>
rect 43 726 95 736
rect 43 448 95 550
rect 2101 726 2153 736
rect 32 392 41 448
rect 97 392 106 448
rect 43 290 95 392
rect 43 104 95 114
rect 2101 290 2153 550
rect 4159 726 4211 736
rect 4159 448 4211 550
rect 4148 392 4157 448
rect 4213 392 4222 448
rect 2101 -29 2153 114
rect 4159 290 4211 392
rect 4159 104 4211 114
rect 2101 -87 2153 -81
<< via2 >>
rect 41 392 97 448
rect 4157 392 4213 448
<< metal3 >>
rect 36 450 102 453
rect 4152 450 4218 453
rect 36 448 4218 450
rect 36 392 41 448
rect 97 392 4157 448
rect 4213 392 4218 448
rect 36 390 4218 392
rect 36 387 102 390
rect 4152 387 4218 390
use sky130_fd_pr__pfet_01v8_LDV24K  sky130_fd_pr__pfet_01v8_LDV24K_0
timestamp 1762704772
transform 1 0 2127 0 1 420
box -2123 -418 2123 418
use sky130_fd_pr__pfet_01v8_P4G5X4  sky130_fd_pr__pfet_01v8_P4G5X4_0
timestamp 1762704772
transform 1 0 4229 0 1 638
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_P4G5X4  sky130_fd_pr__pfet_01v8_P4G5X4_1
timestamp 1762704772
transform 1 0 4229 0 1 202
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_P4G5X4  sky130_fd_pr__pfet_01v8_P4G5X4_2
timestamp 1762704772
transform 1 0 25 0 1 202
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_P4G5X4  sky130_fd_pr__pfet_01v8_P4G5X4_3
timestamp 1762704772
transform 1 0 25 0 1 638
box -109 -162 109 162
<< labels >>
rlabel polycont 7 38 7 38 0 G
port 2 nsew
rlabel polycont 7 802 7 802 0 G
port 2 nsew
rlabel polycont 4247 38 4247 38 0 G
port 2 nsew
rlabel polycont 4247 802 4247 802 0 G
port 2 nsew
flabel metal2 2133 519 2133 519 0 FreeSans 160 0 0 0 vdde
port 3 nsew
flabel metal2 4185 341 4185 341 0 FreeSans 160 0 0 0 d10
port 0 nsew
flabel metal1 2120 797 2120 797 0 FreeSans 160 0 0 0 g10
port 1 nsew
<< end >>
