magic
tech sky130A
magscale 1 2
timestamp 1717913728
<< error_p >>
rect 19 472 77 478
rect 19 438 31 472
rect 19 432 77 438
rect -77 -438 -19 -432
rect -77 -472 -65 -438
rect -77 -478 -19 -472
<< nmos >>
rect -63 -400 -33 400
rect 33 -400 63 400
<< ndiff >>
rect -125 388 -63 400
rect -125 -388 -113 388
rect -79 -388 -63 388
rect -125 -400 -63 -388
rect -33 388 33 400
rect -33 -388 -17 388
rect 17 -388 33 388
rect -33 -400 33 -388
rect 63 388 125 400
rect 63 -388 79 388
rect 113 -388 125 388
rect 63 -400 125 -388
<< ndiffc >>
rect -113 -388 -79 388
rect -17 -388 17 388
rect 79 -388 113 388
<< poly >>
rect 15 472 81 488
rect 15 438 31 472
rect 65 438 81 472
rect -63 400 -33 426
rect 15 422 81 438
rect 33 400 63 422
rect -63 -422 -33 -400
rect -81 -438 -15 -422
rect 33 -426 63 -400
rect -81 -472 -65 -438
rect -31 -472 -15 -438
rect -81 -488 -15 -472
<< polycont >>
rect 31 438 65 472
rect -65 -472 -31 -438
<< locali >>
rect 15 438 31 472
rect 65 438 81 472
rect -113 388 -79 404
rect -113 -404 -79 -388
rect -17 388 17 404
rect -17 -404 17 -388
rect 79 388 113 404
rect 79 -404 113 -388
rect -81 -472 -65 -438
rect -31 -472 -15 -438
<< viali >>
rect 31 438 65 472
rect -113 -388 -79 388
rect -17 -388 17 388
rect 79 -388 113 388
rect -65 -472 -31 -438
<< metal1 >>
rect 19 472 77 478
rect 19 438 31 472
rect 65 438 77 472
rect 19 432 77 438
rect -119 388 -73 400
rect -119 -388 -113 388
rect -79 -388 -73 388
rect -119 -400 -73 -388
rect -23 388 23 400
rect -23 -388 -17 388
rect 17 -388 23 388
rect -23 -400 23 -388
rect 73 388 119 400
rect 73 -388 79 388
rect 113 -388 119 388
rect 73 -400 119 -388
rect -77 -438 -19 -432
rect -77 -472 -65 -438
rect -31 -472 -19 -438
rect -77 -478 -19 -472
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 4 l 0.15 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
