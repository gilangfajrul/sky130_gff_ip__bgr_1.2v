magic
tech sky130A
magscale 1 2
timestamp 1762874782
<< nwell >>
rect 3592 10722 3989 10968
rect 3535 10493 3989 10722
rect 3553 10488 3989 10493
rect 3592 10433 3989 10488
rect 3528 9950 3989 10433
<< metal1 >>
rect 4043 11080 4053 11256
rect 4105 11080 4115 11256
rect 3456 10481 3462 10484
rect 3305 10435 3462 10481
rect 3456 10432 3462 10435
rect 3514 10432 3520 10484
rect 3954 10178 3964 10354
rect 4016 10178 4026 10354
rect 3491 9980 3952 10026
rect -1283 9945 -1231 9951
rect -1283 9114 -1231 9893
rect 3228 9917 3280 9923
rect 3964 9917 4016 9923
rect 3280 9865 3964 9917
rect 3228 9859 3280 9865
rect 3964 9859 4016 9865
rect 3063 9781 3069 9833
rect 3121 9830 3127 9833
rect 8162 9830 8168 9833
rect 3121 9784 8168 9830
rect 3121 9781 3127 9784
rect 8162 9781 8168 9784
rect 8220 9781 8226 9833
rect 3331 9695 3337 9755
rect 3397 9695 3554 9755
rect 3614 9751 4110 9755
rect 3614 9699 4052 9751
rect 4104 9699 4110 9751
rect 3614 9695 4110 9699
rect 3657 9584 3663 9640
rect 3719 9584 3765 9640
rect 3821 9584 3827 9640
rect -841 9063 -718 9114
rect -1283 9056 -1231 9062
rect 5937 9057 5973 9076
rect 2613 8981 2623 9033
rect 2675 8981 2685 9033
rect 6313 8714 6323 8870
rect 6375 8714 6385 8870
rect 2973 8579 3458 8649
rect 4317 8542 4327 8594
rect 4379 8542 4389 8594
rect 8048 8514 8100 8520
rect 3222 8462 3228 8514
rect 3280 8462 8048 8514
rect 8048 8456 8100 8462
rect 3934 8422 3986 8428
rect 2880 8370 2886 8422
rect 2938 8370 3934 8422
rect 3934 8364 3986 8370
rect 6308 8368 6318 8428
rect 6380 8368 8390 8428
rect 8450 8368 8456 8428
rect 4317 8244 4327 8296
rect 4379 8244 4389 8296
rect 3059 8208 3069 8211
rect 2798 8162 3069 8208
rect 3059 8159 3069 8162
rect 3121 8159 3131 8211
<< via1 >>
rect 4053 11080 4105 11256
rect 3462 10432 3514 10484
rect 3964 10178 4016 10354
rect -1283 9893 -1231 9945
rect 3228 9865 3280 9917
rect 3964 9865 4016 9917
rect 3069 9781 3121 9833
rect 8168 9781 8220 9833
rect 3337 9695 3397 9755
rect 3554 9695 3614 9755
rect 4052 9699 4104 9751
rect 3663 9584 3719 9640
rect 3765 9584 3821 9640
rect -1283 9062 -1231 9114
rect 2623 8981 2675 9033
rect 6323 8714 6375 8870
rect 4327 8542 4379 8594
rect 3228 8462 3280 8514
rect 8048 8462 8100 8514
rect 2886 8370 2938 8422
rect 3934 8370 3986 8422
rect 6318 8368 6380 8428
rect 8390 8368 8450 8428
rect 4327 8244 4379 8296
rect 3069 8159 3121 8211
<< metal2 >>
rect 4053 11256 4105 11266
rect 3765 11123 4053 11179
rect 3462 10488 3514 10490
rect 3462 10484 3614 10488
rect 3514 10432 3614 10484
rect 3462 10428 3614 10432
rect 3462 10426 3514 10428
rect -1285 9947 -1229 9957
rect -1289 9893 -1285 9945
rect -1229 9893 -1225 9945
rect -1285 9881 -1229 9891
rect 3222 9865 3228 9917
rect 3280 9865 3286 9917
rect 3069 9833 3121 9839
rect 3069 9775 3121 9781
rect -1289 9062 -1283 9114
rect -1231 9062 -722 9114
rect 2621 9035 2677 9045
rect 2621 8969 2677 8979
rect 2886 8422 2938 8879
rect 2886 8364 2938 8370
rect 3072 8221 3118 9775
rect 3228 8514 3280 9865
rect 3337 9755 3397 9761
rect 3337 9035 3397 9695
rect 3554 9755 3614 10428
rect 3554 9685 3614 9695
rect 3663 9640 3719 9646
rect 3663 9263 3719 9584
rect 3765 9640 3821 11123
rect 4053 11070 4105 11080
rect 3964 10354 4016 10364
rect 3964 9917 4016 10178
rect 3958 9865 3964 9917
rect 4016 9865 4022 9917
rect 4052 9751 4104 10872
rect 8171 9839 8217 10205
rect 8168 9833 8220 9839
rect 8168 9775 8220 9781
rect 4052 9693 4104 9699
rect 3765 9578 3821 9584
rect 6555 9059 6578 9073
rect 3330 8979 3339 9035
rect 3395 8979 3404 9035
rect 3337 8977 3397 8979
rect 6319 8870 6379 8882
rect 6319 8714 6323 8870
rect 6375 8714 6379 8870
rect 3228 8456 3280 8462
rect 4327 8594 4379 8604
rect 3928 8370 3934 8422
rect 3986 8370 3992 8422
rect 3069 8211 3121 8221
rect 3069 8149 3121 8159
rect 3934 8072 3986 8370
rect 4327 8296 4379 8542
rect 6319 8438 6379 8714
rect 8042 8462 8048 8514
rect 8100 8462 8106 8514
rect 6318 8428 6380 8438
rect 6318 8358 6380 8368
rect 4327 8234 4379 8244
rect 8048 7838 8100 8462
rect 8390 8428 8450 8434
rect -294 7724 -238 7734
rect -294 7538 -238 7548
rect 8390 7467 8450 8368
rect 8390 7411 8392 7467
rect 8448 7411 8450 7467
rect 8390 7409 8450 7411
rect 8392 7402 8448 7409
<< via2 >>
rect -1285 9945 -1229 9947
rect -1285 9893 -1283 9945
rect -1283 9893 -1231 9945
rect -1231 9893 -1229 9945
rect -1285 9891 -1229 9893
rect 2621 9033 2677 9035
rect 2621 8981 2623 9033
rect 2623 8981 2675 9033
rect 2675 8981 2677 9033
rect 2621 8979 2677 8981
rect 3339 8979 3395 9035
rect -294 7548 -238 7724
rect 8392 7411 8448 7467
<< metal3 >>
rect -1553 10429 -605 10489
rect -1305 9952 -1205 9969
rect -1305 9886 -1290 9952
rect -1226 9886 -1205 9952
rect -1305 9869 -1205 9886
rect 2611 9037 2687 9040
rect 3334 9037 3400 9040
rect 2611 9035 3710 9037
rect 2611 8979 2621 9035
rect 2677 8979 3339 9035
rect 3395 8979 3710 9035
rect 2611 8977 3710 8979
rect 2611 8974 2687 8977
rect 3334 8974 3400 8977
rect -304 7724 -228 7729
rect -304 7669 -294 7724
rect -1528 7608 -294 7669
rect -304 7548 -294 7608
rect -238 7548 -228 7724
rect -304 7543 -228 7548
rect 8387 7469 8453 7472
rect 8044 7467 8453 7469
rect 8044 7411 8392 7467
rect 8448 7411 8453 7467
rect 8044 7409 8453 7411
rect 8387 7406 8453 7409
<< via3 >>
rect -1290 9947 -1226 9952
rect -1290 9891 -1285 9947
rect -1285 9891 -1229 9947
rect -1229 9891 -1226 9947
rect -1290 9886 -1226 9891
<< metal4 >>
rect -1384 9952 -1207 9967
rect -1384 9886 -1290 9952
rect -1226 9886 -1207 9952
rect -1384 9871 -1207 9886
use cap_op  cap_op_0
timestamp 1762701392
transform 1 0 -5288 0 1 10081
box -4498 -3960 3990 3640
use differential_pair  differential_pair_0
timestamp 1720116957
transform 1 0 4032 0 1 8666
box -606 -124 5240 892
use nmos_tail_current  nmos_tail_current_0
timestamp 1720118050
transform -1 0 8043 0 -1 8158
box -321 -141 8599 1579
use pmos_current_bgr_2  pmos_current_bgr_2_0
timestamp 1720112176
transform -1 0 8259 0 1 11400
box -250 -1450 4496 516
use resistor_op_tt  resistor_op_tt_0
timestamp 1720284839
transform 0 -1 5238 -1 0 9265
box -417 2220 767 6092
use secondstage  secondstage_0
timestamp 1762874024
transform 1 0 -801 0 1 10039
box -172 -89 4426 929
<< labels >>
flabel metal1 3667 9996 3667 9996 0 FreeSans 1600 0 0 0 vdde
port 4 nsew
flabel metal2 6567 9067 6567 9067 0 FreeSans 1600 0 0 0 plus
port 3 nsew
flabel metal1 5954 9068 5954 9068 0 FreeSans 1600 0 0 0 minus
port 1 nsew
flabel metal2 4348 8395 4348 8395 0 FreeSans 1600 0 0 0 AVSS
port 0 nsew
flabel metal3 -1313 10453 -1311 10453 0 FreeSans 1600 0 0 0 out
port 2 nsew
<< end >>
