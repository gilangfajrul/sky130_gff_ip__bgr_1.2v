magic
tech sky130A
magscale 1 2
timestamp 1720952586
<< dnwell >>
rect -17914 13826 9178 22978
rect -17914 226 -1066 13826
rect 330 9996 6378 12566
rect 250 1487 7248 8485
rect 8559 226 9178 13826
rect -17914 -412 9178 226
<< nwell >>
rect -17994 22772 9258 23058
rect -17994 -206 -17708 22772
rect -16736 14678 -2960 17678
rect -16736 14626 -3776 14678
rect 250 12360 6458 12646
rect 250 10202 536 12360
rect 6172 11948 6458 12360
rect 4800 10550 6458 11948
rect 6172 10202 6458 10550
rect 250 9916 6458 10202
rect 8972 -206 9258 22772
rect -17994 -492 9258 -206
<< pwell >>
rect -17561 20831 8723 22741
rect -13185 19267 8723 20831
rect -7201 17703 8723 19267
rect -1328 14640 8723 17703
rect 580 10205 4796 12357
rect 303 8279 1643 8432
rect 303 7245 456 8279
rect 1490 7245 1643 8279
rect 303 7092 1643 7245
rect 1691 8279 3031 8432
rect 1691 7245 1844 8279
rect 2878 7245 3031 8279
rect 1691 7092 3031 7245
rect 3079 8279 4419 8432
rect 3079 7245 3232 8279
rect 4266 7245 4419 8279
rect 3079 7092 4419 7245
rect 4467 8279 5807 8432
rect 4467 7245 4620 8279
rect 5654 7245 5807 8279
rect 4467 7092 5807 7245
rect 5855 8279 7195 8432
rect 5855 7245 6008 8279
rect 7042 7245 7195 8279
rect 5855 7092 7195 7245
rect 303 6891 1643 7044
rect 303 5857 456 6891
rect 1490 5857 1643 6891
rect 303 5704 1643 5857
rect 1691 6891 3031 7044
rect 1691 5857 1844 6891
rect 2878 5857 3031 6891
rect 1691 5704 3031 5857
rect 3079 6891 4419 7044
rect 3079 5857 3232 6891
rect 4266 5857 4419 6891
rect 3079 5704 4419 5857
rect 4467 6891 5807 7044
rect 4467 5857 4620 6891
rect 5654 5857 5807 6891
rect 4467 5704 5807 5857
rect 5855 6891 7195 7044
rect 5855 5857 6008 6891
rect 7042 5857 7195 6891
rect 5855 5704 7195 5857
rect 303 5503 1643 5656
rect 303 4469 456 5503
rect 1490 4469 1643 5503
rect 303 4316 1643 4469
rect 1691 5503 3031 5656
rect 1691 4469 1844 5503
rect 2878 4469 3031 5503
rect 1691 4316 3031 4469
rect 3079 5503 4419 5656
rect 3079 4469 3232 5503
rect 4266 4469 4419 5503
rect 3079 4316 4419 4469
rect 4467 5503 5807 5656
rect 4467 4469 4620 5503
rect 5654 4469 5807 5503
rect 4467 4316 5807 4469
rect 5855 5503 7195 5656
rect 5855 4469 6008 5503
rect 7042 4469 7195 5503
rect 5855 4316 7195 4469
rect 303 4115 1643 4268
rect 303 3081 456 4115
rect 1490 3081 1643 4115
rect 303 2928 1643 3081
rect 1691 4115 3031 4268
rect 1691 3081 1844 4115
rect 2878 3081 3031 4115
rect 1691 2928 3031 3081
rect 3079 4115 4419 4268
rect 3079 3081 3232 4115
rect 4266 3081 4419 4115
rect 3079 2928 4419 3081
rect 4467 4115 5807 4268
rect 4467 3081 4620 4115
rect 5654 3081 5807 4115
rect 4467 2928 5807 3081
rect 5855 4115 7195 4268
rect 5855 3081 6008 4115
rect 7042 3081 7195 4115
rect 5855 2928 7195 3081
rect 303 2727 1643 2880
rect 303 1693 456 2727
rect 1490 1693 1643 2727
rect 303 1540 1643 1693
rect 1691 2727 3031 2880
rect 1691 1693 1844 2727
rect 2878 1693 3031 2727
rect 1691 1540 3031 1693
rect 3079 2727 4419 2880
rect 3079 1693 3232 2727
rect 4266 1693 4419 2727
rect 3079 1540 4419 1693
rect 4467 2727 5807 2880
rect 4467 1693 4620 2727
rect 5654 1693 5807 2727
rect 4467 1540 5807 1693
rect 5855 2727 7195 2880
rect 5855 1693 6008 2727
rect 7042 1693 7195 2727
rect 5855 1540 7195 1693
<< nbase >>
rect 456 7245 1490 8279
rect 1844 7245 2878 8279
rect 3232 7245 4266 8279
rect 4620 7245 5654 8279
rect 6008 7245 7042 8279
rect 456 5857 1490 6891
rect 1844 5857 2878 6891
rect 3232 5857 4266 6891
rect 4620 5857 5654 6891
rect 6008 5857 7042 6891
rect 456 4469 1490 5503
rect 1844 4469 2878 5503
rect 3232 4469 4266 5503
rect 4620 4469 5654 5503
rect 6008 4469 7042 5503
rect 456 3081 1490 4115
rect 1844 3081 2878 4115
rect 3232 3081 4266 4115
rect 4620 3081 5654 4115
rect 6008 3081 7042 4115
rect 456 1693 1490 2727
rect 1844 1693 2878 2727
rect 3232 1693 4266 2727
rect 4620 1693 5654 2727
rect 6008 1693 7042 2727
<< nmos >>
rect -1124 17252 -1094 17452
rect -1036 17252 -836 17452
rect -778 17252 -578 17452
rect -520 17252 -490 17452
rect -1124 16942 -1094 17142
rect -1036 16942 -836 17142
rect -778 16942 -578 17142
rect -520 16942 -490 17142
rect -46 17264 -16 17464
rect 154 17264 4154 17464
rect 4324 17264 8324 17464
rect 8494 17264 8524 17464
rect -46 16870 -16 17070
rect 154 16870 4154 17070
rect 4324 16870 8324 17070
rect 8494 16870 8524 17070
rect -46 16476 -16 16676
rect 154 16476 4154 16676
rect 4324 16476 8324 16676
rect 8494 16476 8524 16676
rect -46 16082 -16 16282
rect 154 16082 4154 16282
rect 4324 16082 8324 16282
rect 8494 16082 8524 16282
rect 3059 15366 3089 15546
rect 3147 15366 5747 15546
rect 5805 15366 8405 15546
rect 8463 15366 8493 15546
rect 3059 14934 3089 15114
rect 3147 14934 5747 15114
rect 5805 14934 8405 15114
rect 8463 14934 8493 15114
<< pmos >>
rect -16471 17266 -16441 17466
rect -16383 17266 -14383 17466
rect -14325 17266 -12325 17466
rect -12267 17266 -10267 17466
rect -10209 17266 -8209 17466
rect -8151 17266 -8121 17466
rect -16471 16787 -16441 16987
rect -16383 16787 -14383 16987
rect -14325 16787 -12325 16987
rect -12267 16787 -10267 16987
rect -10209 16787 -8209 16987
rect -8151 16787 -8121 16987
rect -16471 16317 -16441 16517
rect -16383 16317 -14383 16517
rect -14325 16317 -12325 16517
rect -12267 16317 -10267 16517
rect -10209 16317 -8209 16517
rect -8151 16317 -8121 16517
rect -16471 15838 -16441 16038
rect -16383 15838 -14383 16038
rect -14325 15838 -12325 16038
rect -12267 15838 -10267 16038
rect -10209 15838 -8209 16038
rect -8151 15838 -8121 16038
rect -7450 17172 -7420 17372
rect -7362 17172 -5362 17372
rect -5304 17172 -3304 17372
rect -3246 17172 -3216 17372
rect -7450 16740 -7420 16940
rect -7362 16740 -5362 16940
rect -5304 16740 -3304 16940
rect -3246 16740 -3216 16940
rect -7450 16270 -7420 16470
rect -7362 16270 -5362 16470
rect -5304 16270 -3304 16470
rect -3246 16270 -3216 16470
rect -7450 15838 -7420 16038
rect -7362 15838 -5362 16038
rect -5304 15838 -3304 16038
rect -3246 15838 -3216 16038
rect -12322 15224 -12292 15424
rect -12234 15224 -10234 15424
rect -10176 15224 -8176 15424
rect -8118 15224 -8088 15424
rect -12322 14830 -12292 15030
rect -12234 14830 -10234 15030
rect -10176 14830 -8176 15030
rect -8118 14830 -8088 15030
rect -7416 15289 -7386 15489
rect -7328 15289 -5328 15489
rect -5270 15289 -3270 15489
rect -3212 15289 -3182 15489
rect -7416 14813 -7386 15013
rect -7328 14813 -5328 15013
rect -5270 14813 -3270 15013
rect -3212 14813 -3182 15013
rect 4989 11736 5389 11766
rect 5583 11736 5983 11766
rect 4989 11278 5389 11678
rect 5583 11278 5983 11678
rect 4989 10820 5389 11220
rect 5583 10820 5983 11220
rect 4989 10732 5389 10762
rect 5583 10732 5983 10762
<< nmoslvt >>
rect 750 11378 780 12178
rect 838 11378 1038 12178
rect 1096 11378 1296 12178
rect 1354 11378 1384 12178
rect 750 10384 780 11184
rect 838 10384 1038 11184
rect 1096 10384 1296 11184
rect 1354 10384 1384 11184
rect 1642 11378 1672 12178
rect 1730 11378 1930 12178
rect 1988 11378 2188 12178
rect 2246 11378 2276 12178
rect 1642 10384 1672 11184
rect 1730 10384 1930 11184
rect 1988 10384 2188 11184
rect 2246 10384 2276 11184
rect 2534 11378 2564 12178
rect 2622 11378 2822 12178
rect 2880 11378 3080 12178
rect 3138 11378 3168 12178
rect 2534 10384 2564 11184
rect 2622 10384 2822 11184
rect 2880 10384 3080 11184
rect 3138 10384 3168 11184
rect 3426 11378 3456 12178
rect 3514 11378 3714 12178
rect 3772 11378 3972 12178
rect 4030 11378 4060 12178
rect 3426 10384 3456 11184
rect 3514 10384 3714 11184
rect 3772 10384 3972 11184
rect 4030 10384 4060 11184
rect 4416 12125 4616 12155
rect 4416 11867 4616 12067
rect 4416 11609 4616 11809
rect 4416 11521 4616 11551
rect 4416 11011 4616 11041
rect 4416 10753 4616 10953
rect 4416 10495 4616 10695
rect 4416 10407 4616 10437
<< ndiff >>
rect -1182 17440 -1124 17452
rect -1182 17264 -1170 17440
rect -1136 17264 -1124 17440
rect -1182 17252 -1124 17264
rect -1094 17440 -1036 17452
rect -1094 17264 -1082 17440
rect -1048 17264 -1036 17440
rect -1094 17252 -1036 17264
rect -836 17440 -778 17452
rect -836 17264 -824 17440
rect -790 17264 -778 17440
rect -836 17252 -778 17264
rect -578 17440 -520 17452
rect -578 17264 -566 17440
rect -532 17264 -520 17440
rect -578 17252 -520 17264
rect -490 17440 -432 17452
rect -490 17264 -478 17440
rect -444 17264 -432 17440
rect -490 17252 -432 17264
rect -1182 17130 -1124 17142
rect -1182 16954 -1170 17130
rect -1136 16954 -1124 17130
rect -1182 16942 -1124 16954
rect -1094 17130 -1036 17142
rect -1094 16954 -1082 17130
rect -1048 16954 -1036 17130
rect -1094 16942 -1036 16954
rect -836 17130 -778 17142
rect -836 16954 -824 17130
rect -790 16954 -778 17130
rect -836 16942 -778 16954
rect -578 17130 -520 17142
rect -578 16954 -566 17130
rect -532 16954 -520 17130
rect -578 16942 -520 16954
rect -490 17130 -432 17142
rect -490 16954 -478 17130
rect -444 16954 -432 17130
rect -490 16942 -432 16954
rect -104 17452 -46 17464
rect -104 17276 -92 17452
rect -58 17276 -46 17452
rect -104 17264 -46 17276
rect -16 17452 42 17464
rect -16 17276 -4 17452
rect 30 17276 42 17452
rect -16 17264 42 17276
rect 96 17452 154 17464
rect 96 17276 108 17452
rect 142 17276 154 17452
rect 96 17264 154 17276
rect 4154 17452 4212 17464
rect 4154 17276 4166 17452
rect 4200 17276 4212 17452
rect 4154 17264 4212 17276
rect 4266 17452 4324 17464
rect 4266 17276 4278 17452
rect 4312 17276 4324 17452
rect 4266 17264 4324 17276
rect 8324 17452 8382 17464
rect 8324 17276 8336 17452
rect 8370 17276 8382 17452
rect 8324 17264 8382 17276
rect 8436 17452 8494 17464
rect 8436 17276 8448 17452
rect 8482 17276 8494 17452
rect 8436 17264 8494 17276
rect 8524 17452 8582 17464
rect 8524 17276 8536 17452
rect 8570 17276 8582 17452
rect 8524 17264 8582 17276
rect -104 17058 -46 17070
rect -104 16882 -92 17058
rect -58 16882 -46 17058
rect -104 16870 -46 16882
rect -16 17058 42 17070
rect -16 16882 -4 17058
rect 30 16882 42 17058
rect -16 16870 42 16882
rect 96 17058 154 17070
rect 96 16882 108 17058
rect 142 16882 154 17058
rect 96 16870 154 16882
rect 4154 17058 4212 17070
rect 4154 16882 4166 17058
rect 4200 16882 4212 17058
rect 4154 16870 4212 16882
rect 4266 17058 4324 17070
rect 4266 16882 4278 17058
rect 4312 16882 4324 17058
rect 4266 16870 4324 16882
rect 8324 17058 8382 17070
rect 8324 16882 8336 17058
rect 8370 16882 8382 17058
rect 8324 16870 8382 16882
rect 8436 17058 8494 17070
rect 8436 16882 8448 17058
rect 8482 16882 8494 17058
rect 8436 16870 8494 16882
rect 8524 17058 8582 17070
rect 8524 16882 8536 17058
rect 8570 16882 8582 17058
rect 8524 16870 8582 16882
rect -104 16664 -46 16676
rect -104 16488 -92 16664
rect -58 16488 -46 16664
rect -104 16476 -46 16488
rect -16 16664 42 16676
rect -16 16488 -4 16664
rect 30 16488 42 16664
rect -16 16476 42 16488
rect 96 16664 154 16676
rect 96 16488 108 16664
rect 142 16488 154 16664
rect 96 16476 154 16488
rect 4154 16664 4212 16676
rect 4154 16488 4166 16664
rect 4200 16488 4212 16664
rect 4154 16476 4212 16488
rect 4266 16664 4324 16676
rect 4266 16488 4278 16664
rect 4312 16488 4324 16664
rect 4266 16476 4324 16488
rect 8324 16664 8382 16676
rect 8324 16488 8336 16664
rect 8370 16488 8382 16664
rect 8324 16476 8382 16488
rect 8436 16664 8494 16676
rect 8436 16488 8448 16664
rect 8482 16488 8494 16664
rect 8436 16476 8494 16488
rect 8524 16664 8582 16676
rect 8524 16488 8536 16664
rect 8570 16488 8582 16664
rect 8524 16476 8582 16488
rect -104 16270 -46 16282
rect -104 16094 -92 16270
rect -58 16094 -46 16270
rect -104 16082 -46 16094
rect -16 16270 42 16282
rect -16 16094 -4 16270
rect 30 16094 42 16270
rect -16 16082 42 16094
rect 96 16270 154 16282
rect 96 16094 108 16270
rect 142 16094 154 16270
rect 96 16082 154 16094
rect 4154 16270 4212 16282
rect 4154 16094 4166 16270
rect 4200 16094 4212 16270
rect 4154 16082 4212 16094
rect 4266 16270 4324 16282
rect 4266 16094 4278 16270
rect 4312 16094 4324 16270
rect 4266 16082 4324 16094
rect 8324 16270 8382 16282
rect 8324 16094 8336 16270
rect 8370 16094 8382 16270
rect 8324 16082 8382 16094
rect 8436 16270 8494 16282
rect 8436 16094 8448 16270
rect 8482 16094 8494 16270
rect 8436 16082 8494 16094
rect 8524 16270 8582 16282
rect 8524 16094 8536 16270
rect 8570 16094 8582 16270
rect 8524 16082 8582 16094
rect 3001 15534 3059 15546
rect 3001 15378 3013 15534
rect 3047 15378 3059 15534
rect 3001 15366 3059 15378
rect 3089 15534 3147 15546
rect 3089 15378 3101 15534
rect 3135 15378 3147 15534
rect 3089 15366 3147 15378
rect 5747 15534 5805 15546
rect 5747 15378 5759 15534
rect 5793 15378 5805 15534
rect 5747 15366 5805 15378
rect 8405 15534 8463 15546
rect 8405 15378 8417 15534
rect 8451 15378 8463 15534
rect 8405 15366 8463 15378
rect 8493 15534 8551 15546
rect 8493 15378 8505 15534
rect 8539 15378 8551 15534
rect 8493 15366 8551 15378
rect 3001 15102 3059 15114
rect 3001 14946 3013 15102
rect 3047 14946 3059 15102
rect 3001 14934 3059 14946
rect 3089 15102 3147 15114
rect 3089 14946 3101 15102
rect 3135 14946 3147 15102
rect 3089 14934 3147 14946
rect 5747 15102 5805 15114
rect 5747 14946 5759 15102
rect 5793 14946 5805 15102
rect 5747 14934 5805 14946
rect 8405 15102 8463 15114
rect 8405 14946 8417 15102
rect 8451 14946 8463 15102
rect 8405 14934 8463 14946
rect 8493 15102 8551 15114
rect 8493 14946 8505 15102
rect 8539 14946 8551 15102
rect 8493 14934 8551 14946
rect 692 12166 750 12178
rect 692 11390 704 12166
rect 738 11390 750 12166
rect 692 11378 750 11390
rect 780 12166 838 12178
rect 780 11390 792 12166
rect 826 11390 838 12166
rect 780 11378 838 11390
rect 1038 12166 1096 12178
rect 1038 11390 1050 12166
rect 1084 11390 1096 12166
rect 1038 11378 1096 11390
rect 1296 12166 1354 12178
rect 1296 11390 1308 12166
rect 1342 11390 1354 12166
rect 1296 11378 1354 11390
rect 1384 12166 1442 12178
rect 1384 11390 1396 12166
rect 1430 11390 1442 12166
rect 1384 11378 1442 11390
rect 692 11172 750 11184
rect 692 10396 704 11172
rect 738 10396 750 11172
rect 692 10384 750 10396
rect 780 11172 838 11184
rect 780 10396 792 11172
rect 826 10396 838 11172
rect 780 10384 838 10396
rect 1038 11172 1096 11184
rect 1038 10396 1050 11172
rect 1084 10396 1096 11172
rect 1038 10384 1096 10396
rect 1296 11172 1354 11184
rect 1296 10396 1308 11172
rect 1342 10396 1354 11172
rect 1296 10384 1354 10396
rect 1384 11172 1442 11184
rect 1384 10396 1396 11172
rect 1430 10396 1442 11172
rect 1384 10384 1442 10396
rect 1584 12166 1642 12178
rect 1584 11390 1596 12166
rect 1630 11390 1642 12166
rect 1584 11378 1642 11390
rect 1672 12166 1730 12178
rect 1672 11390 1684 12166
rect 1718 11390 1730 12166
rect 1672 11378 1730 11390
rect 1930 12166 1988 12178
rect 1930 11390 1942 12166
rect 1976 11390 1988 12166
rect 1930 11378 1988 11390
rect 2188 12166 2246 12178
rect 2188 11390 2200 12166
rect 2234 11390 2246 12166
rect 2188 11378 2246 11390
rect 2276 12166 2334 12178
rect 2276 11390 2288 12166
rect 2322 11390 2334 12166
rect 2276 11378 2334 11390
rect 1584 11172 1642 11184
rect 1584 10396 1596 11172
rect 1630 10396 1642 11172
rect 1584 10384 1642 10396
rect 1672 11172 1730 11184
rect 1672 10396 1684 11172
rect 1718 10396 1730 11172
rect 1672 10384 1730 10396
rect 1930 11172 1988 11184
rect 1930 10396 1942 11172
rect 1976 10396 1988 11172
rect 1930 10384 1988 10396
rect 2188 11172 2246 11184
rect 2188 10396 2200 11172
rect 2234 10396 2246 11172
rect 2188 10384 2246 10396
rect 2276 11172 2334 11184
rect 2276 10396 2288 11172
rect 2322 10396 2334 11172
rect 2276 10384 2334 10396
rect 2476 12166 2534 12178
rect 2476 11390 2488 12166
rect 2522 11390 2534 12166
rect 2476 11378 2534 11390
rect 2564 12166 2622 12178
rect 2564 11390 2576 12166
rect 2610 11390 2622 12166
rect 2564 11378 2622 11390
rect 2822 12166 2880 12178
rect 2822 11390 2834 12166
rect 2868 11390 2880 12166
rect 2822 11378 2880 11390
rect 3080 12166 3138 12178
rect 3080 11390 3092 12166
rect 3126 11390 3138 12166
rect 3080 11378 3138 11390
rect 3168 12166 3226 12178
rect 3168 11390 3180 12166
rect 3214 11390 3226 12166
rect 3168 11378 3226 11390
rect 2476 11172 2534 11184
rect 2476 10396 2488 11172
rect 2522 10396 2534 11172
rect 2476 10384 2534 10396
rect 2564 11172 2622 11184
rect 2564 10396 2576 11172
rect 2610 10396 2622 11172
rect 2564 10384 2622 10396
rect 2822 11172 2880 11184
rect 2822 10396 2834 11172
rect 2868 10396 2880 11172
rect 2822 10384 2880 10396
rect 3080 11172 3138 11184
rect 3080 10396 3092 11172
rect 3126 10396 3138 11172
rect 3080 10384 3138 10396
rect 3168 11172 3226 11184
rect 3168 10396 3180 11172
rect 3214 10396 3226 11172
rect 3168 10384 3226 10396
rect 3368 12166 3426 12178
rect 3368 11390 3380 12166
rect 3414 11390 3426 12166
rect 3368 11378 3426 11390
rect 3456 12166 3514 12178
rect 3456 11390 3468 12166
rect 3502 11390 3514 12166
rect 3456 11378 3514 11390
rect 3714 12166 3772 12178
rect 3714 11390 3726 12166
rect 3760 11390 3772 12166
rect 3714 11378 3772 11390
rect 3972 12166 4030 12178
rect 3972 11390 3984 12166
rect 4018 11390 4030 12166
rect 3972 11378 4030 11390
rect 4060 12166 4118 12178
rect 4060 11390 4072 12166
rect 4106 11390 4118 12166
rect 4060 11378 4118 11390
rect 3368 11172 3426 11184
rect 3368 10396 3380 11172
rect 3414 10396 3426 11172
rect 3368 10384 3426 10396
rect 3456 11172 3514 11184
rect 3456 10396 3468 11172
rect 3502 10396 3514 11172
rect 3456 10384 3514 10396
rect 3714 11172 3772 11184
rect 3714 10396 3726 11172
rect 3760 10396 3772 11172
rect 3714 10384 3772 10396
rect 3972 11172 4030 11184
rect 3972 10396 3984 11172
rect 4018 10396 4030 11172
rect 3972 10384 4030 10396
rect 4060 11172 4118 11184
rect 4060 10396 4072 11172
rect 4106 10396 4118 11172
rect 4060 10384 4118 10396
rect 4416 12201 4616 12213
rect 4416 12167 4428 12201
rect 4604 12167 4616 12201
rect 4416 12155 4616 12167
rect 4416 12113 4616 12125
rect 4416 12079 4428 12113
rect 4604 12079 4616 12113
rect 4416 12067 4616 12079
rect 4416 11855 4616 11867
rect 4416 11821 4428 11855
rect 4604 11821 4616 11855
rect 4416 11809 4616 11821
rect 4416 11597 4616 11609
rect 4416 11563 4428 11597
rect 4604 11563 4616 11597
rect 4416 11551 4616 11563
rect 4416 11509 4616 11521
rect 4416 11475 4428 11509
rect 4604 11475 4616 11509
rect 4416 11463 4616 11475
rect 4416 11087 4616 11099
rect 4416 11053 4428 11087
rect 4604 11053 4616 11087
rect 4416 11041 4616 11053
rect 4416 10999 4616 11011
rect 4416 10965 4428 10999
rect 4604 10965 4616 10999
rect 4416 10953 4616 10965
rect 4416 10741 4616 10753
rect 4416 10707 4428 10741
rect 4604 10707 4616 10741
rect 4416 10695 4616 10707
rect 4416 10483 4616 10495
rect 4416 10449 4428 10483
rect 4604 10449 4616 10483
rect 4416 10437 4616 10449
rect 4416 10395 4616 10407
rect 4416 10361 4428 10395
rect 4604 10361 4616 10395
rect 4416 10349 4616 10361
<< pdiff >>
rect -16529 17454 -16471 17466
rect -16529 17278 -16517 17454
rect -16483 17278 -16471 17454
rect -16529 17266 -16471 17278
rect -16441 17454 -16383 17466
rect -16441 17278 -16429 17454
rect -16395 17278 -16383 17454
rect -16441 17266 -16383 17278
rect -14383 17454 -14325 17466
rect -14383 17278 -14371 17454
rect -14337 17278 -14325 17454
rect -14383 17266 -14325 17278
rect -12325 17454 -12267 17466
rect -12325 17278 -12313 17454
rect -12279 17278 -12267 17454
rect -12325 17266 -12267 17278
rect -10267 17454 -10209 17466
rect -10267 17278 -10255 17454
rect -10221 17278 -10209 17454
rect -10267 17266 -10209 17278
rect -8209 17454 -8151 17466
rect -8209 17278 -8197 17454
rect -8163 17278 -8151 17454
rect -8209 17266 -8151 17278
rect -8121 17454 -8063 17466
rect -8121 17278 -8109 17454
rect -8075 17278 -8063 17454
rect -8121 17266 -8063 17278
rect -16529 16975 -16471 16987
rect -16529 16799 -16517 16975
rect -16483 16799 -16471 16975
rect -16529 16787 -16471 16799
rect -16441 16975 -16383 16987
rect -16441 16799 -16429 16975
rect -16395 16799 -16383 16975
rect -16441 16787 -16383 16799
rect -14383 16975 -14325 16987
rect -14383 16799 -14371 16975
rect -14337 16799 -14325 16975
rect -14383 16787 -14325 16799
rect -12325 16975 -12267 16987
rect -12325 16799 -12313 16975
rect -12279 16799 -12267 16975
rect -12325 16787 -12267 16799
rect -10267 16975 -10209 16987
rect -10267 16799 -10255 16975
rect -10221 16799 -10209 16975
rect -10267 16787 -10209 16799
rect -8209 16975 -8151 16987
rect -8209 16799 -8197 16975
rect -8163 16799 -8151 16975
rect -8209 16787 -8151 16799
rect -8121 16975 -8063 16987
rect -8121 16799 -8109 16975
rect -8075 16799 -8063 16975
rect -8121 16787 -8063 16799
rect -16529 16505 -16471 16517
rect -16529 16329 -16517 16505
rect -16483 16329 -16471 16505
rect -16529 16317 -16471 16329
rect -16441 16505 -16383 16517
rect -16441 16329 -16429 16505
rect -16395 16329 -16383 16505
rect -16441 16317 -16383 16329
rect -14383 16505 -14325 16517
rect -14383 16329 -14371 16505
rect -14337 16329 -14325 16505
rect -14383 16317 -14325 16329
rect -12325 16505 -12267 16517
rect -12325 16329 -12313 16505
rect -12279 16329 -12267 16505
rect -12325 16317 -12267 16329
rect -10267 16505 -10209 16517
rect -10267 16329 -10255 16505
rect -10221 16329 -10209 16505
rect -10267 16317 -10209 16329
rect -8209 16505 -8151 16517
rect -8209 16329 -8197 16505
rect -8163 16329 -8151 16505
rect -8209 16317 -8151 16329
rect -8121 16505 -8063 16517
rect -8121 16329 -8109 16505
rect -8075 16329 -8063 16505
rect -8121 16317 -8063 16329
rect -16529 16026 -16471 16038
rect -16529 15850 -16517 16026
rect -16483 15850 -16471 16026
rect -16529 15838 -16471 15850
rect -16441 16026 -16383 16038
rect -16441 15850 -16429 16026
rect -16395 15850 -16383 16026
rect -16441 15838 -16383 15850
rect -14383 16026 -14325 16038
rect -14383 15850 -14371 16026
rect -14337 15850 -14325 16026
rect -14383 15838 -14325 15850
rect -12325 16026 -12267 16038
rect -12325 15850 -12313 16026
rect -12279 15850 -12267 16026
rect -12325 15838 -12267 15850
rect -10267 16026 -10209 16038
rect -10267 15850 -10255 16026
rect -10221 15850 -10209 16026
rect -10267 15838 -10209 15850
rect -8209 16026 -8151 16038
rect -8209 15850 -8197 16026
rect -8163 15850 -8151 16026
rect -8209 15838 -8151 15850
rect -8121 16026 -8063 16038
rect -8121 15850 -8109 16026
rect -8075 15850 -8063 16026
rect -8121 15838 -8063 15850
rect -7508 17360 -7450 17372
rect -7508 17184 -7496 17360
rect -7462 17184 -7450 17360
rect -7508 17172 -7450 17184
rect -7420 17360 -7362 17372
rect -7420 17184 -7408 17360
rect -7374 17184 -7362 17360
rect -7420 17172 -7362 17184
rect -5362 17360 -5304 17372
rect -5362 17184 -5350 17360
rect -5316 17184 -5304 17360
rect -5362 17172 -5304 17184
rect -3304 17360 -3246 17372
rect -3304 17184 -3292 17360
rect -3258 17184 -3246 17360
rect -3304 17172 -3246 17184
rect -3216 17360 -3158 17372
rect -3216 17184 -3204 17360
rect -3170 17184 -3158 17360
rect -3216 17172 -3158 17184
rect -7508 16928 -7450 16940
rect -7508 16752 -7496 16928
rect -7462 16752 -7450 16928
rect -7508 16740 -7450 16752
rect -7420 16928 -7362 16940
rect -7420 16752 -7408 16928
rect -7374 16752 -7362 16928
rect -7420 16740 -7362 16752
rect -5362 16928 -5304 16940
rect -5362 16752 -5350 16928
rect -5316 16752 -5304 16928
rect -5362 16740 -5304 16752
rect -3304 16928 -3246 16940
rect -3304 16752 -3292 16928
rect -3258 16752 -3246 16928
rect -3304 16740 -3246 16752
rect -3216 16928 -3158 16940
rect -3216 16752 -3204 16928
rect -3170 16752 -3158 16928
rect -3216 16740 -3158 16752
rect -7508 16458 -7450 16470
rect -7508 16282 -7496 16458
rect -7462 16282 -7450 16458
rect -7508 16270 -7450 16282
rect -7420 16458 -7362 16470
rect -7420 16282 -7408 16458
rect -7374 16282 -7362 16458
rect -7420 16270 -7362 16282
rect -5362 16458 -5304 16470
rect -5362 16282 -5350 16458
rect -5316 16282 -5304 16458
rect -5362 16270 -5304 16282
rect -3304 16458 -3246 16470
rect -3304 16282 -3292 16458
rect -3258 16282 -3246 16458
rect -3304 16270 -3246 16282
rect -3216 16458 -3158 16470
rect -3216 16282 -3204 16458
rect -3170 16282 -3158 16458
rect -3216 16270 -3158 16282
rect -7508 16026 -7450 16038
rect -7508 15850 -7496 16026
rect -7462 15850 -7450 16026
rect -7508 15838 -7450 15850
rect -7420 16026 -7362 16038
rect -7420 15850 -7408 16026
rect -7374 15850 -7362 16026
rect -7420 15838 -7362 15850
rect -5362 16026 -5304 16038
rect -5362 15850 -5350 16026
rect -5316 15850 -5304 16026
rect -5362 15838 -5304 15850
rect -3304 16026 -3246 16038
rect -3304 15850 -3292 16026
rect -3258 15850 -3246 16026
rect -3304 15838 -3246 15850
rect -3216 16026 -3158 16038
rect -3216 15850 -3204 16026
rect -3170 15850 -3158 16026
rect -3216 15838 -3158 15850
rect -12380 15412 -12322 15424
rect -12380 15236 -12368 15412
rect -12334 15236 -12322 15412
rect -12380 15224 -12322 15236
rect -12292 15412 -12234 15424
rect -12292 15236 -12280 15412
rect -12246 15236 -12234 15412
rect -12292 15224 -12234 15236
rect -10234 15412 -10176 15424
rect -10234 15236 -10222 15412
rect -10188 15236 -10176 15412
rect -10234 15224 -10176 15236
rect -8176 15412 -8118 15424
rect -8176 15236 -8164 15412
rect -8130 15236 -8118 15412
rect -8176 15224 -8118 15236
rect -8088 15412 -8030 15424
rect -8088 15236 -8076 15412
rect -8042 15236 -8030 15412
rect -8088 15224 -8030 15236
rect -12380 15018 -12322 15030
rect -12380 14842 -12368 15018
rect -12334 14842 -12322 15018
rect -12380 14830 -12322 14842
rect -12292 15018 -12234 15030
rect -12292 14842 -12280 15018
rect -12246 14842 -12234 15018
rect -12292 14830 -12234 14842
rect -10234 15018 -10176 15030
rect -10234 14842 -10222 15018
rect -10188 14842 -10176 15018
rect -10234 14830 -10176 14842
rect -8176 15018 -8118 15030
rect -8176 14842 -8164 15018
rect -8130 14842 -8118 15018
rect -8176 14830 -8118 14842
rect -8088 15018 -8030 15030
rect -8088 14842 -8076 15018
rect -8042 14842 -8030 15018
rect -8088 14830 -8030 14842
rect -7474 15477 -7416 15489
rect -7474 15301 -7462 15477
rect -7428 15301 -7416 15477
rect -7474 15289 -7416 15301
rect -7386 15477 -7328 15489
rect -7386 15301 -7374 15477
rect -7340 15301 -7328 15477
rect -7386 15289 -7328 15301
rect -5328 15477 -5270 15489
rect -5328 15301 -5316 15477
rect -5282 15301 -5270 15477
rect -5328 15289 -5270 15301
rect -3270 15477 -3212 15489
rect -3270 15301 -3258 15477
rect -3224 15301 -3212 15477
rect -3270 15289 -3212 15301
rect -3182 15477 -3124 15489
rect -3182 15301 -3170 15477
rect -3136 15301 -3124 15477
rect -3182 15289 -3124 15301
rect -7474 15001 -7416 15013
rect -7474 14825 -7462 15001
rect -7428 14825 -7416 15001
rect -7474 14813 -7416 14825
rect -7386 15001 -7328 15013
rect -7386 14825 -7374 15001
rect -7340 14825 -7328 15001
rect -7386 14813 -7328 14825
rect -5328 15001 -5270 15013
rect -5328 14825 -5316 15001
rect -5282 14825 -5270 15001
rect -5328 14813 -5270 14825
rect -3270 15001 -3212 15013
rect -3270 14825 -3258 15001
rect -3224 14825 -3212 15001
rect -3270 14813 -3212 14825
rect -3182 15001 -3124 15013
rect -3182 14825 -3170 15001
rect -3136 14825 -3124 15001
rect -3182 14813 -3124 14825
rect 4989 11812 5389 11824
rect 4989 11778 5001 11812
rect 5377 11778 5389 11812
rect 4989 11766 5389 11778
rect 5583 11812 5983 11824
rect 5583 11778 5595 11812
rect 5971 11778 5983 11812
rect 5583 11766 5983 11778
rect 4989 11724 5389 11736
rect 4989 11690 5001 11724
rect 5377 11690 5389 11724
rect 4989 11678 5389 11690
rect 5583 11724 5983 11736
rect 5583 11690 5595 11724
rect 5971 11690 5983 11724
rect 5583 11678 5983 11690
rect 4989 11266 5389 11278
rect 4989 11232 5001 11266
rect 5377 11232 5389 11266
rect 4989 11220 5389 11232
rect 5583 11266 5983 11278
rect 5583 11232 5595 11266
rect 5971 11232 5983 11266
rect 5583 11220 5983 11232
rect 4989 10808 5389 10820
rect 4989 10774 5001 10808
rect 5377 10774 5389 10808
rect 4989 10762 5389 10774
rect 5583 10808 5983 10820
rect 5583 10774 5595 10808
rect 5971 10774 5983 10808
rect 5583 10762 5983 10774
rect 4989 10720 5389 10732
rect 4989 10686 5001 10720
rect 5377 10686 5389 10720
rect 4989 10674 5389 10686
rect 5583 10720 5983 10732
rect 5583 10686 5595 10720
rect 5971 10686 5983 10720
rect 5583 10674 5983 10686
rect 633 8050 1313 8102
rect 633 8016 685 8050
rect 719 8016 775 8050
rect 809 8016 865 8050
rect 899 8016 955 8050
rect 989 8016 1045 8050
rect 1079 8016 1135 8050
rect 1169 8016 1225 8050
rect 1259 8016 1313 8050
rect 633 7960 1313 8016
rect 633 7926 685 7960
rect 719 7926 775 7960
rect 809 7926 865 7960
rect 899 7926 955 7960
rect 989 7926 1045 7960
rect 1079 7926 1135 7960
rect 1169 7926 1225 7960
rect 1259 7926 1313 7960
rect 633 7870 1313 7926
rect 633 7836 685 7870
rect 719 7836 775 7870
rect 809 7836 865 7870
rect 899 7836 955 7870
rect 989 7836 1045 7870
rect 1079 7836 1135 7870
rect 1169 7836 1225 7870
rect 1259 7836 1313 7870
rect 633 7780 1313 7836
rect 633 7746 685 7780
rect 719 7746 775 7780
rect 809 7746 865 7780
rect 899 7746 955 7780
rect 989 7746 1045 7780
rect 1079 7746 1135 7780
rect 1169 7746 1225 7780
rect 1259 7746 1313 7780
rect 633 7690 1313 7746
rect 633 7656 685 7690
rect 719 7656 775 7690
rect 809 7656 865 7690
rect 899 7656 955 7690
rect 989 7656 1045 7690
rect 1079 7656 1135 7690
rect 1169 7656 1225 7690
rect 1259 7656 1313 7690
rect 633 7600 1313 7656
rect 633 7566 685 7600
rect 719 7566 775 7600
rect 809 7566 865 7600
rect 899 7566 955 7600
rect 989 7566 1045 7600
rect 1079 7566 1135 7600
rect 1169 7566 1225 7600
rect 1259 7566 1313 7600
rect 633 7510 1313 7566
rect 633 7476 685 7510
rect 719 7476 775 7510
rect 809 7476 865 7510
rect 899 7476 955 7510
rect 989 7476 1045 7510
rect 1079 7476 1135 7510
rect 1169 7476 1225 7510
rect 1259 7476 1313 7510
rect 633 7422 1313 7476
rect 2021 8050 2701 8102
rect 2021 8016 2073 8050
rect 2107 8016 2163 8050
rect 2197 8016 2253 8050
rect 2287 8016 2343 8050
rect 2377 8016 2433 8050
rect 2467 8016 2523 8050
rect 2557 8016 2613 8050
rect 2647 8016 2701 8050
rect 2021 7960 2701 8016
rect 2021 7926 2073 7960
rect 2107 7926 2163 7960
rect 2197 7926 2253 7960
rect 2287 7926 2343 7960
rect 2377 7926 2433 7960
rect 2467 7926 2523 7960
rect 2557 7926 2613 7960
rect 2647 7926 2701 7960
rect 2021 7870 2701 7926
rect 2021 7836 2073 7870
rect 2107 7836 2163 7870
rect 2197 7836 2253 7870
rect 2287 7836 2343 7870
rect 2377 7836 2433 7870
rect 2467 7836 2523 7870
rect 2557 7836 2613 7870
rect 2647 7836 2701 7870
rect 2021 7780 2701 7836
rect 2021 7746 2073 7780
rect 2107 7746 2163 7780
rect 2197 7746 2253 7780
rect 2287 7746 2343 7780
rect 2377 7746 2433 7780
rect 2467 7746 2523 7780
rect 2557 7746 2613 7780
rect 2647 7746 2701 7780
rect 2021 7690 2701 7746
rect 2021 7656 2073 7690
rect 2107 7656 2163 7690
rect 2197 7656 2253 7690
rect 2287 7656 2343 7690
rect 2377 7656 2433 7690
rect 2467 7656 2523 7690
rect 2557 7656 2613 7690
rect 2647 7656 2701 7690
rect 2021 7600 2701 7656
rect 2021 7566 2073 7600
rect 2107 7566 2163 7600
rect 2197 7566 2253 7600
rect 2287 7566 2343 7600
rect 2377 7566 2433 7600
rect 2467 7566 2523 7600
rect 2557 7566 2613 7600
rect 2647 7566 2701 7600
rect 2021 7510 2701 7566
rect 2021 7476 2073 7510
rect 2107 7476 2163 7510
rect 2197 7476 2253 7510
rect 2287 7476 2343 7510
rect 2377 7476 2433 7510
rect 2467 7476 2523 7510
rect 2557 7476 2613 7510
rect 2647 7476 2701 7510
rect 2021 7422 2701 7476
rect 3409 8050 4089 8102
rect 3409 8016 3461 8050
rect 3495 8016 3551 8050
rect 3585 8016 3641 8050
rect 3675 8016 3731 8050
rect 3765 8016 3821 8050
rect 3855 8016 3911 8050
rect 3945 8016 4001 8050
rect 4035 8016 4089 8050
rect 3409 7960 4089 8016
rect 3409 7926 3461 7960
rect 3495 7926 3551 7960
rect 3585 7926 3641 7960
rect 3675 7926 3731 7960
rect 3765 7926 3821 7960
rect 3855 7926 3911 7960
rect 3945 7926 4001 7960
rect 4035 7926 4089 7960
rect 3409 7870 4089 7926
rect 3409 7836 3461 7870
rect 3495 7836 3551 7870
rect 3585 7836 3641 7870
rect 3675 7836 3731 7870
rect 3765 7836 3821 7870
rect 3855 7836 3911 7870
rect 3945 7836 4001 7870
rect 4035 7836 4089 7870
rect 3409 7780 4089 7836
rect 3409 7746 3461 7780
rect 3495 7746 3551 7780
rect 3585 7746 3641 7780
rect 3675 7746 3731 7780
rect 3765 7746 3821 7780
rect 3855 7746 3911 7780
rect 3945 7746 4001 7780
rect 4035 7746 4089 7780
rect 3409 7690 4089 7746
rect 3409 7656 3461 7690
rect 3495 7656 3551 7690
rect 3585 7656 3641 7690
rect 3675 7656 3731 7690
rect 3765 7656 3821 7690
rect 3855 7656 3911 7690
rect 3945 7656 4001 7690
rect 4035 7656 4089 7690
rect 3409 7600 4089 7656
rect 3409 7566 3461 7600
rect 3495 7566 3551 7600
rect 3585 7566 3641 7600
rect 3675 7566 3731 7600
rect 3765 7566 3821 7600
rect 3855 7566 3911 7600
rect 3945 7566 4001 7600
rect 4035 7566 4089 7600
rect 3409 7510 4089 7566
rect 3409 7476 3461 7510
rect 3495 7476 3551 7510
rect 3585 7476 3641 7510
rect 3675 7476 3731 7510
rect 3765 7476 3821 7510
rect 3855 7476 3911 7510
rect 3945 7476 4001 7510
rect 4035 7476 4089 7510
rect 3409 7422 4089 7476
rect 4797 8050 5477 8102
rect 4797 8016 4849 8050
rect 4883 8016 4939 8050
rect 4973 8016 5029 8050
rect 5063 8016 5119 8050
rect 5153 8016 5209 8050
rect 5243 8016 5299 8050
rect 5333 8016 5389 8050
rect 5423 8016 5477 8050
rect 4797 7960 5477 8016
rect 4797 7926 4849 7960
rect 4883 7926 4939 7960
rect 4973 7926 5029 7960
rect 5063 7926 5119 7960
rect 5153 7926 5209 7960
rect 5243 7926 5299 7960
rect 5333 7926 5389 7960
rect 5423 7926 5477 7960
rect 4797 7870 5477 7926
rect 4797 7836 4849 7870
rect 4883 7836 4939 7870
rect 4973 7836 5029 7870
rect 5063 7836 5119 7870
rect 5153 7836 5209 7870
rect 5243 7836 5299 7870
rect 5333 7836 5389 7870
rect 5423 7836 5477 7870
rect 4797 7780 5477 7836
rect 4797 7746 4849 7780
rect 4883 7746 4939 7780
rect 4973 7746 5029 7780
rect 5063 7746 5119 7780
rect 5153 7746 5209 7780
rect 5243 7746 5299 7780
rect 5333 7746 5389 7780
rect 5423 7746 5477 7780
rect 4797 7690 5477 7746
rect 4797 7656 4849 7690
rect 4883 7656 4939 7690
rect 4973 7656 5029 7690
rect 5063 7656 5119 7690
rect 5153 7656 5209 7690
rect 5243 7656 5299 7690
rect 5333 7656 5389 7690
rect 5423 7656 5477 7690
rect 4797 7600 5477 7656
rect 4797 7566 4849 7600
rect 4883 7566 4939 7600
rect 4973 7566 5029 7600
rect 5063 7566 5119 7600
rect 5153 7566 5209 7600
rect 5243 7566 5299 7600
rect 5333 7566 5389 7600
rect 5423 7566 5477 7600
rect 4797 7510 5477 7566
rect 4797 7476 4849 7510
rect 4883 7476 4939 7510
rect 4973 7476 5029 7510
rect 5063 7476 5119 7510
rect 5153 7476 5209 7510
rect 5243 7476 5299 7510
rect 5333 7476 5389 7510
rect 5423 7476 5477 7510
rect 4797 7422 5477 7476
rect 6185 8050 6865 8102
rect 6185 8016 6237 8050
rect 6271 8016 6327 8050
rect 6361 8016 6417 8050
rect 6451 8016 6507 8050
rect 6541 8016 6597 8050
rect 6631 8016 6687 8050
rect 6721 8016 6777 8050
rect 6811 8016 6865 8050
rect 6185 7960 6865 8016
rect 6185 7926 6237 7960
rect 6271 7926 6327 7960
rect 6361 7926 6417 7960
rect 6451 7926 6507 7960
rect 6541 7926 6597 7960
rect 6631 7926 6687 7960
rect 6721 7926 6777 7960
rect 6811 7926 6865 7960
rect 6185 7870 6865 7926
rect 6185 7836 6237 7870
rect 6271 7836 6327 7870
rect 6361 7836 6417 7870
rect 6451 7836 6507 7870
rect 6541 7836 6597 7870
rect 6631 7836 6687 7870
rect 6721 7836 6777 7870
rect 6811 7836 6865 7870
rect 6185 7780 6865 7836
rect 6185 7746 6237 7780
rect 6271 7746 6327 7780
rect 6361 7746 6417 7780
rect 6451 7746 6507 7780
rect 6541 7746 6597 7780
rect 6631 7746 6687 7780
rect 6721 7746 6777 7780
rect 6811 7746 6865 7780
rect 6185 7690 6865 7746
rect 6185 7656 6237 7690
rect 6271 7656 6327 7690
rect 6361 7656 6417 7690
rect 6451 7656 6507 7690
rect 6541 7656 6597 7690
rect 6631 7656 6687 7690
rect 6721 7656 6777 7690
rect 6811 7656 6865 7690
rect 6185 7600 6865 7656
rect 6185 7566 6237 7600
rect 6271 7566 6327 7600
rect 6361 7566 6417 7600
rect 6451 7566 6507 7600
rect 6541 7566 6597 7600
rect 6631 7566 6687 7600
rect 6721 7566 6777 7600
rect 6811 7566 6865 7600
rect 6185 7510 6865 7566
rect 6185 7476 6237 7510
rect 6271 7476 6327 7510
rect 6361 7476 6417 7510
rect 6451 7476 6507 7510
rect 6541 7476 6597 7510
rect 6631 7476 6687 7510
rect 6721 7476 6777 7510
rect 6811 7476 6865 7510
rect 6185 7422 6865 7476
rect 633 6662 1313 6714
rect 633 6628 685 6662
rect 719 6628 775 6662
rect 809 6628 865 6662
rect 899 6628 955 6662
rect 989 6628 1045 6662
rect 1079 6628 1135 6662
rect 1169 6628 1225 6662
rect 1259 6628 1313 6662
rect 633 6572 1313 6628
rect 633 6538 685 6572
rect 719 6538 775 6572
rect 809 6538 865 6572
rect 899 6538 955 6572
rect 989 6538 1045 6572
rect 1079 6538 1135 6572
rect 1169 6538 1225 6572
rect 1259 6538 1313 6572
rect 633 6482 1313 6538
rect 633 6448 685 6482
rect 719 6448 775 6482
rect 809 6448 865 6482
rect 899 6448 955 6482
rect 989 6448 1045 6482
rect 1079 6448 1135 6482
rect 1169 6448 1225 6482
rect 1259 6448 1313 6482
rect 633 6392 1313 6448
rect 633 6358 685 6392
rect 719 6358 775 6392
rect 809 6358 865 6392
rect 899 6358 955 6392
rect 989 6358 1045 6392
rect 1079 6358 1135 6392
rect 1169 6358 1225 6392
rect 1259 6358 1313 6392
rect 633 6302 1313 6358
rect 633 6268 685 6302
rect 719 6268 775 6302
rect 809 6268 865 6302
rect 899 6268 955 6302
rect 989 6268 1045 6302
rect 1079 6268 1135 6302
rect 1169 6268 1225 6302
rect 1259 6268 1313 6302
rect 633 6212 1313 6268
rect 633 6178 685 6212
rect 719 6178 775 6212
rect 809 6178 865 6212
rect 899 6178 955 6212
rect 989 6178 1045 6212
rect 1079 6178 1135 6212
rect 1169 6178 1225 6212
rect 1259 6178 1313 6212
rect 633 6122 1313 6178
rect 633 6088 685 6122
rect 719 6088 775 6122
rect 809 6088 865 6122
rect 899 6088 955 6122
rect 989 6088 1045 6122
rect 1079 6088 1135 6122
rect 1169 6088 1225 6122
rect 1259 6088 1313 6122
rect 633 6034 1313 6088
rect 2021 6662 2701 6714
rect 2021 6628 2073 6662
rect 2107 6628 2163 6662
rect 2197 6628 2253 6662
rect 2287 6628 2343 6662
rect 2377 6628 2433 6662
rect 2467 6628 2523 6662
rect 2557 6628 2613 6662
rect 2647 6628 2701 6662
rect 2021 6572 2701 6628
rect 2021 6538 2073 6572
rect 2107 6538 2163 6572
rect 2197 6538 2253 6572
rect 2287 6538 2343 6572
rect 2377 6538 2433 6572
rect 2467 6538 2523 6572
rect 2557 6538 2613 6572
rect 2647 6538 2701 6572
rect 2021 6482 2701 6538
rect 2021 6448 2073 6482
rect 2107 6448 2163 6482
rect 2197 6448 2253 6482
rect 2287 6448 2343 6482
rect 2377 6448 2433 6482
rect 2467 6448 2523 6482
rect 2557 6448 2613 6482
rect 2647 6448 2701 6482
rect 2021 6392 2701 6448
rect 2021 6358 2073 6392
rect 2107 6358 2163 6392
rect 2197 6358 2253 6392
rect 2287 6358 2343 6392
rect 2377 6358 2433 6392
rect 2467 6358 2523 6392
rect 2557 6358 2613 6392
rect 2647 6358 2701 6392
rect 2021 6302 2701 6358
rect 2021 6268 2073 6302
rect 2107 6268 2163 6302
rect 2197 6268 2253 6302
rect 2287 6268 2343 6302
rect 2377 6268 2433 6302
rect 2467 6268 2523 6302
rect 2557 6268 2613 6302
rect 2647 6268 2701 6302
rect 2021 6212 2701 6268
rect 2021 6178 2073 6212
rect 2107 6178 2163 6212
rect 2197 6178 2253 6212
rect 2287 6178 2343 6212
rect 2377 6178 2433 6212
rect 2467 6178 2523 6212
rect 2557 6178 2613 6212
rect 2647 6178 2701 6212
rect 2021 6122 2701 6178
rect 2021 6088 2073 6122
rect 2107 6088 2163 6122
rect 2197 6088 2253 6122
rect 2287 6088 2343 6122
rect 2377 6088 2433 6122
rect 2467 6088 2523 6122
rect 2557 6088 2613 6122
rect 2647 6088 2701 6122
rect 2021 6034 2701 6088
rect 3409 6662 4089 6714
rect 3409 6628 3461 6662
rect 3495 6628 3551 6662
rect 3585 6628 3641 6662
rect 3675 6628 3731 6662
rect 3765 6628 3821 6662
rect 3855 6628 3911 6662
rect 3945 6628 4001 6662
rect 4035 6628 4089 6662
rect 3409 6572 4089 6628
rect 3409 6538 3461 6572
rect 3495 6538 3551 6572
rect 3585 6538 3641 6572
rect 3675 6538 3731 6572
rect 3765 6538 3821 6572
rect 3855 6538 3911 6572
rect 3945 6538 4001 6572
rect 4035 6538 4089 6572
rect 3409 6482 4089 6538
rect 3409 6448 3461 6482
rect 3495 6448 3551 6482
rect 3585 6448 3641 6482
rect 3675 6448 3731 6482
rect 3765 6448 3821 6482
rect 3855 6448 3911 6482
rect 3945 6448 4001 6482
rect 4035 6448 4089 6482
rect 3409 6392 4089 6448
rect 3409 6358 3461 6392
rect 3495 6358 3551 6392
rect 3585 6358 3641 6392
rect 3675 6358 3731 6392
rect 3765 6358 3821 6392
rect 3855 6358 3911 6392
rect 3945 6358 4001 6392
rect 4035 6358 4089 6392
rect 3409 6302 4089 6358
rect 3409 6268 3461 6302
rect 3495 6268 3551 6302
rect 3585 6268 3641 6302
rect 3675 6268 3731 6302
rect 3765 6268 3821 6302
rect 3855 6268 3911 6302
rect 3945 6268 4001 6302
rect 4035 6268 4089 6302
rect 3409 6212 4089 6268
rect 3409 6178 3461 6212
rect 3495 6178 3551 6212
rect 3585 6178 3641 6212
rect 3675 6178 3731 6212
rect 3765 6178 3821 6212
rect 3855 6178 3911 6212
rect 3945 6178 4001 6212
rect 4035 6178 4089 6212
rect 3409 6122 4089 6178
rect 3409 6088 3461 6122
rect 3495 6088 3551 6122
rect 3585 6088 3641 6122
rect 3675 6088 3731 6122
rect 3765 6088 3821 6122
rect 3855 6088 3911 6122
rect 3945 6088 4001 6122
rect 4035 6088 4089 6122
rect 3409 6034 4089 6088
rect 4797 6662 5477 6714
rect 4797 6628 4849 6662
rect 4883 6628 4939 6662
rect 4973 6628 5029 6662
rect 5063 6628 5119 6662
rect 5153 6628 5209 6662
rect 5243 6628 5299 6662
rect 5333 6628 5389 6662
rect 5423 6628 5477 6662
rect 4797 6572 5477 6628
rect 4797 6538 4849 6572
rect 4883 6538 4939 6572
rect 4973 6538 5029 6572
rect 5063 6538 5119 6572
rect 5153 6538 5209 6572
rect 5243 6538 5299 6572
rect 5333 6538 5389 6572
rect 5423 6538 5477 6572
rect 4797 6482 5477 6538
rect 4797 6448 4849 6482
rect 4883 6448 4939 6482
rect 4973 6448 5029 6482
rect 5063 6448 5119 6482
rect 5153 6448 5209 6482
rect 5243 6448 5299 6482
rect 5333 6448 5389 6482
rect 5423 6448 5477 6482
rect 4797 6392 5477 6448
rect 4797 6358 4849 6392
rect 4883 6358 4939 6392
rect 4973 6358 5029 6392
rect 5063 6358 5119 6392
rect 5153 6358 5209 6392
rect 5243 6358 5299 6392
rect 5333 6358 5389 6392
rect 5423 6358 5477 6392
rect 4797 6302 5477 6358
rect 4797 6268 4849 6302
rect 4883 6268 4939 6302
rect 4973 6268 5029 6302
rect 5063 6268 5119 6302
rect 5153 6268 5209 6302
rect 5243 6268 5299 6302
rect 5333 6268 5389 6302
rect 5423 6268 5477 6302
rect 4797 6212 5477 6268
rect 4797 6178 4849 6212
rect 4883 6178 4939 6212
rect 4973 6178 5029 6212
rect 5063 6178 5119 6212
rect 5153 6178 5209 6212
rect 5243 6178 5299 6212
rect 5333 6178 5389 6212
rect 5423 6178 5477 6212
rect 4797 6122 5477 6178
rect 4797 6088 4849 6122
rect 4883 6088 4939 6122
rect 4973 6088 5029 6122
rect 5063 6088 5119 6122
rect 5153 6088 5209 6122
rect 5243 6088 5299 6122
rect 5333 6088 5389 6122
rect 5423 6088 5477 6122
rect 4797 6034 5477 6088
rect 6185 6662 6865 6714
rect 6185 6628 6237 6662
rect 6271 6628 6327 6662
rect 6361 6628 6417 6662
rect 6451 6628 6507 6662
rect 6541 6628 6597 6662
rect 6631 6628 6687 6662
rect 6721 6628 6777 6662
rect 6811 6628 6865 6662
rect 6185 6572 6865 6628
rect 6185 6538 6237 6572
rect 6271 6538 6327 6572
rect 6361 6538 6417 6572
rect 6451 6538 6507 6572
rect 6541 6538 6597 6572
rect 6631 6538 6687 6572
rect 6721 6538 6777 6572
rect 6811 6538 6865 6572
rect 6185 6482 6865 6538
rect 6185 6448 6237 6482
rect 6271 6448 6327 6482
rect 6361 6448 6417 6482
rect 6451 6448 6507 6482
rect 6541 6448 6597 6482
rect 6631 6448 6687 6482
rect 6721 6448 6777 6482
rect 6811 6448 6865 6482
rect 6185 6392 6865 6448
rect 6185 6358 6237 6392
rect 6271 6358 6327 6392
rect 6361 6358 6417 6392
rect 6451 6358 6507 6392
rect 6541 6358 6597 6392
rect 6631 6358 6687 6392
rect 6721 6358 6777 6392
rect 6811 6358 6865 6392
rect 6185 6302 6865 6358
rect 6185 6268 6237 6302
rect 6271 6268 6327 6302
rect 6361 6268 6417 6302
rect 6451 6268 6507 6302
rect 6541 6268 6597 6302
rect 6631 6268 6687 6302
rect 6721 6268 6777 6302
rect 6811 6268 6865 6302
rect 6185 6212 6865 6268
rect 6185 6178 6237 6212
rect 6271 6178 6327 6212
rect 6361 6178 6417 6212
rect 6451 6178 6507 6212
rect 6541 6178 6597 6212
rect 6631 6178 6687 6212
rect 6721 6178 6777 6212
rect 6811 6178 6865 6212
rect 6185 6122 6865 6178
rect 6185 6088 6237 6122
rect 6271 6088 6327 6122
rect 6361 6088 6417 6122
rect 6451 6088 6507 6122
rect 6541 6088 6597 6122
rect 6631 6088 6687 6122
rect 6721 6088 6777 6122
rect 6811 6088 6865 6122
rect 6185 6034 6865 6088
rect 633 5274 1313 5326
rect 633 5240 685 5274
rect 719 5240 775 5274
rect 809 5240 865 5274
rect 899 5240 955 5274
rect 989 5240 1045 5274
rect 1079 5240 1135 5274
rect 1169 5240 1225 5274
rect 1259 5240 1313 5274
rect 633 5184 1313 5240
rect 633 5150 685 5184
rect 719 5150 775 5184
rect 809 5150 865 5184
rect 899 5150 955 5184
rect 989 5150 1045 5184
rect 1079 5150 1135 5184
rect 1169 5150 1225 5184
rect 1259 5150 1313 5184
rect 633 5094 1313 5150
rect 633 5060 685 5094
rect 719 5060 775 5094
rect 809 5060 865 5094
rect 899 5060 955 5094
rect 989 5060 1045 5094
rect 1079 5060 1135 5094
rect 1169 5060 1225 5094
rect 1259 5060 1313 5094
rect 633 5004 1313 5060
rect 633 4970 685 5004
rect 719 4970 775 5004
rect 809 4970 865 5004
rect 899 4970 955 5004
rect 989 4970 1045 5004
rect 1079 4970 1135 5004
rect 1169 4970 1225 5004
rect 1259 4970 1313 5004
rect 633 4914 1313 4970
rect 633 4880 685 4914
rect 719 4880 775 4914
rect 809 4880 865 4914
rect 899 4880 955 4914
rect 989 4880 1045 4914
rect 1079 4880 1135 4914
rect 1169 4880 1225 4914
rect 1259 4880 1313 4914
rect 633 4824 1313 4880
rect 633 4790 685 4824
rect 719 4790 775 4824
rect 809 4790 865 4824
rect 899 4790 955 4824
rect 989 4790 1045 4824
rect 1079 4790 1135 4824
rect 1169 4790 1225 4824
rect 1259 4790 1313 4824
rect 633 4734 1313 4790
rect 633 4700 685 4734
rect 719 4700 775 4734
rect 809 4700 865 4734
rect 899 4700 955 4734
rect 989 4700 1045 4734
rect 1079 4700 1135 4734
rect 1169 4700 1225 4734
rect 1259 4700 1313 4734
rect 633 4646 1313 4700
rect 2021 5274 2701 5326
rect 2021 5240 2073 5274
rect 2107 5240 2163 5274
rect 2197 5240 2253 5274
rect 2287 5240 2343 5274
rect 2377 5240 2433 5274
rect 2467 5240 2523 5274
rect 2557 5240 2613 5274
rect 2647 5240 2701 5274
rect 2021 5184 2701 5240
rect 2021 5150 2073 5184
rect 2107 5150 2163 5184
rect 2197 5150 2253 5184
rect 2287 5150 2343 5184
rect 2377 5150 2433 5184
rect 2467 5150 2523 5184
rect 2557 5150 2613 5184
rect 2647 5150 2701 5184
rect 2021 5094 2701 5150
rect 2021 5060 2073 5094
rect 2107 5060 2163 5094
rect 2197 5060 2253 5094
rect 2287 5060 2343 5094
rect 2377 5060 2433 5094
rect 2467 5060 2523 5094
rect 2557 5060 2613 5094
rect 2647 5060 2701 5094
rect 2021 5004 2701 5060
rect 2021 4970 2073 5004
rect 2107 4970 2163 5004
rect 2197 4970 2253 5004
rect 2287 4970 2343 5004
rect 2377 4970 2433 5004
rect 2467 4970 2523 5004
rect 2557 4970 2613 5004
rect 2647 4970 2701 5004
rect 2021 4914 2701 4970
rect 2021 4880 2073 4914
rect 2107 4880 2163 4914
rect 2197 4880 2253 4914
rect 2287 4880 2343 4914
rect 2377 4880 2433 4914
rect 2467 4880 2523 4914
rect 2557 4880 2613 4914
rect 2647 4880 2701 4914
rect 2021 4824 2701 4880
rect 2021 4790 2073 4824
rect 2107 4790 2163 4824
rect 2197 4790 2253 4824
rect 2287 4790 2343 4824
rect 2377 4790 2433 4824
rect 2467 4790 2523 4824
rect 2557 4790 2613 4824
rect 2647 4790 2701 4824
rect 2021 4734 2701 4790
rect 2021 4700 2073 4734
rect 2107 4700 2163 4734
rect 2197 4700 2253 4734
rect 2287 4700 2343 4734
rect 2377 4700 2433 4734
rect 2467 4700 2523 4734
rect 2557 4700 2613 4734
rect 2647 4700 2701 4734
rect 2021 4646 2701 4700
rect 3409 5274 4089 5326
rect 3409 5240 3461 5274
rect 3495 5240 3551 5274
rect 3585 5240 3641 5274
rect 3675 5240 3731 5274
rect 3765 5240 3821 5274
rect 3855 5240 3911 5274
rect 3945 5240 4001 5274
rect 4035 5240 4089 5274
rect 3409 5184 4089 5240
rect 3409 5150 3461 5184
rect 3495 5150 3551 5184
rect 3585 5150 3641 5184
rect 3675 5150 3731 5184
rect 3765 5150 3821 5184
rect 3855 5150 3911 5184
rect 3945 5150 4001 5184
rect 4035 5150 4089 5184
rect 3409 5094 4089 5150
rect 3409 5060 3461 5094
rect 3495 5060 3551 5094
rect 3585 5060 3641 5094
rect 3675 5060 3731 5094
rect 3765 5060 3821 5094
rect 3855 5060 3911 5094
rect 3945 5060 4001 5094
rect 4035 5060 4089 5094
rect 3409 5004 4089 5060
rect 3409 4970 3461 5004
rect 3495 4970 3551 5004
rect 3585 4970 3641 5004
rect 3675 4970 3731 5004
rect 3765 4970 3821 5004
rect 3855 4970 3911 5004
rect 3945 4970 4001 5004
rect 4035 4970 4089 5004
rect 3409 4914 4089 4970
rect 3409 4880 3461 4914
rect 3495 4880 3551 4914
rect 3585 4880 3641 4914
rect 3675 4880 3731 4914
rect 3765 4880 3821 4914
rect 3855 4880 3911 4914
rect 3945 4880 4001 4914
rect 4035 4880 4089 4914
rect 3409 4824 4089 4880
rect 3409 4790 3461 4824
rect 3495 4790 3551 4824
rect 3585 4790 3641 4824
rect 3675 4790 3731 4824
rect 3765 4790 3821 4824
rect 3855 4790 3911 4824
rect 3945 4790 4001 4824
rect 4035 4790 4089 4824
rect 3409 4734 4089 4790
rect 3409 4700 3461 4734
rect 3495 4700 3551 4734
rect 3585 4700 3641 4734
rect 3675 4700 3731 4734
rect 3765 4700 3821 4734
rect 3855 4700 3911 4734
rect 3945 4700 4001 4734
rect 4035 4700 4089 4734
rect 3409 4646 4089 4700
rect 4797 5274 5477 5326
rect 4797 5240 4849 5274
rect 4883 5240 4939 5274
rect 4973 5240 5029 5274
rect 5063 5240 5119 5274
rect 5153 5240 5209 5274
rect 5243 5240 5299 5274
rect 5333 5240 5389 5274
rect 5423 5240 5477 5274
rect 4797 5184 5477 5240
rect 4797 5150 4849 5184
rect 4883 5150 4939 5184
rect 4973 5150 5029 5184
rect 5063 5150 5119 5184
rect 5153 5150 5209 5184
rect 5243 5150 5299 5184
rect 5333 5150 5389 5184
rect 5423 5150 5477 5184
rect 4797 5094 5477 5150
rect 4797 5060 4849 5094
rect 4883 5060 4939 5094
rect 4973 5060 5029 5094
rect 5063 5060 5119 5094
rect 5153 5060 5209 5094
rect 5243 5060 5299 5094
rect 5333 5060 5389 5094
rect 5423 5060 5477 5094
rect 4797 5004 5477 5060
rect 4797 4970 4849 5004
rect 4883 4970 4939 5004
rect 4973 4970 5029 5004
rect 5063 4970 5119 5004
rect 5153 4970 5209 5004
rect 5243 4970 5299 5004
rect 5333 4970 5389 5004
rect 5423 4970 5477 5004
rect 4797 4914 5477 4970
rect 4797 4880 4849 4914
rect 4883 4880 4939 4914
rect 4973 4880 5029 4914
rect 5063 4880 5119 4914
rect 5153 4880 5209 4914
rect 5243 4880 5299 4914
rect 5333 4880 5389 4914
rect 5423 4880 5477 4914
rect 4797 4824 5477 4880
rect 4797 4790 4849 4824
rect 4883 4790 4939 4824
rect 4973 4790 5029 4824
rect 5063 4790 5119 4824
rect 5153 4790 5209 4824
rect 5243 4790 5299 4824
rect 5333 4790 5389 4824
rect 5423 4790 5477 4824
rect 4797 4734 5477 4790
rect 4797 4700 4849 4734
rect 4883 4700 4939 4734
rect 4973 4700 5029 4734
rect 5063 4700 5119 4734
rect 5153 4700 5209 4734
rect 5243 4700 5299 4734
rect 5333 4700 5389 4734
rect 5423 4700 5477 4734
rect 4797 4646 5477 4700
rect 6185 5274 6865 5326
rect 6185 5240 6237 5274
rect 6271 5240 6327 5274
rect 6361 5240 6417 5274
rect 6451 5240 6507 5274
rect 6541 5240 6597 5274
rect 6631 5240 6687 5274
rect 6721 5240 6777 5274
rect 6811 5240 6865 5274
rect 6185 5184 6865 5240
rect 6185 5150 6237 5184
rect 6271 5150 6327 5184
rect 6361 5150 6417 5184
rect 6451 5150 6507 5184
rect 6541 5150 6597 5184
rect 6631 5150 6687 5184
rect 6721 5150 6777 5184
rect 6811 5150 6865 5184
rect 6185 5094 6865 5150
rect 6185 5060 6237 5094
rect 6271 5060 6327 5094
rect 6361 5060 6417 5094
rect 6451 5060 6507 5094
rect 6541 5060 6597 5094
rect 6631 5060 6687 5094
rect 6721 5060 6777 5094
rect 6811 5060 6865 5094
rect 6185 5004 6865 5060
rect 6185 4970 6237 5004
rect 6271 4970 6327 5004
rect 6361 4970 6417 5004
rect 6451 4970 6507 5004
rect 6541 4970 6597 5004
rect 6631 4970 6687 5004
rect 6721 4970 6777 5004
rect 6811 4970 6865 5004
rect 6185 4914 6865 4970
rect 6185 4880 6237 4914
rect 6271 4880 6327 4914
rect 6361 4880 6417 4914
rect 6451 4880 6507 4914
rect 6541 4880 6597 4914
rect 6631 4880 6687 4914
rect 6721 4880 6777 4914
rect 6811 4880 6865 4914
rect 6185 4824 6865 4880
rect 6185 4790 6237 4824
rect 6271 4790 6327 4824
rect 6361 4790 6417 4824
rect 6451 4790 6507 4824
rect 6541 4790 6597 4824
rect 6631 4790 6687 4824
rect 6721 4790 6777 4824
rect 6811 4790 6865 4824
rect 6185 4734 6865 4790
rect 6185 4700 6237 4734
rect 6271 4700 6327 4734
rect 6361 4700 6417 4734
rect 6451 4700 6507 4734
rect 6541 4700 6597 4734
rect 6631 4700 6687 4734
rect 6721 4700 6777 4734
rect 6811 4700 6865 4734
rect 6185 4646 6865 4700
rect 633 3886 1313 3938
rect 633 3852 685 3886
rect 719 3852 775 3886
rect 809 3852 865 3886
rect 899 3852 955 3886
rect 989 3852 1045 3886
rect 1079 3852 1135 3886
rect 1169 3852 1225 3886
rect 1259 3852 1313 3886
rect 633 3796 1313 3852
rect 633 3762 685 3796
rect 719 3762 775 3796
rect 809 3762 865 3796
rect 899 3762 955 3796
rect 989 3762 1045 3796
rect 1079 3762 1135 3796
rect 1169 3762 1225 3796
rect 1259 3762 1313 3796
rect 633 3706 1313 3762
rect 633 3672 685 3706
rect 719 3672 775 3706
rect 809 3672 865 3706
rect 899 3672 955 3706
rect 989 3672 1045 3706
rect 1079 3672 1135 3706
rect 1169 3672 1225 3706
rect 1259 3672 1313 3706
rect 633 3616 1313 3672
rect 633 3582 685 3616
rect 719 3582 775 3616
rect 809 3582 865 3616
rect 899 3582 955 3616
rect 989 3582 1045 3616
rect 1079 3582 1135 3616
rect 1169 3582 1225 3616
rect 1259 3582 1313 3616
rect 633 3526 1313 3582
rect 633 3492 685 3526
rect 719 3492 775 3526
rect 809 3492 865 3526
rect 899 3492 955 3526
rect 989 3492 1045 3526
rect 1079 3492 1135 3526
rect 1169 3492 1225 3526
rect 1259 3492 1313 3526
rect 633 3436 1313 3492
rect 633 3402 685 3436
rect 719 3402 775 3436
rect 809 3402 865 3436
rect 899 3402 955 3436
rect 989 3402 1045 3436
rect 1079 3402 1135 3436
rect 1169 3402 1225 3436
rect 1259 3402 1313 3436
rect 633 3346 1313 3402
rect 633 3312 685 3346
rect 719 3312 775 3346
rect 809 3312 865 3346
rect 899 3312 955 3346
rect 989 3312 1045 3346
rect 1079 3312 1135 3346
rect 1169 3312 1225 3346
rect 1259 3312 1313 3346
rect 633 3258 1313 3312
rect 2021 3886 2701 3938
rect 2021 3852 2073 3886
rect 2107 3852 2163 3886
rect 2197 3852 2253 3886
rect 2287 3852 2343 3886
rect 2377 3852 2433 3886
rect 2467 3852 2523 3886
rect 2557 3852 2613 3886
rect 2647 3852 2701 3886
rect 2021 3796 2701 3852
rect 2021 3762 2073 3796
rect 2107 3762 2163 3796
rect 2197 3762 2253 3796
rect 2287 3762 2343 3796
rect 2377 3762 2433 3796
rect 2467 3762 2523 3796
rect 2557 3762 2613 3796
rect 2647 3762 2701 3796
rect 2021 3706 2701 3762
rect 2021 3672 2073 3706
rect 2107 3672 2163 3706
rect 2197 3672 2253 3706
rect 2287 3672 2343 3706
rect 2377 3672 2433 3706
rect 2467 3672 2523 3706
rect 2557 3672 2613 3706
rect 2647 3672 2701 3706
rect 2021 3616 2701 3672
rect 2021 3582 2073 3616
rect 2107 3582 2163 3616
rect 2197 3582 2253 3616
rect 2287 3582 2343 3616
rect 2377 3582 2433 3616
rect 2467 3582 2523 3616
rect 2557 3582 2613 3616
rect 2647 3582 2701 3616
rect 2021 3526 2701 3582
rect 2021 3492 2073 3526
rect 2107 3492 2163 3526
rect 2197 3492 2253 3526
rect 2287 3492 2343 3526
rect 2377 3492 2433 3526
rect 2467 3492 2523 3526
rect 2557 3492 2613 3526
rect 2647 3492 2701 3526
rect 2021 3436 2701 3492
rect 2021 3402 2073 3436
rect 2107 3402 2163 3436
rect 2197 3402 2253 3436
rect 2287 3402 2343 3436
rect 2377 3402 2433 3436
rect 2467 3402 2523 3436
rect 2557 3402 2613 3436
rect 2647 3402 2701 3436
rect 2021 3346 2701 3402
rect 2021 3312 2073 3346
rect 2107 3312 2163 3346
rect 2197 3312 2253 3346
rect 2287 3312 2343 3346
rect 2377 3312 2433 3346
rect 2467 3312 2523 3346
rect 2557 3312 2613 3346
rect 2647 3312 2701 3346
rect 2021 3258 2701 3312
rect 3409 3886 4089 3938
rect 3409 3852 3461 3886
rect 3495 3852 3551 3886
rect 3585 3852 3641 3886
rect 3675 3852 3731 3886
rect 3765 3852 3821 3886
rect 3855 3852 3911 3886
rect 3945 3852 4001 3886
rect 4035 3852 4089 3886
rect 3409 3796 4089 3852
rect 3409 3762 3461 3796
rect 3495 3762 3551 3796
rect 3585 3762 3641 3796
rect 3675 3762 3731 3796
rect 3765 3762 3821 3796
rect 3855 3762 3911 3796
rect 3945 3762 4001 3796
rect 4035 3762 4089 3796
rect 3409 3706 4089 3762
rect 3409 3672 3461 3706
rect 3495 3672 3551 3706
rect 3585 3672 3641 3706
rect 3675 3672 3731 3706
rect 3765 3672 3821 3706
rect 3855 3672 3911 3706
rect 3945 3672 4001 3706
rect 4035 3672 4089 3706
rect 3409 3616 4089 3672
rect 3409 3582 3461 3616
rect 3495 3582 3551 3616
rect 3585 3582 3641 3616
rect 3675 3582 3731 3616
rect 3765 3582 3821 3616
rect 3855 3582 3911 3616
rect 3945 3582 4001 3616
rect 4035 3582 4089 3616
rect 3409 3526 4089 3582
rect 3409 3492 3461 3526
rect 3495 3492 3551 3526
rect 3585 3492 3641 3526
rect 3675 3492 3731 3526
rect 3765 3492 3821 3526
rect 3855 3492 3911 3526
rect 3945 3492 4001 3526
rect 4035 3492 4089 3526
rect 3409 3436 4089 3492
rect 3409 3402 3461 3436
rect 3495 3402 3551 3436
rect 3585 3402 3641 3436
rect 3675 3402 3731 3436
rect 3765 3402 3821 3436
rect 3855 3402 3911 3436
rect 3945 3402 4001 3436
rect 4035 3402 4089 3436
rect 3409 3346 4089 3402
rect 3409 3312 3461 3346
rect 3495 3312 3551 3346
rect 3585 3312 3641 3346
rect 3675 3312 3731 3346
rect 3765 3312 3821 3346
rect 3855 3312 3911 3346
rect 3945 3312 4001 3346
rect 4035 3312 4089 3346
rect 3409 3258 4089 3312
rect 4797 3886 5477 3938
rect 4797 3852 4849 3886
rect 4883 3852 4939 3886
rect 4973 3852 5029 3886
rect 5063 3852 5119 3886
rect 5153 3852 5209 3886
rect 5243 3852 5299 3886
rect 5333 3852 5389 3886
rect 5423 3852 5477 3886
rect 4797 3796 5477 3852
rect 4797 3762 4849 3796
rect 4883 3762 4939 3796
rect 4973 3762 5029 3796
rect 5063 3762 5119 3796
rect 5153 3762 5209 3796
rect 5243 3762 5299 3796
rect 5333 3762 5389 3796
rect 5423 3762 5477 3796
rect 4797 3706 5477 3762
rect 4797 3672 4849 3706
rect 4883 3672 4939 3706
rect 4973 3672 5029 3706
rect 5063 3672 5119 3706
rect 5153 3672 5209 3706
rect 5243 3672 5299 3706
rect 5333 3672 5389 3706
rect 5423 3672 5477 3706
rect 4797 3616 5477 3672
rect 4797 3582 4849 3616
rect 4883 3582 4939 3616
rect 4973 3582 5029 3616
rect 5063 3582 5119 3616
rect 5153 3582 5209 3616
rect 5243 3582 5299 3616
rect 5333 3582 5389 3616
rect 5423 3582 5477 3616
rect 4797 3526 5477 3582
rect 4797 3492 4849 3526
rect 4883 3492 4939 3526
rect 4973 3492 5029 3526
rect 5063 3492 5119 3526
rect 5153 3492 5209 3526
rect 5243 3492 5299 3526
rect 5333 3492 5389 3526
rect 5423 3492 5477 3526
rect 4797 3436 5477 3492
rect 4797 3402 4849 3436
rect 4883 3402 4939 3436
rect 4973 3402 5029 3436
rect 5063 3402 5119 3436
rect 5153 3402 5209 3436
rect 5243 3402 5299 3436
rect 5333 3402 5389 3436
rect 5423 3402 5477 3436
rect 4797 3346 5477 3402
rect 4797 3312 4849 3346
rect 4883 3312 4939 3346
rect 4973 3312 5029 3346
rect 5063 3312 5119 3346
rect 5153 3312 5209 3346
rect 5243 3312 5299 3346
rect 5333 3312 5389 3346
rect 5423 3312 5477 3346
rect 4797 3258 5477 3312
rect 6185 3886 6865 3938
rect 6185 3852 6237 3886
rect 6271 3852 6327 3886
rect 6361 3852 6417 3886
rect 6451 3852 6507 3886
rect 6541 3852 6597 3886
rect 6631 3852 6687 3886
rect 6721 3852 6777 3886
rect 6811 3852 6865 3886
rect 6185 3796 6865 3852
rect 6185 3762 6237 3796
rect 6271 3762 6327 3796
rect 6361 3762 6417 3796
rect 6451 3762 6507 3796
rect 6541 3762 6597 3796
rect 6631 3762 6687 3796
rect 6721 3762 6777 3796
rect 6811 3762 6865 3796
rect 6185 3706 6865 3762
rect 6185 3672 6237 3706
rect 6271 3672 6327 3706
rect 6361 3672 6417 3706
rect 6451 3672 6507 3706
rect 6541 3672 6597 3706
rect 6631 3672 6687 3706
rect 6721 3672 6777 3706
rect 6811 3672 6865 3706
rect 6185 3616 6865 3672
rect 6185 3582 6237 3616
rect 6271 3582 6327 3616
rect 6361 3582 6417 3616
rect 6451 3582 6507 3616
rect 6541 3582 6597 3616
rect 6631 3582 6687 3616
rect 6721 3582 6777 3616
rect 6811 3582 6865 3616
rect 6185 3526 6865 3582
rect 6185 3492 6237 3526
rect 6271 3492 6327 3526
rect 6361 3492 6417 3526
rect 6451 3492 6507 3526
rect 6541 3492 6597 3526
rect 6631 3492 6687 3526
rect 6721 3492 6777 3526
rect 6811 3492 6865 3526
rect 6185 3436 6865 3492
rect 6185 3402 6237 3436
rect 6271 3402 6327 3436
rect 6361 3402 6417 3436
rect 6451 3402 6507 3436
rect 6541 3402 6597 3436
rect 6631 3402 6687 3436
rect 6721 3402 6777 3436
rect 6811 3402 6865 3436
rect 6185 3346 6865 3402
rect 6185 3312 6237 3346
rect 6271 3312 6327 3346
rect 6361 3312 6417 3346
rect 6451 3312 6507 3346
rect 6541 3312 6597 3346
rect 6631 3312 6687 3346
rect 6721 3312 6777 3346
rect 6811 3312 6865 3346
rect 6185 3258 6865 3312
rect 633 2498 1313 2550
rect 633 2464 685 2498
rect 719 2464 775 2498
rect 809 2464 865 2498
rect 899 2464 955 2498
rect 989 2464 1045 2498
rect 1079 2464 1135 2498
rect 1169 2464 1225 2498
rect 1259 2464 1313 2498
rect 633 2408 1313 2464
rect 633 2374 685 2408
rect 719 2374 775 2408
rect 809 2374 865 2408
rect 899 2374 955 2408
rect 989 2374 1045 2408
rect 1079 2374 1135 2408
rect 1169 2374 1225 2408
rect 1259 2374 1313 2408
rect 633 2318 1313 2374
rect 633 2284 685 2318
rect 719 2284 775 2318
rect 809 2284 865 2318
rect 899 2284 955 2318
rect 989 2284 1045 2318
rect 1079 2284 1135 2318
rect 1169 2284 1225 2318
rect 1259 2284 1313 2318
rect 633 2228 1313 2284
rect 633 2194 685 2228
rect 719 2194 775 2228
rect 809 2194 865 2228
rect 899 2194 955 2228
rect 989 2194 1045 2228
rect 1079 2194 1135 2228
rect 1169 2194 1225 2228
rect 1259 2194 1313 2228
rect 633 2138 1313 2194
rect 633 2104 685 2138
rect 719 2104 775 2138
rect 809 2104 865 2138
rect 899 2104 955 2138
rect 989 2104 1045 2138
rect 1079 2104 1135 2138
rect 1169 2104 1225 2138
rect 1259 2104 1313 2138
rect 633 2048 1313 2104
rect 633 2014 685 2048
rect 719 2014 775 2048
rect 809 2014 865 2048
rect 899 2014 955 2048
rect 989 2014 1045 2048
rect 1079 2014 1135 2048
rect 1169 2014 1225 2048
rect 1259 2014 1313 2048
rect 633 1958 1313 2014
rect 633 1924 685 1958
rect 719 1924 775 1958
rect 809 1924 865 1958
rect 899 1924 955 1958
rect 989 1924 1045 1958
rect 1079 1924 1135 1958
rect 1169 1924 1225 1958
rect 1259 1924 1313 1958
rect 633 1870 1313 1924
rect 2021 2498 2701 2550
rect 2021 2464 2073 2498
rect 2107 2464 2163 2498
rect 2197 2464 2253 2498
rect 2287 2464 2343 2498
rect 2377 2464 2433 2498
rect 2467 2464 2523 2498
rect 2557 2464 2613 2498
rect 2647 2464 2701 2498
rect 2021 2408 2701 2464
rect 2021 2374 2073 2408
rect 2107 2374 2163 2408
rect 2197 2374 2253 2408
rect 2287 2374 2343 2408
rect 2377 2374 2433 2408
rect 2467 2374 2523 2408
rect 2557 2374 2613 2408
rect 2647 2374 2701 2408
rect 2021 2318 2701 2374
rect 2021 2284 2073 2318
rect 2107 2284 2163 2318
rect 2197 2284 2253 2318
rect 2287 2284 2343 2318
rect 2377 2284 2433 2318
rect 2467 2284 2523 2318
rect 2557 2284 2613 2318
rect 2647 2284 2701 2318
rect 2021 2228 2701 2284
rect 2021 2194 2073 2228
rect 2107 2194 2163 2228
rect 2197 2194 2253 2228
rect 2287 2194 2343 2228
rect 2377 2194 2433 2228
rect 2467 2194 2523 2228
rect 2557 2194 2613 2228
rect 2647 2194 2701 2228
rect 2021 2138 2701 2194
rect 2021 2104 2073 2138
rect 2107 2104 2163 2138
rect 2197 2104 2253 2138
rect 2287 2104 2343 2138
rect 2377 2104 2433 2138
rect 2467 2104 2523 2138
rect 2557 2104 2613 2138
rect 2647 2104 2701 2138
rect 2021 2048 2701 2104
rect 2021 2014 2073 2048
rect 2107 2014 2163 2048
rect 2197 2014 2253 2048
rect 2287 2014 2343 2048
rect 2377 2014 2433 2048
rect 2467 2014 2523 2048
rect 2557 2014 2613 2048
rect 2647 2014 2701 2048
rect 2021 1958 2701 2014
rect 2021 1924 2073 1958
rect 2107 1924 2163 1958
rect 2197 1924 2253 1958
rect 2287 1924 2343 1958
rect 2377 1924 2433 1958
rect 2467 1924 2523 1958
rect 2557 1924 2613 1958
rect 2647 1924 2701 1958
rect 2021 1870 2701 1924
rect 3409 2498 4089 2550
rect 3409 2464 3461 2498
rect 3495 2464 3551 2498
rect 3585 2464 3641 2498
rect 3675 2464 3731 2498
rect 3765 2464 3821 2498
rect 3855 2464 3911 2498
rect 3945 2464 4001 2498
rect 4035 2464 4089 2498
rect 3409 2408 4089 2464
rect 3409 2374 3461 2408
rect 3495 2374 3551 2408
rect 3585 2374 3641 2408
rect 3675 2374 3731 2408
rect 3765 2374 3821 2408
rect 3855 2374 3911 2408
rect 3945 2374 4001 2408
rect 4035 2374 4089 2408
rect 3409 2318 4089 2374
rect 3409 2284 3461 2318
rect 3495 2284 3551 2318
rect 3585 2284 3641 2318
rect 3675 2284 3731 2318
rect 3765 2284 3821 2318
rect 3855 2284 3911 2318
rect 3945 2284 4001 2318
rect 4035 2284 4089 2318
rect 3409 2228 4089 2284
rect 3409 2194 3461 2228
rect 3495 2194 3551 2228
rect 3585 2194 3641 2228
rect 3675 2194 3731 2228
rect 3765 2194 3821 2228
rect 3855 2194 3911 2228
rect 3945 2194 4001 2228
rect 4035 2194 4089 2228
rect 3409 2138 4089 2194
rect 3409 2104 3461 2138
rect 3495 2104 3551 2138
rect 3585 2104 3641 2138
rect 3675 2104 3731 2138
rect 3765 2104 3821 2138
rect 3855 2104 3911 2138
rect 3945 2104 4001 2138
rect 4035 2104 4089 2138
rect 3409 2048 4089 2104
rect 3409 2014 3461 2048
rect 3495 2014 3551 2048
rect 3585 2014 3641 2048
rect 3675 2014 3731 2048
rect 3765 2014 3821 2048
rect 3855 2014 3911 2048
rect 3945 2014 4001 2048
rect 4035 2014 4089 2048
rect 3409 1958 4089 2014
rect 3409 1924 3461 1958
rect 3495 1924 3551 1958
rect 3585 1924 3641 1958
rect 3675 1924 3731 1958
rect 3765 1924 3821 1958
rect 3855 1924 3911 1958
rect 3945 1924 4001 1958
rect 4035 1924 4089 1958
rect 3409 1870 4089 1924
rect 4797 2498 5477 2550
rect 4797 2464 4849 2498
rect 4883 2464 4939 2498
rect 4973 2464 5029 2498
rect 5063 2464 5119 2498
rect 5153 2464 5209 2498
rect 5243 2464 5299 2498
rect 5333 2464 5389 2498
rect 5423 2464 5477 2498
rect 4797 2408 5477 2464
rect 4797 2374 4849 2408
rect 4883 2374 4939 2408
rect 4973 2374 5029 2408
rect 5063 2374 5119 2408
rect 5153 2374 5209 2408
rect 5243 2374 5299 2408
rect 5333 2374 5389 2408
rect 5423 2374 5477 2408
rect 4797 2318 5477 2374
rect 4797 2284 4849 2318
rect 4883 2284 4939 2318
rect 4973 2284 5029 2318
rect 5063 2284 5119 2318
rect 5153 2284 5209 2318
rect 5243 2284 5299 2318
rect 5333 2284 5389 2318
rect 5423 2284 5477 2318
rect 4797 2228 5477 2284
rect 4797 2194 4849 2228
rect 4883 2194 4939 2228
rect 4973 2194 5029 2228
rect 5063 2194 5119 2228
rect 5153 2194 5209 2228
rect 5243 2194 5299 2228
rect 5333 2194 5389 2228
rect 5423 2194 5477 2228
rect 4797 2138 5477 2194
rect 4797 2104 4849 2138
rect 4883 2104 4939 2138
rect 4973 2104 5029 2138
rect 5063 2104 5119 2138
rect 5153 2104 5209 2138
rect 5243 2104 5299 2138
rect 5333 2104 5389 2138
rect 5423 2104 5477 2138
rect 4797 2048 5477 2104
rect 4797 2014 4849 2048
rect 4883 2014 4939 2048
rect 4973 2014 5029 2048
rect 5063 2014 5119 2048
rect 5153 2014 5209 2048
rect 5243 2014 5299 2048
rect 5333 2014 5389 2048
rect 5423 2014 5477 2048
rect 4797 1958 5477 2014
rect 4797 1924 4849 1958
rect 4883 1924 4939 1958
rect 4973 1924 5029 1958
rect 5063 1924 5119 1958
rect 5153 1924 5209 1958
rect 5243 1924 5299 1958
rect 5333 1924 5389 1958
rect 5423 1924 5477 1958
rect 4797 1870 5477 1924
rect 6185 2498 6865 2550
rect 6185 2464 6237 2498
rect 6271 2464 6327 2498
rect 6361 2464 6417 2498
rect 6451 2464 6507 2498
rect 6541 2464 6597 2498
rect 6631 2464 6687 2498
rect 6721 2464 6777 2498
rect 6811 2464 6865 2498
rect 6185 2408 6865 2464
rect 6185 2374 6237 2408
rect 6271 2374 6327 2408
rect 6361 2374 6417 2408
rect 6451 2374 6507 2408
rect 6541 2374 6597 2408
rect 6631 2374 6687 2408
rect 6721 2374 6777 2408
rect 6811 2374 6865 2408
rect 6185 2318 6865 2374
rect 6185 2284 6237 2318
rect 6271 2284 6327 2318
rect 6361 2284 6417 2318
rect 6451 2284 6507 2318
rect 6541 2284 6597 2318
rect 6631 2284 6687 2318
rect 6721 2284 6777 2318
rect 6811 2284 6865 2318
rect 6185 2228 6865 2284
rect 6185 2194 6237 2228
rect 6271 2194 6327 2228
rect 6361 2194 6417 2228
rect 6451 2194 6507 2228
rect 6541 2194 6597 2228
rect 6631 2194 6687 2228
rect 6721 2194 6777 2228
rect 6811 2194 6865 2228
rect 6185 2138 6865 2194
rect 6185 2104 6237 2138
rect 6271 2104 6327 2138
rect 6361 2104 6417 2138
rect 6451 2104 6507 2138
rect 6541 2104 6597 2138
rect 6631 2104 6687 2138
rect 6721 2104 6777 2138
rect 6811 2104 6865 2138
rect 6185 2048 6865 2104
rect 6185 2014 6237 2048
rect 6271 2014 6327 2048
rect 6361 2014 6417 2048
rect 6451 2014 6507 2048
rect 6541 2014 6597 2048
rect 6631 2014 6687 2048
rect 6721 2014 6777 2048
rect 6811 2014 6865 2048
rect 6185 1958 6865 2014
rect 6185 1924 6237 1958
rect 6271 1924 6327 1958
rect 6361 1924 6417 1958
rect 6451 1924 6507 1958
rect 6541 1924 6597 1958
rect 6631 1924 6687 1958
rect 6721 1924 6777 1958
rect 6811 1924 6865 1958
rect 6185 1870 6865 1924
<< ndiffc >>
rect -1170 17264 -1136 17440
rect -1082 17264 -1048 17440
rect -824 17264 -790 17440
rect -566 17264 -532 17440
rect -478 17264 -444 17440
rect -1170 16954 -1136 17130
rect -1082 16954 -1048 17130
rect -824 16954 -790 17130
rect -566 16954 -532 17130
rect -478 16954 -444 17130
rect -92 17276 -58 17452
rect -4 17276 30 17452
rect 108 17276 142 17452
rect 4166 17276 4200 17452
rect 4278 17276 4312 17452
rect 8336 17276 8370 17452
rect 8448 17276 8482 17452
rect 8536 17276 8570 17452
rect -92 16882 -58 17058
rect -4 16882 30 17058
rect 108 16882 142 17058
rect 4166 16882 4200 17058
rect 4278 16882 4312 17058
rect 8336 16882 8370 17058
rect 8448 16882 8482 17058
rect 8536 16882 8570 17058
rect -92 16488 -58 16664
rect -4 16488 30 16664
rect 108 16488 142 16664
rect 4166 16488 4200 16664
rect 4278 16488 4312 16664
rect 8336 16488 8370 16664
rect 8448 16488 8482 16664
rect 8536 16488 8570 16664
rect -92 16094 -58 16270
rect -4 16094 30 16270
rect 108 16094 142 16270
rect 4166 16094 4200 16270
rect 4278 16094 4312 16270
rect 8336 16094 8370 16270
rect 8448 16094 8482 16270
rect 8536 16094 8570 16270
rect 3013 15378 3047 15534
rect 3101 15378 3135 15534
rect 5759 15378 5793 15534
rect 8417 15378 8451 15534
rect 8505 15378 8539 15534
rect 3013 14946 3047 15102
rect 3101 14946 3135 15102
rect 5759 14946 5793 15102
rect 8417 14946 8451 15102
rect 8505 14946 8539 15102
rect 704 11390 738 12166
rect 792 11390 826 12166
rect 1050 11390 1084 12166
rect 1308 11390 1342 12166
rect 1396 11390 1430 12166
rect 704 10396 738 11172
rect 792 10396 826 11172
rect 1050 10396 1084 11172
rect 1308 10396 1342 11172
rect 1396 10396 1430 11172
rect 1596 11390 1630 12166
rect 1684 11390 1718 12166
rect 1942 11390 1976 12166
rect 2200 11390 2234 12166
rect 2288 11390 2322 12166
rect 1596 10396 1630 11172
rect 1684 10396 1718 11172
rect 1942 10396 1976 11172
rect 2200 10396 2234 11172
rect 2288 10396 2322 11172
rect 2488 11390 2522 12166
rect 2576 11390 2610 12166
rect 2834 11390 2868 12166
rect 3092 11390 3126 12166
rect 3180 11390 3214 12166
rect 2488 10396 2522 11172
rect 2576 10396 2610 11172
rect 2834 10396 2868 11172
rect 3092 10396 3126 11172
rect 3180 10396 3214 11172
rect 3380 11390 3414 12166
rect 3468 11390 3502 12166
rect 3726 11390 3760 12166
rect 3984 11390 4018 12166
rect 4072 11390 4106 12166
rect 3380 10396 3414 11172
rect 3468 10396 3502 11172
rect 3726 10396 3760 11172
rect 3984 10396 4018 11172
rect 4072 10396 4106 11172
rect 4428 12167 4604 12201
rect 4428 12079 4604 12113
rect 4428 11821 4604 11855
rect 4428 11563 4604 11597
rect 4428 11475 4604 11509
rect 4428 11053 4604 11087
rect 4428 10965 4604 10999
rect 4428 10707 4604 10741
rect 4428 10449 4604 10483
rect 4428 10361 4604 10395
<< pdiffc >>
rect -16517 17278 -16483 17454
rect -16429 17278 -16395 17454
rect -14371 17278 -14337 17454
rect -12313 17278 -12279 17454
rect -10255 17278 -10221 17454
rect -8197 17278 -8163 17454
rect -8109 17278 -8075 17454
rect -16517 16799 -16483 16975
rect -16429 16799 -16395 16975
rect -14371 16799 -14337 16975
rect -12313 16799 -12279 16975
rect -10255 16799 -10221 16975
rect -8197 16799 -8163 16975
rect -8109 16799 -8075 16975
rect -16517 16329 -16483 16505
rect -16429 16329 -16395 16505
rect -14371 16329 -14337 16505
rect -12313 16329 -12279 16505
rect -10255 16329 -10221 16505
rect -8197 16329 -8163 16505
rect -8109 16329 -8075 16505
rect -16517 15850 -16483 16026
rect -16429 15850 -16395 16026
rect -14371 15850 -14337 16026
rect -12313 15850 -12279 16026
rect -10255 15850 -10221 16026
rect -8197 15850 -8163 16026
rect -8109 15850 -8075 16026
rect -7496 17184 -7462 17360
rect -7408 17184 -7374 17360
rect -5350 17184 -5316 17360
rect -3292 17184 -3258 17360
rect -3204 17184 -3170 17360
rect -7496 16752 -7462 16928
rect -7408 16752 -7374 16928
rect -5350 16752 -5316 16928
rect -3292 16752 -3258 16928
rect -3204 16752 -3170 16928
rect -7496 16282 -7462 16458
rect -7408 16282 -7374 16458
rect -5350 16282 -5316 16458
rect -3292 16282 -3258 16458
rect -3204 16282 -3170 16458
rect -7496 15850 -7462 16026
rect -7408 15850 -7374 16026
rect -5350 15850 -5316 16026
rect -3292 15850 -3258 16026
rect -3204 15850 -3170 16026
rect -12368 15236 -12334 15412
rect -12280 15236 -12246 15412
rect -10222 15236 -10188 15412
rect -8164 15236 -8130 15412
rect -8076 15236 -8042 15412
rect -12368 14842 -12334 15018
rect -12280 14842 -12246 15018
rect -10222 14842 -10188 15018
rect -8164 14842 -8130 15018
rect -8076 14842 -8042 15018
rect -7462 15301 -7428 15477
rect -7374 15301 -7340 15477
rect -5316 15301 -5282 15477
rect -3258 15301 -3224 15477
rect -3170 15301 -3136 15477
rect -7462 14825 -7428 15001
rect -7374 14825 -7340 15001
rect -5316 14825 -5282 15001
rect -3258 14825 -3224 15001
rect -3170 14825 -3136 15001
rect 5001 11778 5377 11812
rect 5595 11778 5971 11812
rect 5001 11690 5377 11724
rect 5595 11690 5971 11724
rect 5001 11232 5377 11266
rect 5595 11232 5971 11266
rect 5001 10774 5377 10808
rect 5595 10774 5971 10808
rect 5001 10686 5377 10720
rect 5595 10686 5971 10720
rect 685 8016 719 8050
rect 775 8016 809 8050
rect 865 8016 899 8050
rect 955 8016 989 8050
rect 1045 8016 1079 8050
rect 1135 8016 1169 8050
rect 1225 8016 1259 8050
rect 685 7926 719 7960
rect 775 7926 809 7960
rect 865 7926 899 7960
rect 955 7926 989 7960
rect 1045 7926 1079 7960
rect 1135 7926 1169 7960
rect 1225 7926 1259 7960
rect 685 7836 719 7870
rect 775 7836 809 7870
rect 865 7836 899 7870
rect 955 7836 989 7870
rect 1045 7836 1079 7870
rect 1135 7836 1169 7870
rect 1225 7836 1259 7870
rect 685 7746 719 7780
rect 775 7746 809 7780
rect 865 7746 899 7780
rect 955 7746 989 7780
rect 1045 7746 1079 7780
rect 1135 7746 1169 7780
rect 1225 7746 1259 7780
rect 685 7656 719 7690
rect 775 7656 809 7690
rect 865 7656 899 7690
rect 955 7656 989 7690
rect 1045 7656 1079 7690
rect 1135 7656 1169 7690
rect 1225 7656 1259 7690
rect 685 7566 719 7600
rect 775 7566 809 7600
rect 865 7566 899 7600
rect 955 7566 989 7600
rect 1045 7566 1079 7600
rect 1135 7566 1169 7600
rect 1225 7566 1259 7600
rect 685 7476 719 7510
rect 775 7476 809 7510
rect 865 7476 899 7510
rect 955 7476 989 7510
rect 1045 7476 1079 7510
rect 1135 7476 1169 7510
rect 1225 7476 1259 7510
rect 2073 8016 2107 8050
rect 2163 8016 2197 8050
rect 2253 8016 2287 8050
rect 2343 8016 2377 8050
rect 2433 8016 2467 8050
rect 2523 8016 2557 8050
rect 2613 8016 2647 8050
rect 2073 7926 2107 7960
rect 2163 7926 2197 7960
rect 2253 7926 2287 7960
rect 2343 7926 2377 7960
rect 2433 7926 2467 7960
rect 2523 7926 2557 7960
rect 2613 7926 2647 7960
rect 2073 7836 2107 7870
rect 2163 7836 2197 7870
rect 2253 7836 2287 7870
rect 2343 7836 2377 7870
rect 2433 7836 2467 7870
rect 2523 7836 2557 7870
rect 2613 7836 2647 7870
rect 2073 7746 2107 7780
rect 2163 7746 2197 7780
rect 2253 7746 2287 7780
rect 2343 7746 2377 7780
rect 2433 7746 2467 7780
rect 2523 7746 2557 7780
rect 2613 7746 2647 7780
rect 2073 7656 2107 7690
rect 2163 7656 2197 7690
rect 2253 7656 2287 7690
rect 2343 7656 2377 7690
rect 2433 7656 2467 7690
rect 2523 7656 2557 7690
rect 2613 7656 2647 7690
rect 2073 7566 2107 7600
rect 2163 7566 2197 7600
rect 2253 7566 2287 7600
rect 2343 7566 2377 7600
rect 2433 7566 2467 7600
rect 2523 7566 2557 7600
rect 2613 7566 2647 7600
rect 2073 7476 2107 7510
rect 2163 7476 2197 7510
rect 2253 7476 2287 7510
rect 2343 7476 2377 7510
rect 2433 7476 2467 7510
rect 2523 7476 2557 7510
rect 2613 7476 2647 7510
rect 3461 8016 3495 8050
rect 3551 8016 3585 8050
rect 3641 8016 3675 8050
rect 3731 8016 3765 8050
rect 3821 8016 3855 8050
rect 3911 8016 3945 8050
rect 4001 8016 4035 8050
rect 3461 7926 3495 7960
rect 3551 7926 3585 7960
rect 3641 7926 3675 7960
rect 3731 7926 3765 7960
rect 3821 7926 3855 7960
rect 3911 7926 3945 7960
rect 4001 7926 4035 7960
rect 3461 7836 3495 7870
rect 3551 7836 3585 7870
rect 3641 7836 3675 7870
rect 3731 7836 3765 7870
rect 3821 7836 3855 7870
rect 3911 7836 3945 7870
rect 4001 7836 4035 7870
rect 3461 7746 3495 7780
rect 3551 7746 3585 7780
rect 3641 7746 3675 7780
rect 3731 7746 3765 7780
rect 3821 7746 3855 7780
rect 3911 7746 3945 7780
rect 4001 7746 4035 7780
rect 3461 7656 3495 7690
rect 3551 7656 3585 7690
rect 3641 7656 3675 7690
rect 3731 7656 3765 7690
rect 3821 7656 3855 7690
rect 3911 7656 3945 7690
rect 4001 7656 4035 7690
rect 3461 7566 3495 7600
rect 3551 7566 3585 7600
rect 3641 7566 3675 7600
rect 3731 7566 3765 7600
rect 3821 7566 3855 7600
rect 3911 7566 3945 7600
rect 4001 7566 4035 7600
rect 3461 7476 3495 7510
rect 3551 7476 3585 7510
rect 3641 7476 3675 7510
rect 3731 7476 3765 7510
rect 3821 7476 3855 7510
rect 3911 7476 3945 7510
rect 4001 7476 4035 7510
rect 4849 8016 4883 8050
rect 4939 8016 4973 8050
rect 5029 8016 5063 8050
rect 5119 8016 5153 8050
rect 5209 8016 5243 8050
rect 5299 8016 5333 8050
rect 5389 8016 5423 8050
rect 4849 7926 4883 7960
rect 4939 7926 4973 7960
rect 5029 7926 5063 7960
rect 5119 7926 5153 7960
rect 5209 7926 5243 7960
rect 5299 7926 5333 7960
rect 5389 7926 5423 7960
rect 4849 7836 4883 7870
rect 4939 7836 4973 7870
rect 5029 7836 5063 7870
rect 5119 7836 5153 7870
rect 5209 7836 5243 7870
rect 5299 7836 5333 7870
rect 5389 7836 5423 7870
rect 4849 7746 4883 7780
rect 4939 7746 4973 7780
rect 5029 7746 5063 7780
rect 5119 7746 5153 7780
rect 5209 7746 5243 7780
rect 5299 7746 5333 7780
rect 5389 7746 5423 7780
rect 4849 7656 4883 7690
rect 4939 7656 4973 7690
rect 5029 7656 5063 7690
rect 5119 7656 5153 7690
rect 5209 7656 5243 7690
rect 5299 7656 5333 7690
rect 5389 7656 5423 7690
rect 4849 7566 4883 7600
rect 4939 7566 4973 7600
rect 5029 7566 5063 7600
rect 5119 7566 5153 7600
rect 5209 7566 5243 7600
rect 5299 7566 5333 7600
rect 5389 7566 5423 7600
rect 4849 7476 4883 7510
rect 4939 7476 4973 7510
rect 5029 7476 5063 7510
rect 5119 7476 5153 7510
rect 5209 7476 5243 7510
rect 5299 7476 5333 7510
rect 5389 7476 5423 7510
rect 6237 8016 6271 8050
rect 6327 8016 6361 8050
rect 6417 8016 6451 8050
rect 6507 8016 6541 8050
rect 6597 8016 6631 8050
rect 6687 8016 6721 8050
rect 6777 8016 6811 8050
rect 6237 7926 6271 7960
rect 6327 7926 6361 7960
rect 6417 7926 6451 7960
rect 6507 7926 6541 7960
rect 6597 7926 6631 7960
rect 6687 7926 6721 7960
rect 6777 7926 6811 7960
rect 6237 7836 6271 7870
rect 6327 7836 6361 7870
rect 6417 7836 6451 7870
rect 6507 7836 6541 7870
rect 6597 7836 6631 7870
rect 6687 7836 6721 7870
rect 6777 7836 6811 7870
rect 6237 7746 6271 7780
rect 6327 7746 6361 7780
rect 6417 7746 6451 7780
rect 6507 7746 6541 7780
rect 6597 7746 6631 7780
rect 6687 7746 6721 7780
rect 6777 7746 6811 7780
rect 6237 7656 6271 7690
rect 6327 7656 6361 7690
rect 6417 7656 6451 7690
rect 6507 7656 6541 7690
rect 6597 7656 6631 7690
rect 6687 7656 6721 7690
rect 6777 7656 6811 7690
rect 6237 7566 6271 7600
rect 6327 7566 6361 7600
rect 6417 7566 6451 7600
rect 6507 7566 6541 7600
rect 6597 7566 6631 7600
rect 6687 7566 6721 7600
rect 6777 7566 6811 7600
rect 6237 7476 6271 7510
rect 6327 7476 6361 7510
rect 6417 7476 6451 7510
rect 6507 7476 6541 7510
rect 6597 7476 6631 7510
rect 6687 7476 6721 7510
rect 6777 7476 6811 7510
rect 685 6628 719 6662
rect 775 6628 809 6662
rect 865 6628 899 6662
rect 955 6628 989 6662
rect 1045 6628 1079 6662
rect 1135 6628 1169 6662
rect 1225 6628 1259 6662
rect 685 6538 719 6572
rect 775 6538 809 6572
rect 865 6538 899 6572
rect 955 6538 989 6572
rect 1045 6538 1079 6572
rect 1135 6538 1169 6572
rect 1225 6538 1259 6572
rect 685 6448 719 6482
rect 775 6448 809 6482
rect 865 6448 899 6482
rect 955 6448 989 6482
rect 1045 6448 1079 6482
rect 1135 6448 1169 6482
rect 1225 6448 1259 6482
rect 685 6358 719 6392
rect 775 6358 809 6392
rect 865 6358 899 6392
rect 955 6358 989 6392
rect 1045 6358 1079 6392
rect 1135 6358 1169 6392
rect 1225 6358 1259 6392
rect 685 6268 719 6302
rect 775 6268 809 6302
rect 865 6268 899 6302
rect 955 6268 989 6302
rect 1045 6268 1079 6302
rect 1135 6268 1169 6302
rect 1225 6268 1259 6302
rect 685 6178 719 6212
rect 775 6178 809 6212
rect 865 6178 899 6212
rect 955 6178 989 6212
rect 1045 6178 1079 6212
rect 1135 6178 1169 6212
rect 1225 6178 1259 6212
rect 685 6088 719 6122
rect 775 6088 809 6122
rect 865 6088 899 6122
rect 955 6088 989 6122
rect 1045 6088 1079 6122
rect 1135 6088 1169 6122
rect 1225 6088 1259 6122
rect 2073 6628 2107 6662
rect 2163 6628 2197 6662
rect 2253 6628 2287 6662
rect 2343 6628 2377 6662
rect 2433 6628 2467 6662
rect 2523 6628 2557 6662
rect 2613 6628 2647 6662
rect 2073 6538 2107 6572
rect 2163 6538 2197 6572
rect 2253 6538 2287 6572
rect 2343 6538 2377 6572
rect 2433 6538 2467 6572
rect 2523 6538 2557 6572
rect 2613 6538 2647 6572
rect 2073 6448 2107 6482
rect 2163 6448 2197 6482
rect 2253 6448 2287 6482
rect 2343 6448 2377 6482
rect 2433 6448 2467 6482
rect 2523 6448 2557 6482
rect 2613 6448 2647 6482
rect 2073 6358 2107 6392
rect 2163 6358 2197 6392
rect 2253 6358 2287 6392
rect 2343 6358 2377 6392
rect 2433 6358 2467 6392
rect 2523 6358 2557 6392
rect 2613 6358 2647 6392
rect 2073 6268 2107 6302
rect 2163 6268 2197 6302
rect 2253 6268 2287 6302
rect 2343 6268 2377 6302
rect 2433 6268 2467 6302
rect 2523 6268 2557 6302
rect 2613 6268 2647 6302
rect 2073 6178 2107 6212
rect 2163 6178 2197 6212
rect 2253 6178 2287 6212
rect 2343 6178 2377 6212
rect 2433 6178 2467 6212
rect 2523 6178 2557 6212
rect 2613 6178 2647 6212
rect 2073 6088 2107 6122
rect 2163 6088 2197 6122
rect 2253 6088 2287 6122
rect 2343 6088 2377 6122
rect 2433 6088 2467 6122
rect 2523 6088 2557 6122
rect 2613 6088 2647 6122
rect 3461 6628 3495 6662
rect 3551 6628 3585 6662
rect 3641 6628 3675 6662
rect 3731 6628 3765 6662
rect 3821 6628 3855 6662
rect 3911 6628 3945 6662
rect 4001 6628 4035 6662
rect 3461 6538 3495 6572
rect 3551 6538 3585 6572
rect 3641 6538 3675 6572
rect 3731 6538 3765 6572
rect 3821 6538 3855 6572
rect 3911 6538 3945 6572
rect 4001 6538 4035 6572
rect 3461 6448 3495 6482
rect 3551 6448 3585 6482
rect 3641 6448 3675 6482
rect 3731 6448 3765 6482
rect 3821 6448 3855 6482
rect 3911 6448 3945 6482
rect 4001 6448 4035 6482
rect 3461 6358 3495 6392
rect 3551 6358 3585 6392
rect 3641 6358 3675 6392
rect 3731 6358 3765 6392
rect 3821 6358 3855 6392
rect 3911 6358 3945 6392
rect 4001 6358 4035 6392
rect 3461 6268 3495 6302
rect 3551 6268 3585 6302
rect 3641 6268 3675 6302
rect 3731 6268 3765 6302
rect 3821 6268 3855 6302
rect 3911 6268 3945 6302
rect 4001 6268 4035 6302
rect 3461 6178 3495 6212
rect 3551 6178 3585 6212
rect 3641 6178 3675 6212
rect 3731 6178 3765 6212
rect 3821 6178 3855 6212
rect 3911 6178 3945 6212
rect 4001 6178 4035 6212
rect 3461 6088 3495 6122
rect 3551 6088 3585 6122
rect 3641 6088 3675 6122
rect 3731 6088 3765 6122
rect 3821 6088 3855 6122
rect 3911 6088 3945 6122
rect 4001 6088 4035 6122
rect 4849 6628 4883 6662
rect 4939 6628 4973 6662
rect 5029 6628 5063 6662
rect 5119 6628 5153 6662
rect 5209 6628 5243 6662
rect 5299 6628 5333 6662
rect 5389 6628 5423 6662
rect 4849 6538 4883 6572
rect 4939 6538 4973 6572
rect 5029 6538 5063 6572
rect 5119 6538 5153 6572
rect 5209 6538 5243 6572
rect 5299 6538 5333 6572
rect 5389 6538 5423 6572
rect 4849 6448 4883 6482
rect 4939 6448 4973 6482
rect 5029 6448 5063 6482
rect 5119 6448 5153 6482
rect 5209 6448 5243 6482
rect 5299 6448 5333 6482
rect 5389 6448 5423 6482
rect 4849 6358 4883 6392
rect 4939 6358 4973 6392
rect 5029 6358 5063 6392
rect 5119 6358 5153 6392
rect 5209 6358 5243 6392
rect 5299 6358 5333 6392
rect 5389 6358 5423 6392
rect 4849 6268 4883 6302
rect 4939 6268 4973 6302
rect 5029 6268 5063 6302
rect 5119 6268 5153 6302
rect 5209 6268 5243 6302
rect 5299 6268 5333 6302
rect 5389 6268 5423 6302
rect 4849 6178 4883 6212
rect 4939 6178 4973 6212
rect 5029 6178 5063 6212
rect 5119 6178 5153 6212
rect 5209 6178 5243 6212
rect 5299 6178 5333 6212
rect 5389 6178 5423 6212
rect 4849 6088 4883 6122
rect 4939 6088 4973 6122
rect 5029 6088 5063 6122
rect 5119 6088 5153 6122
rect 5209 6088 5243 6122
rect 5299 6088 5333 6122
rect 5389 6088 5423 6122
rect 6237 6628 6271 6662
rect 6327 6628 6361 6662
rect 6417 6628 6451 6662
rect 6507 6628 6541 6662
rect 6597 6628 6631 6662
rect 6687 6628 6721 6662
rect 6777 6628 6811 6662
rect 6237 6538 6271 6572
rect 6327 6538 6361 6572
rect 6417 6538 6451 6572
rect 6507 6538 6541 6572
rect 6597 6538 6631 6572
rect 6687 6538 6721 6572
rect 6777 6538 6811 6572
rect 6237 6448 6271 6482
rect 6327 6448 6361 6482
rect 6417 6448 6451 6482
rect 6507 6448 6541 6482
rect 6597 6448 6631 6482
rect 6687 6448 6721 6482
rect 6777 6448 6811 6482
rect 6237 6358 6271 6392
rect 6327 6358 6361 6392
rect 6417 6358 6451 6392
rect 6507 6358 6541 6392
rect 6597 6358 6631 6392
rect 6687 6358 6721 6392
rect 6777 6358 6811 6392
rect 6237 6268 6271 6302
rect 6327 6268 6361 6302
rect 6417 6268 6451 6302
rect 6507 6268 6541 6302
rect 6597 6268 6631 6302
rect 6687 6268 6721 6302
rect 6777 6268 6811 6302
rect 6237 6178 6271 6212
rect 6327 6178 6361 6212
rect 6417 6178 6451 6212
rect 6507 6178 6541 6212
rect 6597 6178 6631 6212
rect 6687 6178 6721 6212
rect 6777 6178 6811 6212
rect 6237 6088 6271 6122
rect 6327 6088 6361 6122
rect 6417 6088 6451 6122
rect 6507 6088 6541 6122
rect 6597 6088 6631 6122
rect 6687 6088 6721 6122
rect 6777 6088 6811 6122
rect 685 5240 719 5274
rect 775 5240 809 5274
rect 865 5240 899 5274
rect 955 5240 989 5274
rect 1045 5240 1079 5274
rect 1135 5240 1169 5274
rect 1225 5240 1259 5274
rect 685 5150 719 5184
rect 775 5150 809 5184
rect 865 5150 899 5184
rect 955 5150 989 5184
rect 1045 5150 1079 5184
rect 1135 5150 1169 5184
rect 1225 5150 1259 5184
rect 685 5060 719 5094
rect 775 5060 809 5094
rect 865 5060 899 5094
rect 955 5060 989 5094
rect 1045 5060 1079 5094
rect 1135 5060 1169 5094
rect 1225 5060 1259 5094
rect 685 4970 719 5004
rect 775 4970 809 5004
rect 865 4970 899 5004
rect 955 4970 989 5004
rect 1045 4970 1079 5004
rect 1135 4970 1169 5004
rect 1225 4970 1259 5004
rect 685 4880 719 4914
rect 775 4880 809 4914
rect 865 4880 899 4914
rect 955 4880 989 4914
rect 1045 4880 1079 4914
rect 1135 4880 1169 4914
rect 1225 4880 1259 4914
rect 685 4790 719 4824
rect 775 4790 809 4824
rect 865 4790 899 4824
rect 955 4790 989 4824
rect 1045 4790 1079 4824
rect 1135 4790 1169 4824
rect 1225 4790 1259 4824
rect 685 4700 719 4734
rect 775 4700 809 4734
rect 865 4700 899 4734
rect 955 4700 989 4734
rect 1045 4700 1079 4734
rect 1135 4700 1169 4734
rect 1225 4700 1259 4734
rect 2073 5240 2107 5274
rect 2163 5240 2197 5274
rect 2253 5240 2287 5274
rect 2343 5240 2377 5274
rect 2433 5240 2467 5274
rect 2523 5240 2557 5274
rect 2613 5240 2647 5274
rect 2073 5150 2107 5184
rect 2163 5150 2197 5184
rect 2253 5150 2287 5184
rect 2343 5150 2377 5184
rect 2433 5150 2467 5184
rect 2523 5150 2557 5184
rect 2613 5150 2647 5184
rect 2073 5060 2107 5094
rect 2163 5060 2197 5094
rect 2253 5060 2287 5094
rect 2343 5060 2377 5094
rect 2433 5060 2467 5094
rect 2523 5060 2557 5094
rect 2613 5060 2647 5094
rect 2073 4970 2107 5004
rect 2163 4970 2197 5004
rect 2253 4970 2287 5004
rect 2343 4970 2377 5004
rect 2433 4970 2467 5004
rect 2523 4970 2557 5004
rect 2613 4970 2647 5004
rect 2073 4880 2107 4914
rect 2163 4880 2197 4914
rect 2253 4880 2287 4914
rect 2343 4880 2377 4914
rect 2433 4880 2467 4914
rect 2523 4880 2557 4914
rect 2613 4880 2647 4914
rect 2073 4790 2107 4824
rect 2163 4790 2197 4824
rect 2253 4790 2287 4824
rect 2343 4790 2377 4824
rect 2433 4790 2467 4824
rect 2523 4790 2557 4824
rect 2613 4790 2647 4824
rect 2073 4700 2107 4734
rect 2163 4700 2197 4734
rect 2253 4700 2287 4734
rect 2343 4700 2377 4734
rect 2433 4700 2467 4734
rect 2523 4700 2557 4734
rect 2613 4700 2647 4734
rect 3461 5240 3495 5274
rect 3551 5240 3585 5274
rect 3641 5240 3675 5274
rect 3731 5240 3765 5274
rect 3821 5240 3855 5274
rect 3911 5240 3945 5274
rect 4001 5240 4035 5274
rect 3461 5150 3495 5184
rect 3551 5150 3585 5184
rect 3641 5150 3675 5184
rect 3731 5150 3765 5184
rect 3821 5150 3855 5184
rect 3911 5150 3945 5184
rect 4001 5150 4035 5184
rect 3461 5060 3495 5094
rect 3551 5060 3585 5094
rect 3641 5060 3675 5094
rect 3731 5060 3765 5094
rect 3821 5060 3855 5094
rect 3911 5060 3945 5094
rect 4001 5060 4035 5094
rect 3461 4970 3495 5004
rect 3551 4970 3585 5004
rect 3641 4970 3675 5004
rect 3731 4970 3765 5004
rect 3821 4970 3855 5004
rect 3911 4970 3945 5004
rect 4001 4970 4035 5004
rect 3461 4880 3495 4914
rect 3551 4880 3585 4914
rect 3641 4880 3675 4914
rect 3731 4880 3765 4914
rect 3821 4880 3855 4914
rect 3911 4880 3945 4914
rect 4001 4880 4035 4914
rect 3461 4790 3495 4824
rect 3551 4790 3585 4824
rect 3641 4790 3675 4824
rect 3731 4790 3765 4824
rect 3821 4790 3855 4824
rect 3911 4790 3945 4824
rect 4001 4790 4035 4824
rect 3461 4700 3495 4734
rect 3551 4700 3585 4734
rect 3641 4700 3675 4734
rect 3731 4700 3765 4734
rect 3821 4700 3855 4734
rect 3911 4700 3945 4734
rect 4001 4700 4035 4734
rect 4849 5240 4883 5274
rect 4939 5240 4973 5274
rect 5029 5240 5063 5274
rect 5119 5240 5153 5274
rect 5209 5240 5243 5274
rect 5299 5240 5333 5274
rect 5389 5240 5423 5274
rect 4849 5150 4883 5184
rect 4939 5150 4973 5184
rect 5029 5150 5063 5184
rect 5119 5150 5153 5184
rect 5209 5150 5243 5184
rect 5299 5150 5333 5184
rect 5389 5150 5423 5184
rect 4849 5060 4883 5094
rect 4939 5060 4973 5094
rect 5029 5060 5063 5094
rect 5119 5060 5153 5094
rect 5209 5060 5243 5094
rect 5299 5060 5333 5094
rect 5389 5060 5423 5094
rect 4849 4970 4883 5004
rect 4939 4970 4973 5004
rect 5029 4970 5063 5004
rect 5119 4970 5153 5004
rect 5209 4970 5243 5004
rect 5299 4970 5333 5004
rect 5389 4970 5423 5004
rect 4849 4880 4883 4914
rect 4939 4880 4973 4914
rect 5029 4880 5063 4914
rect 5119 4880 5153 4914
rect 5209 4880 5243 4914
rect 5299 4880 5333 4914
rect 5389 4880 5423 4914
rect 4849 4790 4883 4824
rect 4939 4790 4973 4824
rect 5029 4790 5063 4824
rect 5119 4790 5153 4824
rect 5209 4790 5243 4824
rect 5299 4790 5333 4824
rect 5389 4790 5423 4824
rect 4849 4700 4883 4734
rect 4939 4700 4973 4734
rect 5029 4700 5063 4734
rect 5119 4700 5153 4734
rect 5209 4700 5243 4734
rect 5299 4700 5333 4734
rect 5389 4700 5423 4734
rect 6237 5240 6271 5274
rect 6327 5240 6361 5274
rect 6417 5240 6451 5274
rect 6507 5240 6541 5274
rect 6597 5240 6631 5274
rect 6687 5240 6721 5274
rect 6777 5240 6811 5274
rect 6237 5150 6271 5184
rect 6327 5150 6361 5184
rect 6417 5150 6451 5184
rect 6507 5150 6541 5184
rect 6597 5150 6631 5184
rect 6687 5150 6721 5184
rect 6777 5150 6811 5184
rect 6237 5060 6271 5094
rect 6327 5060 6361 5094
rect 6417 5060 6451 5094
rect 6507 5060 6541 5094
rect 6597 5060 6631 5094
rect 6687 5060 6721 5094
rect 6777 5060 6811 5094
rect 6237 4970 6271 5004
rect 6327 4970 6361 5004
rect 6417 4970 6451 5004
rect 6507 4970 6541 5004
rect 6597 4970 6631 5004
rect 6687 4970 6721 5004
rect 6777 4970 6811 5004
rect 6237 4880 6271 4914
rect 6327 4880 6361 4914
rect 6417 4880 6451 4914
rect 6507 4880 6541 4914
rect 6597 4880 6631 4914
rect 6687 4880 6721 4914
rect 6777 4880 6811 4914
rect 6237 4790 6271 4824
rect 6327 4790 6361 4824
rect 6417 4790 6451 4824
rect 6507 4790 6541 4824
rect 6597 4790 6631 4824
rect 6687 4790 6721 4824
rect 6777 4790 6811 4824
rect 6237 4700 6271 4734
rect 6327 4700 6361 4734
rect 6417 4700 6451 4734
rect 6507 4700 6541 4734
rect 6597 4700 6631 4734
rect 6687 4700 6721 4734
rect 6777 4700 6811 4734
rect 685 3852 719 3886
rect 775 3852 809 3886
rect 865 3852 899 3886
rect 955 3852 989 3886
rect 1045 3852 1079 3886
rect 1135 3852 1169 3886
rect 1225 3852 1259 3886
rect 685 3762 719 3796
rect 775 3762 809 3796
rect 865 3762 899 3796
rect 955 3762 989 3796
rect 1045 3762 1079 3796
rect 1135 3762 1169 3796
rect 1225 3762 1259 3796
rect 685 3672 719 3706
rect 775 3672 809 3706
rect 865 3672 899 3706
rect 955 3672 989 3706
rect 1045 3672 1079 3706
rect 1135 3672 1169 3706
rect 1225 3672 1259 3706
rect 685 3582 719 3616
rect 775 3582 809 3616
rect 865 3582 899 3616
rect 955 3582 989 3616
rect 1045 3582 1079 3616
rect 1135 3582 1169 3616
rect 1225 3582 1259 3616
rect 685 3492 719 3526
rect 775 3492 809 3526
rect 865 3492 899 3526
rect 955 3492 989 3526
rect 1045 3492 1079 3526
rect 1135 3492 1169 3526
rect 1225 3492 1259 3526
rect 685 3402 719 3436
rect 775 3402 809 3436
rect 865 3402 899 3436
rect 955 3402 989 3436
rect 1045 3402 1079 3436
rect 1135 3402 1169 3436
rect 1225 3402 1259 3436
rect 685 3312 719 3346
rect 775 3312 809 3346
rect 865 3312 899 3346
rect 955 3312 989 3346
rect 1045 3312 1079 3346
rect 1135 3312 1169 3346
rect 1225 3312 1259 3346
rect 2073 3852 2107 3886
rect 2163 3852 2197 3886
rect 2253 3852 2287 3886
rect 2343 3852 2377 3886
rect 2433 3852 2467 3886
rect 2523 3852 2557 3886
rect 2613 3852 2647 3886
rect 2073 3762 2107 3796
rect 2163 3762 2197 3796
rect 2253 3762 2287 3796
rect 2343 3762 2377 3796
rect 2433 3762 2467 3796
rect 2523 3762 2557 3796
rect 2613 3762 2647 3796
rect 2073 3672 2107 3706
rect 2163 3672 2197 3706
rect 2253 3672 2287 3706
rect 2343 3672 2377 3706
rect 2433 3672 2467 3706
rect 2523 3672 2557 3706
rect 2613 3672 2647 3706
rect 2073 3582 2107 3616
rect 2163 3582 2197 3616
rect 2253 3582 2287 3616
rect 2343 3582 2377 3616
rect 2433 3582 2467 3616
rect 2523 3582 2557 3616
rect 2613 3582 2647 3616
rect 2073 3492 2107 3526
rect 2163 3492 2197 3526
rect 2253 3492 2287 3526
rect 2343 3492 2377 3526
rect 2433 3492 2467 3526
rect 2523 3492 2557 3526
rect 2613 3492 2647 3526
rect 2073 3402 2107 3436
rect 2163 3402 2197 3436
rect 2253 3402 2287 3436
rect 2343 3402 2377 3436
rect 2433 3402 2467 3436
rect 2523 3402 2557 3436
rect 2613 3402 2647 3436
rect 2073 3312 2107 3346
rect 2163 3312 2197 3346
rect 2253 3312 2287 3346
rect 2343 3312 2377 3346
rect 2433 3312 2467 3346
rect 2523 3312 2557 3346
rect 2613 3312 2647 3346
rect 3461 3852 3495 3886
rect 3551 3852 3585 3886
rect 3641 3852 3675 3886
rect 3731 3852 3765 3886
rect 3821 3852 3855 3886
rect 3911 3852 3945 3886
rect 4001 3852 4035 3886
rect 3461 3762 3495 3796
rect 3551 3762 3585 3796
rect 3641 3762 3675 3796
rect 3731 3762 3765 3796
rect 3821 3762 3855 3796
rect 3911 3762 3945 3796
rect 4001 3762 4035 3796
rect 3461 3672 3495 3706
rect 3551 3672 3585 3706
rect 3641 3672 3675 3706
rect 3731 3672 3765 3706
rect 3821 3672 3855 3706
rect 3911 3672 3945 3706
rect 4001 3672 4035 3706
rect 3461 3582 3495 3616
rect 3551 3582 3585 3616
rect 3641 3582 3675 3616
rect 3731 3582 3765 3616
rect 3821 3582 3855 3616
rect 3911 3582 3945 3616
rect 4001 3582 4035 3616
rect 3461 3492 3495 3526
rect 3551 3492 3585 3526
rect 3641 3492 3675 3526
rect 3731 3492 3765 3526
rect 3821 3492 3855 3526
rect 3911 3492 3945 3526
rect 4001 3492 4035 3526
rect 3461 3402 3495 3436
rect 3551 3402 3585 3436
rect 3641 3402 3675 3436
rect 3731 3402 3765 3436
rect 3821 3402 3855 3436
rect 3911 3402 3945 3436
rect 4001 3402 4035 3436
rect 3461 3312 3495 3346
rect 3551 3312 3585 3346
rect 3641 3312 3675 3346
rect 3731 3312 3765 3346
rect 3821 3312 3855 3346
rect 3911 3312 3945 3346
rect 4001 3312 4035 3346
rect 4849 3852 4883 3886
rect 4939 3852 4973 3886
rect 5029 3852 5063 3886
rect 5119 3852 5153 3886
rect 5209 3852 5243 3886
rect 5299 3852 5333 3886
rect 5389 3852 5423 3886
rect 4849 3762 4883 3796
rect 4939 3762 4973 3796
rect 5029 3762 5063 3796
rect 5119 3762 5153 3796
rect 5209 3762 5243 3796
rect 5299 3762 5333 3796
rect 5389 3762 5423 3796
rect 4849 3672 4883 3706
rect 4939 3672 4973 3706
rect 5029 3672 5063 3706
rect 5119 3672 5153 3706
rect 5209 3672 5243 3706
rect 5299 3672 5333 3706
rect 5389 3672 5423 3706
rect 4849 3582 4883 3616
rect 4939 3582 4973 3616
rect 5029 3582 5063 3616
rect 5119 3582 5153 3616
rect 5209 3582 5243 3616
rect 5299 3582 5333 3616
rect 5389 3582 5423 3616
rect 4849 3492 4883 3526
rect 4939 3492 4973 3526
rect 5029 3492 5063 3526
rect 5119 3492 5153 3526
rect 5209 3492 5243 3526
rect 5299 3492 5333 3526
rect 5389 3492 5423 3526
rect 4849 3402 4883 3436
rect 4939 3402 4973 3436
rect 5029 3402 5063 3436
rect 5119 3402 5153 3436
rect 5209 3402 5243 3436
rect 5299 3402 5333 3436
rect 5389 3402 5423 3436
rect 4849 3312 4883 3346
rect 4939 3312 4973 3346
rect 5029 3312 5063 3346
rect 5119 3312 5153 3346
rect 5209 3312 5243 3346
rect 5299 3312 5333 3346
rect 5389 3312 5423 3346
rect 6237 3852 6271 3886
rect 6327 3852 6361 3886
rect 6417 3852 6451 3886
rect 6507 3852 6541 3886
rect 6597 3852 6631 3886
rect 6687 3852 6721 3886
rect 6777 3852 6811 3886
rect 6237 3762 6271 3796
rect 6327 3762 6361 3796
rect 6417 3762 6451 3796
rect 6507 3762 6541 3796
rect 6597 3762 6631 3796
rect 6687 3762 6721 3796
rect 6777 3762 6811 3796
rect 6237 3672 6271 3706
rect 6327 3672 6361 3706
rect 6417 3672 6451 3706
rect 6507 3672 6541 3706
rect 6597 3672 6631 3706
rect 6687 3672 6721 3706
rect 6777 3672 6811 3706
rect 6237 3582 6271 3616
rect 6327 3582 6361 3616
rect 6417 3582 6451 3616
rect 6507 3582 6541 3616
rect 6597 3582 6631 3616
rect 6687 3582 6721 3616
rect 6777 3582 6811 3616
rect 6237 3492 6271 3526
rect 6327 3492 6361 3526
rect 6417 3492 6451 3526
rect 6507 3492 6541 3526
rect 6597 3492 6631 3526
rect 6687 3492 6721 3526
rect 6777 3492 6811 3526
rect 6237 3402 6271 3436
rect 6327 3402 6361 3436
rect 6417 3402 6451 3436
rect 6507 3402 6541 3436
rect 6597 3402 6631 3436
rect 6687 3402 6721 3436
rect 6777 3402 6811 3436
rect 6237 3312 6271 3346
rect 6327 3312 6361 3346
rect 6417 3312 6451 3346
rect 6507 3312 6541 3346
rect 6597 3312 6631 3346
rect 6687 3312 6721 3346
rect 6777 3312 6811 3346
rect 685 2464 719 2498
rect 775 2464 809 2498
rect 865 2464 899 2498
rect 955 2464 989 2498
rect 1045 2464 1079 2498
rect 1135 2464 1169 2498
rect 1225 2464 1259 2498
rect 685 2374 719 2408
rect 775 2374 809 2408
rect 865 2374 899 2408
rect 955 2374 989 2408
rect 1045 2374 1079 2408
rect 1135 2374 1169 2408
rect 1225 2374 1259 2408
rect 685 2284 719 2318
rect 775 2284 809 2318
rect 865 2284 899 2318
rect 955 2284 989 2318
rect 1045 2284 1079 2318
rect 1135 2284 1169 2318
rect 1225 2284 1259 2318
rect 685 2194 719 2228
rect 775 2194 809 2228
rect 865 2194 899 2228
rect 955 2194 989 2228
rect 1045 2194 1079 2228
rect 1135 2194 1169 2228
rect 1225 2194 1259 2228
rect 685 2104 719 2138
rect 775 2104 809 2138
rect 865 2104 899 2138
rect 955 2104 989 2138
rect 1045 2104 1079 2138
rect 1135 2104 1169 2138
rect 1225 2104 1259 2138
rect 685 2014 719 2048
rect 775 2014 809 2048
rect 865 2014 899 2048
rect 955 2014 989 2048
rect 1045 2014 1079 2048
rect 1135 2014 1169 2048
rect 1225 2014 1259 2048
rect 685 1924 719 1958
rect 775 1924 809 1958
rect 865 1924 899 1958
rect 955 1924 989 1958
rect 1045 1924 1079 1958
rect 1135 1924 1169 1958
rect 1225 1924 1259 1958
rect 2073 2464 2107 2498
rect 2163 2464 2197 2498
rect 2253 2464 2287 2498
rect 2343 2464 2377 2498
rect 2433 2464 2467 2498
rect 2523 2464 2557 2498
rect 2613 2464 2647 2498
rect 2073 2374 2107 2408
rect 2163 2374 2197 2408
rect 2253 2374 2287 2408
rect 2343 2374 2377 2408
rect 2433 2374 2467 2408
rect 2523 2374 2557 2408
rect 2613 2374 2647 2408
rect 2073 2284 2107 2318
rect 2163 2284 2197 2318
rect 2253 2284 2287 2318
rect 2343 2284 2377 2318
rect 2433 2284 2467 2318
rect 2523 2284 2557 2318
rect 2613 2284 2647 2318
rect 2073 2194 2107 2228
rect 2163 2194 2197 2228
rect 2253 2194 2287 2228
rect 2343 2194 2377 2228
rect 2433 2194 2467 2228
rect 2523 2194 2557 2228
rect 2613 2194 2647 2228
rect 2073 2104 2107 2138
rect 2163 2104 2197 2138
rect 2253 2104 2287 2138
rect 2343 2104 2377 2138
rect 2433 2104 2467 2138
rect 2523 2104 2557 2138
rect 2613 2104 2647 2138
rect 2073 2014 2107 2048
rect 2163 2014 2197 2048
rect 2253 2014 2287 2048
rect 2343 2014 2377 2048
rect 2433 2014 2467 2048
rect 2523 2014 2557 2048
rect 2613 2014 2647 2048
rect 2073 1924 2107 1958
rect 2163 1924 2197 1958
rect 2253 1924 2287 1958
rect 2343 1924 2377 1958
rect 2433 1924 2467 1958
rect 2523 1924 2557 1958
rect 2613 1924 2647 1958
rect 3461 2464 3495 2498
rect 3551 2464 3585 2498
rect 3641 2464 3675 2498
rect 3731 2464 3765 2498
rect 3821 2464 3855 2498
rect 3911 2464 3945 2498
rect 4001 2464 4035 2498
rect 3461 2374 3495 2408
rect 3551 2374 3585 2408
rect 3641 2374 3675 2408
rect 3731 2374 3765 2408
rect 3821 2374 3855 2408
rect 3911 2374 3945 2408
rect 4001 2374 4035 2408
rect 3461 2284 3495 2318
rect 3551 2284 3585 2318
rect 3641 2284 3675 2318
rect 3731 2284 3765 2318
rect 3821 2284 3855 2318
rect 3911 2284 3945 2318
rect 4001 2284 4035 2318
rect 3461 2194 3495 2228
rect 3551 2194 3585 2228
rect 3641 2194 3675 2228
rect 3731 2194 3765 2228
rect 3821 2194 3855 2228
rect 3911 2194 3945 2228
rect 4001 2194 4035 2228
rect 3461 2104 3495 2138
rect 3551 2104 3585 2138
rect 3641 2104 3675 2138
rect 3731 2104 3765 2138
rect 3821 2104 3855 2138
rect 3911 2104 3945 2138
rect 4001 2104 4035 2138
rect 3461 2014 3495 2048
rect 3551 2014 3585 2048
rect 3641 2014 3675 2048
rect 3731 2014 3765 2048
rect 3821 2014 3855 2048
rect 3911 2014 3945 2048
rect 4001 2014 4035 2048
rect 3461 1924 3495 1958
rect 3551 1924 3585 1958
rect 3641 1924 3675 1958
rect 3731 1924 3765 1958
rect 3821 1924 3855 1958
rect 3911 1924 3945 1958
rect 4001 1924 4035 1958
rect 4849 2464 4883 2498
rect 4939 2464 4973 2498
rect 5029 2464 5063 2498
rect 5119 2464 5153 2498
rect 5209 2464 5243 2498
rect 5299 2464 5333 2498
rect 5389 2464 5423 2498
rect 4849 2374 4883 2408
rect 4939 2374 4973 2408
rect 5029 2374 5063 2408
rect 5119 2374 5153 2408
rect 5209 2374 5243 2408
rect 5299 2374 5333 2408
rect 5389 2374 5423 2408
rect 4849 2284 4883 2318
rect 4939 2284 4973 2318
rect 5029 2284 5063 2318
rect 5119 2284 5153 2318
rect 5209 2284 5243 2318
rect 5299 2284 5333 2318
rect 5389 2284 5423 2318
rect 4849 2194 4883 2228
rect 4939 2194 4973 2228
rect 5029 2194 5063 2228
rect 5119 2194 5153 2228
rect 5209 2194 5243 2228
rect 5299 2194 5333 2228
rect 5389 2194 5423 2228
rect 4849 2104 4883 2138
rect 4939 2104 4973 2138
rect 5029 2104 5063 2138
rect 5119 2104 5153 2138
rect 5209 2104 5243 2138
rect 5299 2104 5333 2138
rect 5389 2104 5423 2138
rect 4849 2014 4883 2048
rect 4939 2014 4973 2048
rect 5029 2014 5063 2048
rect 5119 2014 5153 2048
rect 5209 2014 5243 2048
rect 5299 2014 5333 2048
rect 5389 2014 5423 2048
rect 4849 1924 4883 1958
rect 4939 1924 4973 1958
rect 5029 1924 5063 1958
rect 5119 1924 5153 1958
rect 5209 1924 5243 1958
rect 5299 1924 5333 1958
rect 5389 1924 5423 1958
rect 6237 2464 6271 2498
rect 6327 2464 6361 2498
rect 6417 2464 6451 2498
rect 6507 2464 6541 2498
rect 6597 2464 6631 2498
rect 6687 2464 6721 2498
rect 6777 2464 6811 2498
rect 6237 2374 6271 2408
rect 6327 2374 6361 2408
rect 6417 2374 6451 2408
rect 6507 2374 6541 2408
rect 6597 2374 6631 2408
rect 6687 2374 6721 2408
rect 6777 2374 6811 2408
rect 6237 2284 6271 2318
rect 6327 2284 6361 2318
rect 6417 2284 6451 2318
rect 6507 2284 6541 2318
rect 6597 2284 6631 2318
rect 6687 2284 6721 2318
rect 6777 2284 6811 2318
rect 6237 2194 6271 2228
rect 6327 2194 6361 2228
rect 6417 2194 6451 2228
rect 6507 2194 6541 2228
rect 6597 2194 6631 2228
rect 6687 2194 6721 2228
rect 6777 2194 6811 2228
rect 6237 2104 6271 2138
rect 6327 2104 6361 2138
rect 6417 2104 6451 2138
rect 6507 2104 6541 2138
rect 6597 2104 6631 2138
rect 6687 2104 6721 2138
rect 6777 2104 6811 2138
rect 6237 2014 6271 2048
rect 6327 2014 6361 2048
rect 6417 2014 6451 2048
rect 6507 2014 6541 2048
rect 6597 2014 6631 2048
rect 6687 2014 6721 2048
rect 6777 2014 6811 2048
rect 6237 1924 6271 1958
rect 6327 1924 6361 1958
rect 6417 1924 6451 1958
rect 6507 1924 6541 1958
rect 6597 1924 6631 1958
rect 6687 1924 6721 1958
rect 6777 1924 6811 1958
<< psubdiff >>
rect -17500 22657 -17440 22691
rect 8642 22657 8702 22691
rect -17500 22631 -17466 22657
rect 8668 22631 8702 22657
rect -17500 20886 -17466 20912
rect 8668 20886 8702 20912
rect -17500 20852 -17440 20886
rect 8642 20852 8702 20886
rect -13149 20761 -13053 20795
rect 8591 20761 8687 20795
rect -13149 20699 -13115 20761
rect 8653 20699 8687 20761
rect -13149 19337 -13115 19399
rect 8653 19337 8687 19399
rect -13149 19303 -13053 19337
rect 8591 19303 8687 19337
rect -7165 19197 -7069 19231
rect 8591 19197 8687 19231
rect -7165 19135 -7131 19197
rect 8653 19135 8687 19197
rect -7165 17773 -7131 17835
rect 8653 17773 8687 17835
rect -7165 17739 -7069 17773
rect 8591 17739 8687 17773
rect -1270 17574 -1210 17608
rect -404 17574 -344 17608
rect -1270 17541 -1236 17574
rect -378 17541 -344 17574
rect -1270 16820 -1236 16854
rect -378 16820 -344 16843
rect -1270 16786 -1210 16820
rect -404 16786 -344 16820
rect -209 17587 -149 17621
rect 8627 17587 8687 17621
rect -209 17539 -175 17587
rect 8653 17539 8687 17587
rect -209 15959 -175 15985
rect 8653 15959 8687 15985
rect -209 15925 -149 15959
rect 8627 15925 8687 15959
rect -1220 15829 -1160 15863
rect 2568 15829 2628 15863
rect -1220 15803 -1186 15829
rect 2594 15803 2628 15829
rect -1220 14737 -1186 14763
rect 2865 15744 2927 15778
rect 8625 15744 8687 15778
rect 2865 15703 2899 15744
rect 8653 15703 8687 15744
rect 2865 14820 2899 14861
rect 8653 14820 8687 14861
rect 2865 14786 2927 14820
rect 8625 14786 8687 14820
rect 2594 14737 2628 14763
rect -1220 14703 -1160 14737
rect 2568 14703 2628 14737
rect 604 12297 664 12331
rect 1470 12297 1556 12331
rect 2362 12297 2448 12331
rect 3254 12297 3340 12331
rect 4146 12297 4206 12331
rect 604 12271 638 12297
rect 1496 12271 1530 12297
rect 604 10265 638 10291
rect 2388 12271 2422 12297
rect 1496 10265 1530 10291
rect 3280 12271 3314 12297
rect 2388 10265 2422 10291
rect 4172 12271 4206 12297
rect 3280 10265 3314 10291
rect 4260 12267 4320 12301
rect 4712 12267 4772 12301
rect 4260 12241 4294 12267
rect 4738 12241 4772 12267
rect 4260 11409 4294 11435
rect 4738 11409 4772 11435
rect 4260 11375 4320 11409
rect 4712 11375 4772 11409
rect 4172 10265 4206 10291
rect 604 10231 664 10265
rect 1470 10231 1556 10265
rect 2362 10231 2448 10265
rect 3254 10231 3340 10265
rect 4146 10231 4206 10265
rect 4260 11153 4320 11187
rect 4712 11153 4772 11187
rect 4260 11127 4294 11153
rect 4738 11127 4772 11153
rect 4260 10295 4294 10321
rect 4738 10295 4772 10321
rect 4260 10261 4320 10295
rect 4712 10261 4772 10295
rect 329 8373 1617 8406
rect 329 8339 387 8373
rect 421 8339 477 8373
rect 511 8339 567 8373
rect 601 8339 657 8373
rect 691 8339 747 8373
rect 781 8339 837 8373
rect 871 8339 927 8373
rect 961 8339 1017 8373
rect 1051 8339 1107 8373
rect 1141 8339 1197 8373
rect 1231 8339 1287 8373
rect 1321 8339 1377 8373
rect 1411 8339 1467 8373
rect 1501 8339 1617 8373
rect 329 8305 1617 8339
rect 329 8272 430 8305
rect 329 8238 364 8272
rect 398 8238 430 8272
rect 1516 8272 1617 8305
rect 329 8182 430 8238
rect 329 8148 364 8182
rect 398 8148 430 8182
rect 329 8092 430 8148
rect 329 8058 364 8092
rect 398 8058 430 8092
rect 329 8002 430 8058
rect 329 7968 364 8002
rect 398 7968 430 8002
rect 329 7912 430 7968
rect 329 7878 364 7912
rect 398 7878 430 7912
rect 329 7822 430 7878
rect 329 7788 364 7822
rect 398 7788 430 7822
rect 329 7732 430 7788
rect 329 7698 364 7732
rect 398 7698 430 7732
rect 329 7642 430 7698
rect 329 7608 364 7642
rect 398 7608 430 7642
rect 329 7552 430 7608
rect 329 7518 364 7552
rect 398 7518 430 7552
rect 329 7462 430 7518
rect 329 7428 364 7462
rect 398 7428 430 7462
rect 329 7372 430 7428
rect 329 7338 364 7372
rect 398 7338 430 7372
rect 329 7282 430 7338
rect 329 7248 364 7282
rect 398 7248 430 7282
rect 1516 8238 1551 8272
rect 1585 8238 1617 8272
rect 1516 8182 1617 8238
rect 1516 8148 1551 8182
rect 1585 8148 1617 8182
rect 1516 8092 1617 8148
rect 1516 8058 1551 8092
rect 1585 8058 1617 8092
rect 1516 8002 1617 8058
rect 1516 7968 1551 8002
rect 1585 7968 1617 8002
rect 1516 7912 1617 7968
rect 1516 7878 1551 7912
rect 1585 7878 1617 7912
rect 1516 7822 1617 7878
rect 1516 7788 1551 7822
rect 1585 7788 1617 7822
rect 1516 7732 1617 7788
rect 1516 7698 1551 7732
rect 1585 7698 1617 7732
rect 1516 7642 1617 7698
rect 1516 7608 1551 7642
rect 1585 7608 1617 7642
rect 1516 7552 1617 7608
rect 1516 7518 1551 7552
rect 1585 7518 1617 7552
rect 1516 7462 1617 7518
rect 1516 7428 1551 7462
rect 1585 7428 1617 7462
rect 1516 7372 1617 7428
rect 1516 7338 1551 7372
rect 1585 7338 1617 7372
rect 1516 7282 1617 7338
rect 329 7219 430 7248
rect 1516 7248 1551 7282
rect 1585 7248 1617 7282
rect 1516 7219 1617 7248
rect 329 7186 1617 7219
rect 329 7152 387 7186
rect 421 7152 477 7186
rect 511 7152 567 7186
rect 601 7152 657 7186
rect 691 7152 747 7186
rect 781 7152 837 7186
rect 871 7152 927 7186
rect 961 7152 1017 7186
rect 1051 7152 1107 7186
rect 1141 7152 1197 7186
rect 1231 7152 1287 7186
rect 1321 7152 1377 7186
rect 1411 7152 1467 7186
rect 1501 7152 1617 7186
rect 329 7118 1617 7152
rect 1717 8373 3005 8406
rect 1717 8339 1775 8373
rect 1809 8339 1865 8373
rect 1899 8339 1955 8373
rect 1989 8339 2045 8373
rect 2079 8339 2135 8373
rect 2169 8339 2225 8373
rect 2259 8339 2315 8373
rect 2349 8339 2405 8373
rect 2439 8339 2495 8373
rect 2529 8339 2585 8373
rect 2619 8339 2675 8373
rect 2709 8339 2765 8373
rect 2799 8339 2855 8373
rect 2889 8339 3005 8373
rect 1717 8305 3005 8339
rect 1717 8272 1818 8305
rect 1717 8238 1752 8272
rect 1786 8238 1818 8272
rect 2904 8272 3005 8305
rect 1717 8182 1818 8238
rect 1717 8148 1752 8182
rect 1786 8148 1818 8182
rect 1717 8092 1818 8148
rect 1717 8058 1752 8092
rect 1786 8058 1818 8092
rect 1717 8002 1818 8058
rect 1717 7968 1752 8002
rect 1786 7968 1818 8002
rect 1717 7912 1818 7968
rect 1717 7878 1752 7912
rect 1786 7878 1818 7912
rect 1717 7822 1818 7878
rect 1717 7788 1752 7822
rect 1786 7788 1818 7822
rect 1717 7732 1818 7788
rect 1717 7698 1752 7732
rect 1786 7698 1818 7732
rect 1717 7642 1818 7698
rect 1717 7608 1752 7642
rect 1786 7608 1818 7642
rect 1717 7552 1818 7608
rect 1717 7518 1752 7552
rect 1786 7518 1818 7552
rect 1717 7462 1818 7518
rect 1717 7428 1752 7462
rect 1786 7428 1818 7462
rect 1717 7372 1818 7428
rect 1717 7338 1752 7372
rect 1786 7338 1818 7372
rect 1717 7282 1818 7338
rect 1717 7248 1752 7282
rect 1786 7248 1818 7282
rect 2904 8238 2939 8272
rect 2973 8238 3005 8272
rect 2904 8182 3005 8238
rect 2904 8148 2939 8182
rect 2973 8148 3005 8182
rect 2904 8092 3005 8148
rect 2904 8058 2939 8092
rect 2973 8058 3005 8092
rect 2904 8002 3005 8058
rect 2904 7968 2939 8002
rect 2973 7968 3005 8002
rect 2904 7912 3005 7968
rect 2904 7878 2939 7912
rect 2973 7878 3005 7912
rect 2904 7822 3005 7878
rect 2904 7788 2939 7822
rect 2973 7788 3005 7822
rect 2904 7732 3005 7788
rect 2904 7698 2939 7732
rect 2973 7698 3005 7732
rect 2904 7642 3005 7698
rect 2904 7608 2939 7642
rect 2973 7608 3005 7642
rect 2904 7552 3005 7608
rect 2904 7518 2939 7552
rect 2973 7518 3005 7552
rect 2904 7462 3005 7518
rect 2904 7428 2939 7462
rect 2973 7428 3005 7462
rect 2904 7372 3005 7428
rect 2904 7338 2939 7372
rect 2973 7338 3005 7372
rect 2904 7282 3005 7338
rect 1717 7219 1818 7248
rect 2904 7248 2939 7282
rect 2973 7248 3005 7282
rect 2904 7219 3005 7248
rect 1717 7186 3005 7219
rect 1717 7152 1775 7186
rect 1809 7152 1865 7186
rect 1899 7152 1955 7186
rect 1989 7152 2045 7186
rect 2079 7152 2135 7186
rect 2169 7152 2225 7186
rect 2259 7152 2315 7186
rect 2349 7152 2405 7186
rect 2439 7152 2495 7186
rect 2529 7152 2585 7186
rect 2619 7152 2675 7186
rect 2709 7152 2765 7186
rect 2799 7152 2855 7186
rect 2889 7152 3005 7186
rect 1717 7118 3005 7152
rect 3105 8373 4393 8406
rect 3105 8339 3163 8373
rect 3197 8339 3253 8373
rect 3287 8339 3343 8373
rect 3377 8339 3433 8373
rect 3467 8339 3523 8373
rect 3557 8339 3613 8373
rect 3647 8339 3703 8373
rect 3737 8339 3793 8373
rect 3827 8339 3883 8373
rect 3917 8339 3973 8373
rect 4007 8339 4063 8373
rect 4097 8339 4153 8373
rect 4187 8339 4243 8373
rect 4277 8339 4393 8373
rect 3105 8305 4393 8339
rect 3105 8272 3206 8305
rect 3105 8238 3140 8272
rect 3174 8238 3206 8272
rect 4292 8272 4393 8305
rect 3105 8182 3206 8238
rect 3105 8148 3140 8182
rect 3174 8148 3206 8182
rect 3105 8092 3206 8148
rect 3105 8058 3140 8092
rect 3174 8058 3206 8092
rect 3105 8002 3206 8058
rect 3105 7968 3140 8002
rect 3174 7968 3206 8002
rect 3105 7912 3206 7968
rect 3105 7878 3140 7912
rect 3174 7878 3206 7912
rect 3105 7822 3206 7878
rect 3105 7788 3140 7822
rect 3174 7788 3206 7822
rect 3105 7732 3206 7788
rect 3105 7698 3140 7732
rect 3174 7698 3206 7732
rect 3105 7642 3206 7698
rect 3105 7608 3140 7642
rect 3174 7608 3206 7642
rect 3105 7552 3206 7608
rect 3105 7518 3140 7552
rect 3174 7518 3206 7552
rect 3105 7462 3206 7518
rect 3105 7428 3140 7462
rect 3174 7428 3206 7462
rect 3105 7372 3206 7428
rect 3105 7338 3140 7372
rect 3174 7338 3206 7372
rect 3105 7282 3206 7338
rect 3105 7248 3140 7282
rect 3174 7248 3206 7282
rect 4292 8238 4327 8272
rect 4361 8238 4393 8272
rect 4292 8182 4393 8238
rect 4292 8148 4327 8182
rect 4361 8148 4393 8182
rect 4292 8092 4393 8148
rect 4292 8058 4327 8092
rect 4361 8058 4393 8092
rect 4292 8002 4393 8058
rect 4292 7968 4327 8002
rect 4361 7968 4393 8002
rect 4292 7912 4393 7968
rect 4292 7878 4327 7912
rect 4361 7878 4393 7912
rect 4292 7822 4393 7878
rect 4292 7788 4327 7822
rect 4361 7788 4393 7822
rect 4292 7732 4393 7788
rect 4292 7698 4327 7732
rect 4361 7698 4393 7732
rect 4292 7642 4393 7698
rect 4292 7608 4327 7642
rect 4361 7608 4393 7642
rect 4292 7552 4393 7608
rect 4292 7518 4327 7552
rect 4361 7518 4393 7552
rect 4292 7462 4393 7518
rect 4292 7428 4327 7462
rect 4361 7428 4393 7462
rect 4292 7372 4393 7428
rect 4292 7338 4327 7372
rect 4361 7338 4393 7372
rect 4292 7282 4393 7338
rect 3105 7219 3206 7248
rect 4292 7248 4327 7282
rect 4361 7248 4393 7282
rect 4292 7219 4393 7248
rect 3105 7186 4393 7219
rect 3105 7152 3163 7186
rect 3197 7152 3253 7186
rect 3287 7152 3343 7186
rect 3377 7152 3433 7186
rect 3467 7152 3523 7186
rect 3557 7152 3613 7186
rect 3647 7152 3703 7186
rect 3737 7152 3793 7186
rect 3827 7152 3883 7186
rect 3917 7152 3973 7186
rect 4007 7152 4063 7186
rect 4097 7152 4153 7186
rect 4187 7152 4243 7186
rect 4277 7152 4393 7186
rect 3105 7118 4393 7152
rect 4493 8373 5781 8406
rect 4493 8339 4551 8373
rect 4585 8339 4641 8373
rect 4675 8339 4731 8373
rect 4765 8339 4821 8373
rect 4855 8339 4911 8373
rect 4945 8339 5001 8373
rect 5035 8339 5091 8373
rect 5125 8339 5181 8373
rect 5215 8339 5271 8373
rect 5305 8339 5361 8373
rect 5395 8339 5451 8373
rect 5485 8339 5541 8373
rect 5575 8339 5631 8373
rect 5665 8339 5781 8373
rect 4493 8305 5781 8339
rect 4493 8272 4594 8305
rect 4493 8238 4528 8272
rect 4562 8238 4594 8272
rect 5680 8272 5781 8305
rect 4493 8182 4594 8238
rect 4493 8148 4528 8182
rect 4562 8148 4594 8182
rect 4493 8092 4594 8148
rect 4493 8058 4528 8092
rect 4562 8058 4594 8092
rect 4493 8002 4594 8058
rect 4493 7968 4528 8002
rect 4562 7968 4594 8002
rect 4493 7912 4594 7968
rect 4493 7878 4528 7912
rect 4562 7878 4594 7912
rect 4493 7822 4594 7878
rect 4493 7788 4528 7822
rect 4562 7788 4594 7822
rect 4493 7732 4594 7788
rect 4493 7698 4528 7732
rect 4562 7698 4594 7732
rect 4493 7642 4594 7698
rect 4493 7608 4528 7642
rect 4562 7608 4594 7642
rect 4493 7552 4594 7608
rect 4493 7518 4528 7552
rect 4562 7518 4594 7552
rect 4493 7462 4594 7518
rect 4493 7428 4528 7462
rect 4562 7428 4594 7462
rect 4493 7372 4594 7428
rect 4493 7338 4528 7372
rect 4562 7338 4594 7372
rect 4493 7282 4594 7338
rect 4493 7248 4528 7282
rect 4562 7248 4594 7282
rect 5680 8238 5715 8272
rect 5749 8238 5781 8272
rect 5680 8182 5781 8238
rect 5680 8148 5715 8182
rect 5749 8148 5781 8182
rect 5680 8092 5781 8148
rect 5680 8058 5715 8092
rect 5749 8058 5781 8092
rect 5680 8002 5781 8058
rect 5680 7968 5715 8002
rect 5749 7968 5781 8002
rect 5680 7912 5781 7968
rect 5680 7878 5715 7912
rect 5749 7878 5781 7912
rect 5680 7822 5781 7878
rect 5680 7788 5715 7822
rect 5749 7788 5781 7822
rect 5680 7732 5781 7788
rect 5680 7698 5715 7732
rect 5749 7698 5781 7732
rect 5680 7642 5781 7698
rect 5680 7608 5715 7642
rect 5749 7608 5781 7642
rect 5680 7552 5781 7608
rect 5680 7518 5715 7552
rect 5749 7518 5781 7552
rect 5680 7462 5781 7518
rect 5680 7428 5715 7462
rect 5749 7428 5781 7462
rect 5680 7372 5781 7428
rect 5680 7338 5715 7372
rect 5749 7338 5781 7372
rect 5680 7282 5781 7338
rect 4493 7219 4594 7248
rect 5680 7248 5715 7282
rect 5749 7248 5781 7282
rect 5680 7219 5781 7248
rect 4493 7186 5781 7219
rect 4493 7152 4551 7186
rect 4585 7152 4641 7186
rect 4675 7152 4731 7186
rect 4765 7152 4821 7186
rect 4855 7152 4911 7186
rect 4945 7152 5001 7186
rect 5035 7152 5091 7186
rect 5125 7152 5181 7186
rect 5215 7152 5271 7186
rect 5305 7152 5361 7186
rect 5395 7152 5451 7186
rect 5485 7152 5541 7186
rect 5575 7152 5631 7186
rect 5665 7152 5781 7186
rect 4493 7118 5781 7152
rect 5881 8373 7169 8406
rect 5881 8339 5939 8373
rect 5973 8339 6029 8373
rect 6063 8339 6119 8373
rect 6153 8339 6209 8373
rect 6243 8339 6299 8373
rect 6333 8339 6389 8373
rect 6423 8339 6479 8373
rect 6513 8339 6569 8373
rect 6603 8339 6659 8373
rect 6693 8339 6749 8373
rect 6783 8339 6839 8373
rect 6873 8339 6929 8373
rect 6963 8339 7019 8373
rect 7053 8339 7169 8373
rect 5881 8305 7169 8339
rect 5881 8272 5982 8305
rect 5881 8238 5916 8272
rect 5950 8238 5982 8272
rect 7068 8272 7169 8305
rect 5881 8182 5982 8238
rect 5881 8148 5916 8182
rect 5950 8148 5982 8182
rect 5881 8092 5982 8148
rect 5881 8058 5916 8092
rect 5950 8058 5982 8092
rect 5881 8002 5982 8058
rect 5881 7968 5916 8002
rect 5950 7968 5982 8002
rect 5881 7912 5982 7968
rect 5881 7878 5916 7912
rect 5950 7878 5982 7912
rect 5881 7822 5982 7878
rect 5881 7788 5916 7822
rect 5950 7788 5982 7822
rect 5881 7732 5982 7788
rect 5881 7698 5916 7732
rect 5950 7698 5982 7732
rect 5881 7642 5982 7698
rect 5881 7608 5916 7642
rect 5950 7608 5982 7642
rect 5881 7552 5982 7608
rect 5881 7518 5916 7552
rect 5950 7518 5982 7552
rect 5881 7462 5982 7518
rect 5881 7428 5916 7462
rect 5950 7428 5982 7462
rect 5881 7372 5982 7428
rect 5881 7338 5916 7372
rect 5950 7338 5982 7372
rect 5881 7282 5982 7338
rect 5881 7248 5916 7282
rect 5950 7248 5982 7282
rect 7068 8238 7103 8272
rect 7137 8238 7169 8272
rect 7068 8182 7169 8238
rect 7068 8148 7103 8182
rect 7137 8148 7169 8182
rect 7068 8092 7169 8148
rect 7068 8058 7103 8092
rect 7137 8058 7169 8092
rect 7068 8002 7169 8058
rect 7068 7968 7103 8002
rect 7137 7968 7169 8002
rect 7068 7912 7169 7968
rect 7068 7878 7103 7912
rect 7137 7878 7169 7912
rect 7068 7822 7169 7878
rect 7068 7788 7103 7822
rect 7137 7788 7169 7822
rect 7068 7732 7169 7788
rect 7068 7698 7103 7732
rect 7137 7698 7169 7732
rect 7068 7642 7169 7698
rect 7068 7608 7103 7642
rect 7137 7608 7169 7642
rect 7068 7552 7169 7608
rect 7068 7518 7103 7552
rect 7137 7518 7169 7552
rect 7068 7462 7169 7518
rect 7068 7428 7103 7462
rect 7137 7428 7169 7462
rect 7068 7372 7169 7428
rect 7068 7338 7103 7372
rect 7137 7338 7169 7372
rect 7068 7282 7169 7338
rect 5881 7219 5982 7248
rect 7068 7248 7103 7282
rect 7137 7248 7169 7282
rect 7068 7219 7169 7248
rect 5881 7186 7169 7219
rect 5881 7152 5939 7186
rect 5973 7152 6029 7186
rect 6063 7152 6119 7186
rect 6153 7152 6209 7186
rect 6243 7152 6299 7186
rect 6333 7152 6389 7186
rect 6423 7152 6479 7186
rect 6513 7152 6569 7186
rect 6603 7152 6659 7186
rect 6693 7152 6749 7186
rect 6783 7152 6839 7186
rect 6873 7152 6929 7186
rect 6963 7152 7019 7186
rect 7053 7152 7169 7186
rect 5881 7118 7169 7152
rect 329 6985 1617 7018
rect 329 6951 387 6985
rect 421 6951 477 6985
rect 511 6951 567 6985
rect 601 6951 657 6985
rect 691 6951 747 6985
rect 781 6951 837 6985
rect 871 6951 927 6985
rect 961 6951 1017 6985
rect 1051 6951 1107 6985
rect 1141 6951 1197 6985
rect 1231 6951 1287 6985
rect 1321 6951 1377 6985
rect 1411 6951 1467 6985
rect 1501 6951 1617 6985
rect 329 6917 1617 6951
rect 329 6884 430 6917
rect 329 6850 364 6884
rect 398 6850 430 6884
rect 1516 6884 1617 6917
rect 329 6794 430 6850
rect 329 6760 364 6794
rect 398 6760 430 6794
rect 329 6704 430 6760
rect 329 6670 364 6704
rect 398 6670 430 6704
rect 329 6614 430 6670
rect 329 6580 364 6614
rect 398 6580 430 6614
rect 329 6524 430 6580
rect 329 6490 364 6524
rect 398 6490 430 6524
rect 329 6434 430 6490
rect 329 6400 364 6434
rect 398 6400 430 6434
rect 329 6344 430 6400
rect 329 6310 364 6344
rect 398 6310 430 6344
rect 329 6254 430 6310
rect 329 6220 364 6254
rect 398 6220 430 6254
rect 329 6164 430 6220
rect 329 6130 364 6164
rect 398 6130 430 6164
rect 329 6074 430 6130
rect 329 6040 364 6074
rect 398 6040 430 6074
rect 329 5984 430 6040
rect 329 5950 364 5984
rect 398 5950 430 5984
rect 329 5894 430 5950
rect 329 5860 364 5894
rect 398 5860 430 5894
rect 1516 6850 1551 6884
rect 1585 6850 1617 6884
rect 1516 6794 1617 6850
rect 1516 6760 1551 6794
rect 1585 6760 1617 6794
rect 1516 6704 1617 6760
rect 1516 6670 1551 6704
rect 1585 6670 1617 6704
rect 1516 6614 1617 6670
rect 1516 6580 1551 6614
rect 1585 6580 1617 6614
rect 1516 6524 1617 6580
rect 1516 6490 1551 6524
rect 1585 6490 1617 6524
rect 1516 6434 1617 6490
rect 1516 6400 1551 6434
rect 1585 6400 1617 6434
rect 1516 6344 1617 6400
rect 1516 6310 1551 6344
rect 1585 6310 1617 6344
rect 1516 6254 1617 6310
rect 1516 6220 1551 6254
rect 1585 6220 1617 6254
rect 1516 6164 1617 6220
rect 1516 6130 1551 6164
rect 1585 6130 1617 6164
rect 1516 6074 1617 6130
rect 1516 6040 1551 6074
rect 1585 6040 1617 6074
rect 1516 5984 1617 6040
rect 1516 5950 1551 5984
rect 1585 5950 1617 5984
rect 1516 5894 1617 5950
rect 329 5831 430 5860
rect 1516 5860 1551 5894
rect 1585 5860 1617 5894
rect 1516 5831 1617 5860
rect 329 5798 1617 5831
rect 329 5764 387 5798
rect 421 5764 477 5798
rect 511 5764 567 5798
rect 601 5764 657 5798
rect 691 5764 747 5798
rect 781 5764 837 5798
rect 871 5764 927 5798
rect 961 5764 1017 5798
rect 1051 5764 1107 5798
rect 1141 5764 1197 5798
rect 1231 5764 1287 5798
rect 1321 5764 1377 5798
rect 1411 5764 1467 5798
rect 1501 5764 1617 5798
rect 329 5730 1617 5764
rect 1717 6985 3005 7018
rect 1717 6951 1775 6985
rect 1809 6951 1865 6985
rect 1899 6951 1955 6985
rect 1989 6951 2045 6985
rect 2079 6951 2135 6985
rect 2169 6951 2225 6985
rect 2259 6951 2315 6985
rect 2349 6951 2405 6985
rect 2439 6951 2495 6985
rect 2529 6951 2585 6985
rect 2619 6951 2675 6985
rect 2709 6951 2765 6985
rect 2799 6951 2855 6985
rect 2889 6951 3005 6985
rect 1717 6917 3005 6951
rect 1717 6884 1818 6917
rect 1717 6850 1752 6884
rect 1786 6850 1818 6884
rect 2904 6884 3005 6917
rect 1717 6794 1818 6850
rect 1717 6760 1752 6794
rect 1786 6760 1818 6794
rect 1717 6704 1818 6760
rect 1717 6670 1752 6704
rect 1786 6670 1818 6704
rect 1717 6614 1818 6670
rect 1717 6580 1752 6614
rect 1786 6580 1818 6614
rect 1717 6524 1818 6580
rect 1717 6490 1752 6524
rect 1786 6490 1818 6524
rect 1717 6434 1818 6490
rect 1717 6400 1752 6434
rect 1786 6400 1818 6434
rect 1717 6344 1818 6400
rect 1717 6310 1752 6344
rect 1786 6310 1818 6344
rect 1717 6254 1818 6310
rect 1717 6220 1752 6254
rect 1786 6220 1818 6254
rect 1717 6164 1818 6220
rect 1717 6130 1752 6164
rect 1786 6130 1818 6164
rect 1717 6074 1818 6130
rect 1717 6040 1752 6074
rect 1786 6040 1818 6074
rect 1717 5984 1818 6040
rect 1717 5950 1752 5984
rect 1786 5950 1818 5984
rect 1717 5894 1818 5950
rect 1717 5860 1752 5894
rect 1786 5860 1818 5894
rect 2904 6850 2939 6884
rect 2973 6850 3005 6884
rect 2904 6794 3005 6850
rect 2904 6760 2939 6794
rect 2973 6760 3005 6794
rect 2904 6704 3005 6760
rect 2904 6670 2939 6704
rect 2973 6670 3005 6704
rect 2904 6614 3005 6670
rect 2904 6580 2939 6614
rect 2973 6580 3005 6614
rect 2904 6524 3005 6580
rect 2904 6490 2939 6524
rect 2973 6490 3005 6524
rect 2904 6434 3005 6490
rect 2904 6400 2939 6434
rect 2973 6400 3005 6434
rect 2904 6344 3005 6400
rect 2904 6310 2939 6344
rect 2973 6310 3005 6344
rect 2904 6254 3005 6310
rect 2904 6220 2939 6254
rect 2973 6220 3005 6254
rect 2904 6164 3005 6220
rect 2904 6130 2939 6164
rect 2973 6130 3005 6164
rect 2904 6074 3005 6130
rect 2904 6040 2939 6074
rect 2973 6040 3005 6074
rect 2904 5984 3005 6040
rect 2904 5950 2939 5984
rect 2973 5950 3005 5984
rect 2904 5894 3005 5950
rect 1717 5831 1818 5860
rect 2904 5860 2939 5894
rect 2973 5860 3005 5894
rect 2904 5831 3005 5860
rect 1717 5798 3005 5831
rect 1717 5764 1775 5798
rect 1809 5764 1865 5798
rect 1899 5764 1955 5798
rect 1989 5764 2045 5798
rect 2079 5764 2135 5798
rect 2169 5764 2225 5798
rect 2259 5764 2315 5798
rect 2349 5764 2405 5798
rect 2439 5764 2495 5798
rect 2529 5764 2585 5798
rect 2619 5764 2675 5798
rect 2709 5764 2765 5798
rect 2799 5764 2855 5798
rect 2889 5764 3005 5798
rect 1717 5730 3005 5764
rect 3105 6985 4393 7018
rect 3105 6951 3163 6985
rect 3197 6951 3253 6985
rect 3287 6951 3343 6985
rect 3377 6951 3433 6985
rect 3467 6951 3523 6985
rect 3557 6951 3613 6985
rect 3647 6951 3703 6985
rect 3737 6951 3793 6985
rect 3827 6951 3883 6985
rect 3917 6951 3973 6985
rect 4007 6951 4063 6985
rect 4097 6951 4153 6985
rect 4187 6951 4243 6985
rect 4277 6951 4393 6985
rect 3105 6917 4393 6951
rect 3105 6884 3206 6917
rect 3105 6850 3140 6884
rect 3174 6850 3206 6884
rect 4292 6884 4393 6917
rect 3105 6794 3206 6850
rect 3105 6760 3140 6794
rect 3174 6760 3206 6794
rect 3105 6704 3206 6760
rect 3105 6670 3140 6704
rect 3174 6670 3206 6704
rect 3105 6614 3206 6670
rect 3105 6580 3140 6614
rect 3174 6580 3206 6614
rect 3105 6524 3206 6580
rect 3105 6490 3140 6524
rect 3174 6490 3206 6524
rect 3105 6434 3206 6490
rect 3105 6400 3140 6434
rect 3174 6400 3206 6434
rect 3105 6344 3206 6400
rect 3105 6310 3140 6344
rect 3174 6310 3206 6344
rect 3105 6254 3206 6310
rect 3105 6220 3140 6254
rect 3174 6220 3206 6254
rect 3105 6164 3206 6220
rect 3105 6130 3140 6164
rect 3174 6130 3206 6164
rect 3105 6074 3206 6130
rect 3105 6040 3140 6074
rect 3174 6040 3206 6074
rect 3105 5984 3206 6040
rect 3105 5950 3140 5984
rect 3174 5950 3206 5984
rect 3105 5894 3206 5950
rect 3105 5860 3140 5894
rect 3174 5860 3206 5894
rect 4292 6850 4327 6884
rect 4361 6850 4393 6884
rect 4292 6794 4393 6850
rect 4292 6760 4327 6794
rect 4361 6760 4393 6794
rect 4292 6704 4393 6760
rect 4292 6670 4327 6704
rect 4361 6670 4393 6704
rect 4292 6614 4393 6670
rect 4292 6580 4327 6614
rect 4361 6580 4393 6614
rect 4292 6524 4393 6580
rect 4292 6490 4327 6524
rect 4361 6490 4393 6524
rect 4292 6434 4393 6490
rect 4292 6400 4327 6434
rect 4361 6400 4393 6434
rect 4292 6344 4393 6400
rect 4292 6310 4327 6344
rect 4361 6310 4393 6344
rect 4292 6254 4393 6310
rect 4292 6220 4327 6254
rect 4361 6220 4393 6254
rect 4292 6164 4393 6220
rect 4292 6130 4327 6164
rect 4361 6130 4393 6164
rect 4292 6074 4393 6130
rect 4292 6040 4327 6074
rect 4361 6040 4393 6074
rect 4292 5984 4393 6040
rect 4292 5950 4327 5984
rect 4361 5950 4393 5984
rect 4292 5894 4393 5950
rect 3105 5831 3206 5860
rect 4292 5860 4327 5894
rect 4361 5860 4393 5894
rect 4292 5831 4393 5860
rect 3105 5798 4393 5831
rect 3105 5764 3163 5798
rect 3197 5764 3253 5798
rect 3287 5764 3343 5798
rect 3377 5764 3433 5798
rect 3467 5764 3523 5798
rect 3557 5764 3613 5798
rect 3647 5764 3703 5798
rect 3737 5764 3793 5798
rect 3827 5764 3883 5798
rect 3917 5764 3973 5798
rect 4007 5764 4063 5798
rect 4097 5764 4153 5798
rect 4187 5764 4243 5798
rect 4277 5764 4393 5798
rect 3105 5730 4393 5764
rect 4493 6985 5781 7018
rect 4493 6951 4551 6985
rect 4585 6951 4641 6985
rect 4675 6951 4731 6985
rect 4765 6951 4821 6985
rect 4855 6951 4911 6985
rect 4945 6951 5001 6985
rect 5035 6951 5091 6985
rect 5125 6951 5181 6985
rect 5215 6951 5271 6985
rect 5305 6951 5361 6985
rect 5395 6951 5451 6985
rect 5485 6951 5541 6985
rect 5575 6951 5631 6985
rect 5665 6951 5781 6985
rect 4493 6917 5781 6951
rect 4493 6884 4594 6917
rect 4493 6850 4528 6884
rect 4562 6850 4594 6884
rect 5680 6884 5781 6917
rect 4493 6794 4594 6850
rect 4493 6760 4528 6794
rect 4562 6760 4594 6794
rect 4493 6704 4594 6760
rect 4493 6670 4528 6704
rect 4562 6670 4594 6704
rect 4493 6614 4594 6670
rect 4493 6580 4528 6614
rect 4562 6580 4594 6614
rect 4493 6524 4594 6580
rect 4493 6490 4528 6524
rect 4562 6490 4594 6524
rect 4493 6434 4594 6490
rect 4493 6400 4528 6434
rect 4562 6400 4594 6434
rect 4493 6344 4594 6400
rect 4493 6310 4528 6344
rect 4562 6310 4594 6344
rect 4493 6254 4594 6310
rect 4493 6220 4528 6254
rect 4562 6220 4594 6254
rect 4493 6164 4594 6220
rect 4493 6130 4528 6164
rect 4562 6130 4594 6164
rect 4493 6074 4594 6130
rect 4493 6040 4528 6074
rect 4562 6040 4594 6074
rect 4493 5984 4594 6040
rect 4493 5950 4528 5984
rect 4562 5950 4594 5984
rect 4493 5894 4594 5950
rect 4493 5860 4528 5894
rect 4562 5860 4594 5894
rect 5680 6850 5715 6884
rect 5749 6850 5781 6884
rect 5680 6794 5781 6850
rect 5680 6760 5715 6794
rect 5749 6760 5781 6794
rect 5680 6704 5781 6760
rect 5680 6670 5715 6704
rect 5749 6670 5781 6704
rect 5680 6614 5781 6670
rect 5680 6580 5715 6614
rect 5749 6580 5781 6614
rect 5680 6524 5781 6580
rect 5680 6490 5715 6524
rect 5749 6490 5781 6524
rect 5680 6434 5781 6490
rect 5680 6400 5715 6434
rect 5749 6400 5781 6434
rect 5680 6344 5781 6400
rect 5680 6310 5715 6344
rect 5749 6310 5781 6344
rect 5680 6254 5781 6310
rect 5680 6220 5715 6254
rect 5749 6220 5781 6254
rect 5680 6164 5781 6220
rect 5680 6130 5715 6164
rect 5749 6130 5781 6164
rect 5680 6074 5781 6130
rect 5680 6040 5715 6074
rect 5749 6040 5781 6074
rect 5680 5984 5781 6040
rect 5680 5950 5715 5984
rect 5749 5950 5781 5984
rect 5680 5894 5781 5950
rect 4493 5831 4594 5860
rect 5680 5860 5715 5894
rect 5749 5860 5781 5894
rect 5680 5831 5781 5860
rect 4493 5798 5781 5831
rect 4493 5764 4551 5798
rect 4585 5764 4641 5798
rect 4675 5764 4731 5798
rect 4765 5764 4821 5798
rect 4855 5764 4911 5798
rect 4945 5764 5001 5798
rect 5035 5764 5091 5798
rect 5125 5764 5181 5798
rect 5215 5764 5271 5798
rect 5305 5764 5361 5798
rect 5395 5764 5451 5798
rect 5485 5764 5541 5798
rect 5575 5764 5631 5798
rect 5665 5764 5781 5798
rect 4493 5730 5781 5764
rect 5881 6985 7169 7018
rect 5881 6951 5939 6985
rect 5973 6951 6029 6985
rect 6063 6951 6119 6985
rect 6153 6951 6209 6985
rect 6243 6951 6299 6985
rect 6333 6951 6389 6985
rect 6423 6951 6479 6985
rect 6513 6951 6569 6985
rect 6603 6951 6659 6985
rect 6693 6951 6749 6985
rect 6783 6951 6839 6985
rect 6873 6951 6929 6985
rect 6963 6951 7019 6985
rect 7053 6951 7169 6985
rect 5881 6917 7169 6951
rect 5881 6884 5982 6917
rect 5881 6850 5916 6884
rect 5950 6850 5982 6884
rect 7068 6884 7169 6917
rect 5881 6794 5982 6850
rect 5881 6760 5916 6794
rect 5950 6760 5982 6794
rect 5881 6704 5982 6760
rect 5881 6670 5916 6704
rect 5950 6670 5982 6704
rect 5881 6614 5982 6670
rect 5881 6580 5916 6614
rect 5950 6580 5982 6614
rect 5881 6524 5982 6580
rect 5881 6490 5916 6524
rect 5950 6490 5982 6524
rect 5881 6434 5982 6490
rect 5881 6400 5916 6434
rect 5950 6400 5982 6434
rect 5881 6344 5982 6400
rect 5881 6310 5916 6344
rect 5950 6310 5982 6344
rect 5881 6254 5982 6310
rect 5881 6220 5916 6254
rect 5950 6220 5982 6254
rect 5881 6164 5982 6220
rect 5881 6130 5916 6164
rect 5950 6130 5982 6164
rect 5881 6074 5982 6130
rect 5881 6040 5916 6074
rect 5950 6040 5982 6074
rect 5881 5984 5982 6040
rect 5881 5950 5916 5984
rect 5950 5950 5982 5984
rect 5881 5894 5982 5950
rect 5881 5860 5916 5894
rect 5950 5860 5982 5894
rect 7068 6850 7103 6884
rect 7137 6850 7169 6884
rect 7068 6794 7169 6850
rect 7068 6760 7103 6794
rect 7137 6760 7169 6794
rect 7068 6704 7169 6760
rect 7068 6670 7103 6704
rect 7137 6670 7169 6704
rect 7068 6614 7169 6670
rect 7068 6580 7103 6614
rect 7137 6580 7169 6614
rect 7068 6524 7169 6580
rect 7068 6490 7103 6524
rect 7137 6490 7169 6524
rect 7068 6434 7169 6490
rect 7068 6400 7103 6434
rect 7137 6400 7169 6434
rect 7068 6344 7169 6400
rect 7068 6310 7103 6344
rect 7137 6310 7169 6344
rect 7068 6254 7169 6310
rect 7068 6220 7103 6254
rect 7137 6220 7169 6254
rect 7068 6164 7169 6220
rect 7068 6130 7103 6164
rect 7137 6130 7169 6164
rect 7068 6074 7169 6130
rect 7068 6040 7103 6074
rect 7137 6040 7169 6074
rect 7068 5984 7169 6040
rect 7068 5950 7103 5984
rect 7137 5950 7169 5984
rect 7068 5894 7169 5950
rect 5881 5831 5982 5860
rect 7068 5860 7103 5894
rect 7137 5860 7169 5894
rect 7068 5831 7169 5860
rect 5881 5798 7169 5831
rect 5881 5764 5939 5798
rect 5973 5764 6029 5798
rect 6063 5764 6119 5798
rect 6153 5764 6209 5798
rect 6243 5764 6299 5798
rect 6333 5764 6389 5798
rect 6423 5764 6479 5798
rect 6513 5764 6569 5798
rect 6603 5764 6659 5798
rect 6693 5764 6749 5798
rect 6783 5764 6839 5798
rect 6873 5764 6929 5798
rect 6963 5764 7019 5798
rect 7053 5764 7169 5798
rect 5881 5730 7169 5764
rect 329 5597 1617 5630
rect 329 5563 387 5597
rect 421 5563 477 5597
rect 511 5563 567 5597
rect 601 5563 657 5597
rect 691 5563 747 5597
rect 781 5563 837 5597
rect 871 5563 927 5597
rect 961 5563 1017 5597
rect 1051 5563 1107 5597
rect 1141 5563 1197 5597
rect 1231 5563 1287 5597
rect 1321 5563 1377 5597
rect 1411 5563 1467 5597
rect 1501 5563 1617 5597
rect 329 5529 1617 5563
rect 329 5496 430 5529
rect 329 5462 364 5496
rect 398 5462 430 5496
rect 1516 5496 1617 5529
rect 329 5406 430 5462
rect 329 5372 364 5406
rect 398 5372 430 5406
rect 329 5316 430 5372
rect 329 5282 364 5316
rect 398 5282 430 5316
rect 329 5226 430 5282
rect 329 5192 364 5226
rect 398 5192 430 5226
rect 329 5136 430 5192
rect 329 5102 364 5136
rect 398 5102 430 5136
rect 329 5046 430 5102
rect 329 5012 364 5046
rect 398 5012 430 5046
rect 329 4956 430 5012
rect 329 4922 364 4956
rect 398 4922 430 4956
rect 329 4866 430 4922
rect 329 4832 364 4866
rect 398 4832 430 4866
rect 329 4776 430 4832
rect 329 4742 364 4776
rect 398 4742 430 4776
rect 329 4686 430 4742
rect 329 4652 364 4686
rect 398 4652 430 4686
rect 329 4596 430 4652
rect 329 4562 364 4596
rect 398 4562 430 4596
rect 329 4506 430 4562
rect 329 4472 364 4506
rect 398 4472 430 4506
rect 1516 5462 1551 5496
rect 1585 5462 1617 5496
rect 1516 5406 1617 5462
rect 1516 5372 1551 5406
rect 1585 5372 1617 5406
rect 1516 5316 1617 5372
rect 1516 5282 1551 5316
rect 1585 5282 1617 5316
rect 1516 5226 1617 5282
rect 1516 5192 1551 5226
rect 1585 5192 1617 5226
rect 1516 5136 1617 5192
rect 1516 5102 1551 5136
rect 1585 5102 1617 5136
rect 1516 5046 1617 5102
rect 1516 5012 1551 5046
rect 1585 5012 1617 5046
rect 1516 4956 1617 5012
rect 1516 4922 1551 4956
rect 1585 4922 1617 4956
rect 1516 4866 1617 4922
rect 1516 4832 1551 4866
rect 1585 4832 1617 4866
rect 1516 4776 1617 4832
rect 1516 4742 1551 4776
rect 1585 4742 1617 4776
rect 1516 4686 1617 4742
rect 1516 4652 1551 4686
rect 1585 4652 1617 4686
rect 1516 4596 1617 4652
rect 1516 4562 1551 4596
rect 1585 4562 1617 4596
rect 1516 4506 1617 4562
rect 329 4443 430 4472
rect 1516 4472 1551 4506
rect 1585 4472 1617 4506
rect 1516 4443 1617 4472
rect 329 4410 1617 4443
rect 329 4376 387 4410
rect 421 4376 477 4410
rect 511 4376 567 4410
rect 601 4376 657 4410
rect 691 4376 747 4410
rect 781 4376 837 4410
rect 871 4376 927 4410
rect 961 4376 1017 4410
rect 1051 4376 1107 4410
rect 1141 4376 1197 4410
rect 1231 4376 1287 4410
rect 1321 4376 1377 4410
rect 1411 4376 1467 4410
rect 1501 4376 1617 4410
rect 329 4342 1617 4376
rect 1717 5597 3005 5630
rect 1717 5563 1775 5597
rect 1809 5563 1865 5597
rect 1899 5563 1955 5597
rect 1989 5563 2045 5597
rect 2079 5563 2135 5597
rect 2169 5563 2225 5597
rect 2259 5563 2315 5597
rect 2349 5563 2405 5597
rect 2439 5563 2495 5597
rect 2529 5563 2585 5597
rect 2619 5563 2675 5597
rect 2709 5563 2765 5597
rect 2799 5563 2855 5597
rect 2889 5563 3005 5597
rect 1717 5529 3005 5563
rect 1717 5496 1818 5529
rect 1717 5462 1752 5496
rect 1786 5462 1818 5496
rect 2904 5496 3005 5529
rect 1717 5406 1818 5462
rect 1717 5372 1752 5406
rect 1786 5372 1818 5406
rect 1717 5316 1818 5372
rect 1717 5282 1752 5316
rect 1786 5282 1818 5316
rect 1717 5226 1818 5282
rect 1717 5192 1752 5226
rect 1786 5192 1818 5226
rect 1717 5136 1818 5192
rect 1717 5102 1752 5136
rect 1786 5102 1818 5136
rect 1717 5046 1818 5102
rect 1717 5012 1752 5046
rect 1786 5012 1818 5046
rect 1717 4956 1818 5012
rect 1717 4922 1752 4956
rect 1786 4922 1818 4956
rect 1717 4866 1818 4922
rect 1717 4832 1752 4866
rect 1786 4832 1818 4866
rect 1717 4776 1818 4832
rect 1717 4742 1752 4776
rect 1786 4742 1818 4776
rect 1717 4686 1818 4742
rect 1717 4652 1752 4686
rect 1786 4652 1818 4686
rect 1717 4596 1818 4652
rect 1717 4562 1752 4596
rect 1786 4562 1818 4596
rect 1717 4506 1818 4562
rect 1717 4472 1752 4506
rect 1786 4472 1818 4506
rect 2904 5462 2939 5496
rect 2973 5462 3005 5496
rect 2904 5406 3005 5462
rect 2904 5372 2939 5406
rect 2973 5372 3005 5406
rect 2904 5316 3005 5372
rect 2904 5282 2939 5316
rect 2973 5282 3005 5316
rect 2904 5226 3005 5282
rect 2904 5192 2939 5226
rect 2973 5192 3005 5226
rect 2904 5136 3005 5192
rect 2904 5102 2939 5136
rect 2973 5102 3005 5136
rect 2904 5046 3005 5102
rect 2904 5012 2939 5046
rect 2973 5012 3005 5046
rect 2904 4956 3005 5012
rect 2904 4922 2939 4956
rect 2973 4922 3005 4956
rect 2904 4866 3005 4922
rect 2904 4832 2939 4866
rect 2973 4832 3005 4866
rect 2904 4776 3005 4832
rect 2904 4742 2939 4776
rect 2973 4742 3005 4776
rect 2904 4686 3005 4742
rect 2904 4652 2939 4686
rect 2973 4652 3005 4686
rect 2904 4596 3005 4652
rect 2904 4562 2939 4596
rect 2973 4562 3005 4596
rect 2904 4506 3005 4562
rect 1717 4443 1818 4472
rect 2904 4472 2939 4506
rect 2973 4472 3005 4506
rect 2904 4443 3005 4472
rect 1717 4410 3005 4443
rect 1717 4376 1775 4410
rect 1809 4376 1865 4410
rect 1899 4376 1955 4410
rect 1989 4376 2045 4410
rect 2079 4376 2135 4410
rect 2169 4376 2225 4410
rect 2259 4376 2315 4410
rect 2349 4376 2405 4410
rect 2439 4376 2495 4410
rect 2529 4376 2585 4410
rect 2619 4376 2675 4410
rect 2709 4376 2765 4410
rect 2799 4376 2855 4410
rect 2889 4376 3005 4410
rect 1717 4342 3005 4376
rect 3105 5597 4393 5630
rect 3105 5563 3163 5597
rect 3197 5563 3253 5597
rect 3287 5563 3343 5597
rect 3377 5563 3433 5597
rect 3467 5563 3523 5597
rect 3557 5563 3613 5597
rect 3647 5563 3703 5597
rect 3737 5563 3793 5597
rect 3827 5563 3883 5597
rect 3917 5563 3973 5597
rect 4007 5563 4063 5597
rect 4097 5563 4153 5597
rect 4187 5563 4243 5597
rect 4277 5563 4393 5597
rect 3105 5529 4393 5563
rect 3105 5496 3206 5529
rect 3105 5462 3140 5496
rect 3174 5462 3206 5496
rect 4292 5496 4393 5529
rect 3105 5406 3206 5462
rect 3105 5372 3140 5406
rect 3174 5372 3206 5406
rect 3105 5316 3206 5372
rect 3105 5282 3140 5316
rect 3174 5282 3206 5316
rect 3105 5226 3206 5282
rect 3105 5192 3140 5226
rect 3174 5192 3206 5226
rect 3105 5136 3206 5192
rect 3105 5102 3140 5136
rect 3174 5102 3206 5136
rect 3105 5046 3206 5102
rect 3105 5012 3140 5046
rect 3174 5012 3206 5046
rect 3105 4956 3206 5012
rect 3105 4922 3140 4956
rect 3174 4922 3206 4956
rect 3105 4866 3206 4922
rect 3105 4832 3140 4866
rect 3174 4832 3206 4866
rect 3105 4776 3206 4832
rect 3105 4742 3140 4776
rect 3174 4742 3206 4776
rect 3105 4686 3206 4742
rect 3105 4652 3140 4686
rect 3174 4652 3206 4686
rect 3105 4596 3206 4652
rect 3105 4562 3140 4596
rect 3174 4562 3206 4596
rect 3105 4506 3206 4562
rect 3105 4472 3140 4506
rect 3174 4472 3206 4506
rect 4292 5462 4327 5496
rect 4361 5462 4393 5496
rect 4292 5406 4393 5462
rect 4292 5372 4327 5406
rect 4361 5372 4393 5406
rect 4292 5316 4393 5372
rect 4292 5282 4327 5316
rect 4361 5282 4393 5316
rect 4292 5226 4393 5282
rect 4292 5192 4327 5226
rect 4361 5192 4393 5226
rect 4292 5136 4393 5192
rect 4292 5102 4327 5136
rect 4361 5102 4393 5136
rect 4292 5046 4393 5102
rect 4292 5012 4327 5046
rect 4361 5012 4393 5046
rect 4292 4956 4393 5012
rect 4292 4922 4327 4956
rect 4361 4922 4393 4956
rect 4292 4866 4393 4922
rect 4292 4832 4327 4866
rect 4361 4832 4393 4866
rect 4292 4776 4393 4832
rect 4292 4742 4327 4776
rect 4361 4742 4393 4776
rect 4292 4686 4393 4742
rect 4292 4652 4327 4686
rect 4361 4652 4393 4686
rect 4292 4596 4393 4652
rect 4292 4562 4327 4596
rect 4361 4562 4393 4596
rect 4292 4506 4393 4562
rect 3105 4443 3206 4472
rect 4292 4472 4327 4506
rect 4361 4472 4393 4506
rect 4292 4443 4393 4472
rect 3105 4410 4393 4443
rect 3105 4376 3163 4410
rect 3197 4376 3253 4410
rect 3287 4376 3343 4410
rect 3377 4376 3433 4410
rect 3467 4376 3523 4410
rect 3557 4376 3613 4410
rect 3647 4376 3703 4410
rect 3737 4376 3793 4410
rect 3827 4376 3883 4410
rect 3917 4376 3973 4410
rect 4007 4376 4063 4410
rect 4097 4376 4153 4410
rect 4187 4376 4243 4410
rect 4277 4376 4393 4410
rect 3105 4342 4393 4376
rect 4493 5597 5781 5630
rect 4493 5563 4551 5597
rect 4585 5563 4641 5597
rect 4675 5563 4731 5597
rect 4765 5563 4821 5597
rect 4855 5563 4911 5597
rect 4945 5563 5001 5597
rect 5035 5563 5091 5597
rect 5125 5563 5181 5597
rect 5215 5563 5271 5597
rect 5305 5563 5361 5597
rect 5395 5563 5451 5597
rect 5485 5563 5541 5597
rect 5575 5563 5631 5597
rect 5665 5563 5781 5597
rect 4493 5529 5781 5563
rect 4493 5496 4594 5529
rect 4493 5462 4528 5496
rect 4562 5462 4594 5496
rect 5680 5496 5781 5529
rect 4493 5406 4594 5462
rect 4493 5372 4528 5406
rect 4562 5372 4594 5406
rect 4493 5316 4594 5372
rect 4493 5282 4528 5316
rect 4562 5282 4594 5316
rect 4493 5226 4594 5282
rect 4493 5192 4528 5226
rect 4562 5192 4594 5226
rect 4493 5136 4594 5192
rect 4493 5102 4528 5136
rect 4562 5102 4594 5136
rect 4493 5046 4594 5102
rect 4493 5012 4528 5046
rect 4562 5012 4594 5046
rect 4493 4956 4594 5012
rect 4493 4922 4528 4956
rect 4562 4922 4594 4956
rect 4493 4866 4594 4922
rect 4493 4832 4528 4866
rect 4562 4832 4594 4866
rect 4493 4776 4594 4832
rect 4493 4742 4528 4776
rect 4562 4742 4594 4776
rect 4493 4686 4594 4742
rect 4493 4652 4528 4686
rect 4562 4652 4594 4686
rect 4493 4596 4594 4652
rect 4493 4562 4528 4596
rect 4562 4562 4594 4596
rect 4493 4506 4594 4562
rect 4493 4472 4528 4506
rect 4562 4472 4594 4506
rect 5680 5462 5715 5496
rect 5749 5462 5781 5496
rect 5680 5406 5781 5462
rect 5680 5372 5715 5406
rect 5749 5372 5781 5406
rect 5680 5316 5781 5372
rect 5680 5282 5715 5316
rect 5749 5282 5781 5316
rect 5680 5226 5781 5282
rect 5680 5192 5715 5226
rect 5749 5192 5781 5226
rect 5680 5136 5781 5192
rect 5680 5102 5715 5136
rect 5749 5102 5781 5136
rect 5680 5046 5781 5102
rect 5680 5012 5715 5046
rect 5749 5012 5781 5046
rect 5680 4956 5781 5012
rect 5680 4922 5715 4956
rect 5749 4922 5781 4956
rect 5680 4866 5781 4922
rect 5680 4832 5715 4866
rect 5749 4832 5781 4866
rect 5680 4776 5781 4832
rect 5680 4742 5715 4776
rect 5749 4742 5781 4776
rect 5680 4686 5781 4742
rect 5680 4652 5715 4686
rect 5749 4652 5781 4686
rect 5680 4596 5781 4652
rect 5680 4562 5715 4596
rect 5749 4562 5781 4596
rect 5680 4506 5781 4562
rect 4493 4443 4594 4472
rect 5680 4472 5715 4506
rect 5749 4472 5781 4506
rect 5680 4443 5781 4472
rect 4493 4410 5781 4443
rect 4493 4376 4551 4410
rect 4585 4376 4641 4410
rect 4675 4376 4731 4410
rect 4765 4376 4821 4410
rect 4855 4376 4911 4410
rect 4945 4376 5001 4410
rect 5035 4376 5091 4410
rect 5125 4376 5181 4410
rect 5215 4376 5271 4410
rect 5305 4376 5361 4410
rect 5395 4376 5451 4410
rect 5485 4376 5541 4410
rect 5575 4376 5631 4410
rect 5665 4376 5781 4410
rect 4493 4342 5781 4376
rect 5881 5597 7169 5630
rect 5881 5563 5939 5597
rect 5973 5563 6029 5597
rect 6063 5563 6119 5597
rect 6153 5563 6209 5597
rect 6243 5563 6299 5597
rect 6333 5563 6389 5597
rect 6423 5563 6479 5597
rect 6513 5563 6569 5597
rect 6603 5563 6659 5597
rect 6693 5563 6749 5597
rect 6783 5563 6839 5597
rect 6873 5563 6929 5597
rect 6963 5563 7019 5597
rect 7053 5563 7169 5597
rect 5881 5529 7169 5563
rect 5881 5496 5982 5529
rect 5881 5462 5916 5496
rect 5950 5462 5982 5496
rect 7068 5496 7169 5529
rect 5881 5406 5982 5462
rect 5881 5372 5916 5406
rect 5950 5372 5982 5406
rect 5881 5316 5982 5372
rect 5881 5282 5916 5316
rect 5950 5282 5982 5316
rect 5881 5226 5982 5282
rect 5881 5192 5916 5226
rect 5950 5192 5982 5226
rect 5881 5136 5982 5192
rect 5881 5102 5916 5136
rect 5950 5102 5982 5136
rect 5881 5046 5982 5102
rect 5881 5012 5916 5046
rect 5950 5012 5982 5046
rect 5881 4956 5982 5012
rect 5881 4922 5916 4956
rect 5950 4922 5982 4956
rect 5881 4866 5982 4922
rect 5881 4832 5916 4866
rect 5950 4832 5982 4866
rect 5881 4776 5982 4832
rect 5881 4742 5916 4776
rect 5950 4742 5982 4776
rect 5881 4686 5982 4742
rect 5881 4652 5916 4686
rect 5950 4652 5982 4686
rect 5881 4596 5982 4652
rect 5881 4562 5916 4596
rect 5950 4562 5982 4596
rect 5881 4506 5982 4562
rect 5881 4472 5916 4506
rect 5950 4472 5982 4506
rect 7068 5462 7103 5496
rect 7137 5462 7169 5496
rect 7068 5406 7169 5462
rect 7068 5372 7103 5406
rect 7137 5372 7169 5406
rect 7068 5316 7169 5372
rect 7068 5282 7103 5316
rect 7137 5282 7169 5316
rect 7068 5226 7169 5282
rect 7068 5192 7103 5226
rect 7137 5192 7169 5226
rect 7068 5136 7169 5192
rect 7068 5102 7103 5136
rect 7137 5102 7169 5136
rect 7068 5046 7169 5102
rect 7068 5012 7103 5046
rect 7137 5012 7169 5046
rect 7068 4956 7169 5012
rect 7068 4922 7103 4956
rect 7137 4922 7169 4956
rect 7068 4866 7169 4922
rect 7068 4832 7103 4866
rect 7137 4832 7169 4866
rect 7068 4776 7169 4832
rect 7068 4742 7103 4776
rect 7137 4742 7169 4776
rect 7068 4686 7169 4742
rect 7068 4652 7103 4686
rect 7137 4652 7169 4686
rect 7068 4596 7169 4652
rect 7068 4562 7103 4596
rect 7137 4562 7169 4596
rect 7068 4506 7169 4562
rect 5881 4443 5982 4472
rect 7068 4472 7103 4506
rect 7137 4472 7169 4506
rect 7068 4443 7169 4472
rect 5881 4410 7169 4443
rect 5881 4376 5939 4410
rect 5973 4376 6029 4410
rect 6063 4376 6119 4410
rect 6153 4376 6209 4410
rect 6243 4376 6299 4410
rect 6333 4376 6389 4410
rect 6423 4376 6479 4410
rect 6513 4376 6569 4410
rect 6603 4376 6659 4410
rect 6693 4376 6749 4410
rect 6783 4376 6839 4410
rect 6873 4376 6929 4410
rect 6963 4376 7019 4410
rect 7053 4376 7169 4410
rect 5881 4342 7169 4376
rect 329 4209 1617 4242
rect 329 4175 387 4209
rect 421 4175 477 4209
rect 511 4175 567 4209
rect 601 4175 657 4209
rect 691 4175 747 4209
rect 781 4175 837 4209
rect 871 4175 927 4209
rect 961 4175 1017 4209
rect 1051 4175 1107 4209
rect 1141 4175 1197 4209
rect 1231 4175 1287 4209
rect 1321 4175 1377 4209
rect 1411 4175 1467 4209
rect 1501 4175 1617 4209
rect 329 4141 1617 4175
rect 329 4108 430 4141
rect 329 4074 364 4108
rect 398 4074 430 4108
rect 1516 4108 1617 4141
rect 329 4018 430 4074
rect 329 3984 364 4018
rect 398 3984 430 4018
rect 329 3928 430 3984
rect 329 3894 364 3928
rect 398 3894 430 3928
rect 329 3838 430 3894
rect 329 3804 364 3838
rect 398 3804 430 3838
rect 329 3748 430 3804
rect 329 3714 364 3748
rect 398 3714 430 3748
rect 329 3658 430 3714
rect 329 3624 364 3658
rect 398 3624 430 3658
rect 329 3568 430 3624
rect 329 3534 364 3568
rect 398 3534 430 3568
rect 329 3478 430 3534
rect 329 3444 364 3478
rect 398 3444 430 3478
rect 329 3388 430 3444
rect 329 3354 364 3388
rect 398 3354 430 3388
rect 329 3298 430 3354
rect 329 3264 364 3298
rect 398 3264 430 3298
rect 329 3208 430 3264
rect 329 3174 364 3208
rect 398 3174 430 3208
rect 329 3118 430 3174
rect 329 3084 364 3118
rect 398 3084 430 3118
rect 1516 4074 1551 4108
rect 1585 4074 1617 4108
rect 1516 4018 1617 4074
rect 1516 3984 1551 4018
rect 1585 3984 1617 4018
rect 1516 3928 1617 3984
rect 1516 3894 1551 3928
rect 1585 3894 1617 3928
rect 1516 3838 1617 3894
rect 1516 3804 1551 3838
rect 1585 3804 1617 3838
rect 1516 3748 1617 3804
rect 1516 3714 1551 3748
rect 1585 3714 1617 3748
rect 1516 3658 1617 3714
rect 1516 3624 1551 3658
rect 1585 3624 1617 3658
rect 1516 3568 1617 3624
rect 1516 3534 1551 3568
rect 1585 3534 1617 3568
rect 1516 3478 1617 3534
rect 1516 3444 1551 3478
rect 1585 3444 1617 3478
rect 1516 3388 1617 3444
rect 1516 3354 1551 3388
rect 1585 3354 1617 3388
rect 1516 3298 1617 3354
rect 1516 3264 1551 3298
rect 1585 3264 1617 3298
rect 1516 3208 1617 3264
rect 1516 3174 1551 3208
rect 1585 3174 1617 3208
rect 1516 3118 1617 3174
rect 329 3055 430 3084
rect 1516 3084 1551 3118
rect 1585 3084 1617 3118
rect 1516 3055 1617 3084
rect 329 3022 1617 3055
rect 329 2988 387 3022
rect 421 2988 477 3022
rect 511 2988 567 3022
rect 601 2988 657 3022
rect 691 2988 747 3022
rect 781 2988 837 3022
rect 871 2988 927 3022
rect 961 2988 1017 3022
rect 1051 2988 1107 3022
rect 1141 2988 1197 3022
rect 1231 2988 1287 3022
rect 1321 2988 1377 3022
rect 1411 2988 1467 3022
rect 1501 2988 1617 3022
rect 329 2954 1617 2988
rect 1717 4209 3005 4242
rect 1717 4175 1775 4209
rect 1809 4175 1865 4209
rect 1899 4175 1955 4209
rect 1989 4175 2045 4209
rect 2079 4175 2135 4209
rect 2169 4175 2225 4209
rect 2259 4175 2315 4209
rect 2349 4175 2405 4209
rect 2439 4175 2495 4209
rect 2529 4175 2585 4209
rect 2619 4175 2675 4209
rect 2709 4175 2765 4209
rect 2799 4175 2855 4209
rect 2889 4175 3005 4209
rect 1717 4141 3005 4175
rect 1717 4108 1818 4141
rect 1717 4074 1752 4108
rect 1786 4074 1818 4108
rect 2904 4108 3005 4141
rect 1717 4018 1818 4074
rect 1717 3984 1752 4018
rect 1786 3984 1818 4018
rect 1717 3928 1818 3984
rect 1717 3894 1752 3928
rect 1786 3894 1818 3928
rect 1717 3838 1818 3894
rect 1717 3804 1752 3838
rect 1786 3804 1818 3838
rect 1717 3748 1818 3804
rect 1717 3714 1752 3748
rect 1786 3714 1818 3748
rect 1717 3658 1818 3714
rect 1717 3624 1752 3658
rect 1786 3624 1818 3658
rect 1717 3568 1818 3624
rect 1717 3534 1752 3568
rect 1786 3534 1818 3568
rect 1717 3478 1818 3534
rect 1717 3444 1752 3478
rect 1786 3444 1818 3478
rect 1717 3388 1818 3444
rect 1717 3354 1752 3388
rect 1786 3354 1818 3388
rect 1717 3298 1818 3354
rect 1717 3264 1752 3298
rect 1786 3264 1818 3298
rect 1717 3208 1818 3264
rect 1717 3174 1752 3208
rect 1786 3174 1818 3208
rect 1717 3118 1818 3174
rect 1717 3084 1752 3118
rect 1786 3084 1818 3118
rect 2904 4074 2939 4108
rect 2973 4074 3005 4108
rect 2904 4018 3005 4074
rect 2904 3984 2939 4018
rect 2973 3984 3005 4018
rect 2904 3928 3005 3984
rect 2904 3894 2939 3928
rect 2973 3894 3005 3928
rect 2904 3838 3005 3894
rect 2904 3804 2939 3838
rect 2973 3804 3005 3838
rect 2904 3748 3005 3804
rect 2904 3714 2939 3748
rect 2973 3714 3005 3748
rect 2904 3658 3005 3714
rect 2904 3624 2939 3658
rect 2973 3624 3005 3658
rect 2904 3568 3005 3624
rect 2904 3534 2939 3568
rect 2973 3534 3005 3568
rect 2904 3478 3005 3534
rect 2904 3444 2939 3478
rect 2973 3444 3005 3478
rect 2904 3388 3005 3444
rect 2904 3354 2939 3388
rect 2973 3354 3005 3388
rect 2904 3298 3005 3354
rect 2904 3264 2939 3298
rect 2973 3264 3005 3298
rect 2904 3208 3005 3264
rect 2904 3174 2939 3208
rect 2973 3174 3005 3208
rect 2904 3118 3005 3174
rect 1717 3055 1818 3084
rect 2904 3084 2939 3118
rect 2973 3084 3005 3118
rect 2904 3055 3005 3084
rect 1717 3022 3005 3055
rect 1717 2988 1775 3022
rect 1809 2988 1865 3022
rect 1899 2988 1955 3022
rect 1989 2988 2045 3022
rect 2079 2988 2135 3022
rect 2169 2988 2225 3022
rect 2259 2988 2315 3022
rect 2349 2988 2405 3022
rect 2439 2988 2495 3022
rect 2529 2988 2585 3022
rect 2619 2988 2675 3022
rect 2709 2988 2765 3022
rect 2799 2988 2855 3022
rect 2889 2988 3005 3022
rect 1717 2954 3005 2988
rect 3105 4209 4393 4242
rect 3105 4175 3163 4209
rect 3197 4175 3253 4209
rect 3287 4175 3343 4209
rect 3377 4175 3433 4209
rect 3467 4175 3523 4209
rect 3557 4175 3613 4209
rect 3647 4175 3703 4209
rect 3737 4175 3793 4209
rect 3827 4175 3883 4209
rect 3917 4175 3973 4209
rect 4007 4175 4063 4209
rect 4097 4175 4153 4209
rect 4187 4175 4243 4209
rect 4277 4175 4393 4209
rect 3105 4141 4393 4175
rect 3105 4108 3206 4141
rect 3105 4074 3140 4108
rect 3174 4074 3206 4108
rect 4292 4108 4393 4141
rect 3105 4018 3206 4074
rect 3105 3984 3140 4018
rect 3174 3984 3206 4018
rect 3105 3928 3206 3984
rect 3105 3894 3140 3928
rect 3174 3894 3206 3928
rect 3105 3838 3206 3894
rect 3105 3804 3140 3838
rect 3174 3804 3206 3838
rect 3105 3748 3206 3804
rect 3105 3714 3140 3748
rect 3174 3714 3206 3748
rect 3105 3658 3206 3714
rect 3105 3624 3140 3658
rect 3174 3624 3206 3658
rect 3105 3568 3206 3624
rect 3105 3534 3140 3568
rect 3174 3534 3206 3568
rect 3105 3478 3206 3534
rect 3105 3444 3140 3478
rect 3174 3444 3206 3478
rect 3105 3388 3206 3444
rect 3105 3354 3140 3388
rect 3174 3354 3206 3388
rect 3105 3298 3206 3354
rect 3105 3264 3140 3298
rect 3174 3264 3206 3298
rect 3105 3208 3206 3264
rect 3105 3174 3140 3208
rect 3174 3174 3206 3208
rect 3105 3118 3206 3174
rect 3105 3084 3140 3118
rect 3174 3084 3206 3118
rect 4292 4074 4327 4108
rect 4361 4074 4393 4108
rect 4292 4018 4393 4074
rect 4292 3984 4327 4018
rect 4361 3984 4393 4018
rect 4292 3928 4393 3984
rect 4292 3894 4327 3928
rect 4361 3894 4393 3928
rect 4292 3838 4393 3894
rect 4292 3804 4327 3838
rect 4361 3804 4393 3838
rect 4292 3748 4393 3804
rect 4292 3714 4327 3748
rect 4361 3714 4393 3748
rect 4292 3658 4393 3714
rect 4292 3624 4327 3658
rect 4361 3624 4393 3658
rect 4292 3568 4393 3624
rect 4292 3534 4327 3568
rect 4361 3534 4393 3568
rect 4292 3478 4393 3534
rect 4292 3444 4327 3478
rect 4361 3444 4393 3478
rect 4292 3388 4393 3444
rect 4292 3354 4327 3388
rect 4361 3354 4393 3388
rect 4292 3298 4393 3354
rect 4292 3264 4327 3298
rect 4361 3264 4393 3298
rect 4292 3208 4393 3264
rect 4292 3174 4327 3208
rect 4361 3174 4393 3208
rect 4292 3118 4393 3174
rect 3105 3055 3206 3084
rect 4292 3084 4327 3118
rect 4361 3084 4393 3118
rect 4292 3055 4393 3084
rect 3105 3022 4393 3055
rect 3105 2988 3163 3022
rect 3197 2988 3253 3022
rect 3287 2988 3343 3022
rect 3377 2988 3433 3022
rect 3467 2988 3523 3022
rect 3557 2988 3613 3022
rect 3647 2988 3703 3022
rect 3737 2988 3793 3022
rect 3827 2988 3883 3022
rect 3917 2988 3973 3022
rect 4007 2988 4063 3022
rect 4097 2988 4153 3022
rect 4187 2988 4243 3022
rect 4277 2988 4393 3022
rect 3105 2954 4393 2988
rect 4493 4209 5781 4242
rect 4493 4175 4551 4209
rect 4585 4175 4641 4209
rect 4675 4175 4731 4209
rect 4765 4175 4821 4209
rect 4855 4175 4911 4209
rect 4945 4175 5001 4209
rect 5035 4175 5091 4209
rect 5125 4175 5181 4209
rect 5215 4175 5271 4209
rect 5305 4175 5361 4209
rect 5395 4175 5451 4209
rect 5485 4175 5541 4209
rect 5575 4175 5631 4209
rect 5665 4175 5781 4209
rect 4493 4141 5781 4175
rect 4493 4108 4594 4141
rect 4493 4074 4528 4108
rect 4562 4074 4594 4108
rect 5680 4108 5781 4141
rect 4493 4018 4594 4074
rect 4493 3984 4528 4018
rect 4562 3984 4594 4018
rect 4493 3928 4594 3984
rect 4493 3894 4528 3928
rect 4562 3894 4594 3928
rect 4493 3838 4594 3894
rect 4493 3804 4528 3838
rect 4562 3804 4594 3838
rect 4493 3748 4594 3804
rect 4493 3714 4528 3748
rect 4562 3714 4594 3748
rect 4493 3658 4594 3714
rect 4493 3624 4528 3658
rect 4562 3624 4594 3658
rect 4493 3568 4594 3624
rect 4493 3534 4528 3568
rect 4562 3534 4594 3568
rect 4493 3478 4594 3534
rect 4493 3444 4528 3478
rect 4562 3444 4594 3478
rect 4493 3388 4594 3444
rect 4493 3354 4528 3388
rect 4562 3354 4594 3388
rect 4493 3298 4594 3354
rect 4493 3264 4528 3298
rect 4562 3264 4594 3298
rect 4493 3208 4594 3264
rect 4493 3174 4528 3208
rect 4562 3174 4594 3208
rect 4493 3118 4594 3174
rect 4493 3084 4528 3118
rect 4562 3084 4594 3118
rect 5680 4074 5715 4108
rect 5749 4074 5781 4108
rect 5680 4018 5781 4074
rect 5680 3984 5715 4018
rect 5749 3984 5781 4018
rect 5680 3928 5781 3984
rect 5680 3894 5715 3928
rect 5749 3894 5781 3928
rect 5680 3838 5781 3894
rect 5680 3804 5715 3838
rect 5749 3804 5781 3838
rect 5680 3748 5781 3804
rect 5680 3714 5715 3748
rect 5749 3714 5781 3748
rect 5680 3658 5781 3714
rect 5680 3624 5715 3658
rect 5749 3624 5781 3658
rect 5680 3568 5781 3624
rect 5680 3534 5715 3568
rect 5749 3534 5781 3568
rect 5680 3478 5781 3534
rect 5680 3444 5715 3478
rect 5749 3444 5781 3478
rect 5680 3388 5781 3444
rect 5680 3354 5715 3388
rect 5749 3354 5781 3388
rect 5680 3298 5781 3354
rect 5680 3264 5715 3298
rect 5749 3264 5781 3298
rect 5680 3208 5781 3264
rect 5680 3174 5715 3208
rect 5749 3174 5781 3208
rect 5680 3118 5781 3174
rect 4493 3055 4594 3084
rect 5680 3084 5715 3118
rect 5749 3084 5781 3118
rect 5680 3055 5781 3084
rect 4493 3022 5781 3055
rect 4493 2988 4551 3022
rect 4585 2988 4641 3022
rect 4675 2988 4731 3022
rect 4765 2988 4821 3022
rect 4855 2988 4911 3022
rect 4945 2988 5001 3022
rect 5035 2988 5091 3022
rect 5125 2988 5181 3022
rect 5215 2988 5271 3022
rect 5305 2988 5361 3022
rect 5395 2988 5451 3022
rect 5485 2988 5541 3022
rect 5575 2988 5631 3022
rect 5665 2988 5781 3022
rect 4493 2954 5781 2988
rect 5881 4209 7169 4242
rect 5881 4175 5939 4209
rect 5973 4175 6029 4209
rect 6063 4175 6119 4209
rect 6153 4175 6209 4209
rect 6243 4175 6299 4209
rect 6333 4175 6389 4209
rect 6423 4175 6479 4209
rect 6513 4175 6569 4209
rect 6603 4175 6659 4209
rect 6693 4175 6749 4209
rect 6783 4175 6839 4209
rect 6873 4175 6929 4209
rect 6963 4175 7019 4209
rect 7053 4175 7169 4209
rect 5881 4141 7169 4175
rect 5881 4108 5982 4141
rect 5881 4074 5916 4108
rect 5950 4074 5982 4108
rect 7068 4108 7169 4141
rect 5881 4018 5982 4074
rect 5881 3984 5916 4018
rect 5950 3984 5982 4018
rect 5881 3928 5982 3984
rect 5881 3894 5916 3928
rect 5950 3894 5982 3928
rect 5881 3838 5982 3894
rect 5881 3804 5916 3838
rect 5950 3804 5982 3838
rect 5881 3748 5982 3804
rect 5881 3714 5916 3748
rect 5950 3714 5982 3748
rect 5881 3658 5982 3714
rect 5881 3624 5916 3658
rect 5950 3624 5982 3658
rect 5881 3568 5982 3624
rect 5881 3534 5916 3568
rect 5950 3534 5982 3568
rect 5881 3478 5982 3534
rect 5881 3444 5916 3478
rect 5950 3444 5982 3478
rect 5881 3388 5982 3444
rect 5881 3354 5916 3388
rect 5950 3354 5982 3388
rect 5881 3298 5982 3354
rect 5881 3264 5916 3298
rect 5950 3264 5982 3298
rect 5881 3208 5982 3264
rect 5881 3174 5916 3208
rect 5950 3174 5982 3208
rect 5881 3118 5982 3174
rect 5881 3084 5916 3118
rect 5950 3084 5982 3118
rect 7068 4074 7103 4108
rect 7137 4074 7169 4108
rect 7068 4018 7169 4074
rect 7068 3984 7103 4018
rect 7137 3984 7169 4018
rect 7068 3928 7169 3984
rect 7068 3894 7103 3928
rect 7137 3894 7169 3928
rect 7068 3838 7169 3894
rect 7068 3804 7103 3838
rect 7137 3804 7169 3838
rect 7068 3748 7169 3804
rect 7068 3714 7103 3748
rect 7137 3714 7169 3748
rect 7068 3658 7169 3714
rect 7068 3624 7103 3658
rect 7137 3624 7169 3658
rect 7068 3568 7169 3624
rect 7068 3534 7103 3568
rect 7137 3534 7169 3568
rect 7068 3478 7169 3534
rect 7068 3444 7103 3478
rect 7137 3444 7169 3478
rect 7068 3388 7169 3444
rect 7068 3354 7103 3388
rect 7137 3354 7169 3388
rect 7068 3298 7169 3354
rect 7068 3264 7103 3298
rect 7137 3264 7169 3298
rect 7068 3208 7169 3264
rect 7068 3174 7103 3208
rect 7137 3174 7169 3208
rect 7068 3118 7169 3174
rect 5881 3055 5982 3084
rect 7068 3084 7103 3118
rect 7137 3084 7169 3118
rect 7068 3055 7169 3084
rect 5881 3022 7169 3055
rect 5881 2988 5939 3022
rect 5973 2988 6029 3022
rect 6063 2988 6119 3022
rect 6153 2988 6209 3022
rect 6243 2988 6299 3022
rect 6333 2988 6389 3022
rect 6423 2988 6479 3022
rect 6513 2988 6569 3022
rect 6603 2988 6659 3022
rect 6693 2988 6749 3022
rect 6783 2988 6839 3022
rect 6873 2988 6929 3022
rect 6963 2988 7019 3022
rect 7053 2988 7169 3022
rect 5881 2954 7169 2988
rect 329 2821 1617 2854
rect 329 2787 387 2821
rect 421 2787 477 2821
rect 511 2787 567 2821
rect 601 2787 657 2821
rect 691 2787 747 2821
rect 781 2787 837 2821
rect 871 2787 927 2821
rect 961 2787 1017 2821
rect 1051 2787 1107 2821
rect 1141 2787 1197 2821
rect 1231 2787 1287 2821
rect 1321 2787 1377 2821
rect 1411 2787 1467 2821
rect 1501 2787 1617 2821
rect 329 2753 1617 2787
rect 329 2720 430 2753
rect 329 2686 364 2720
rect 398 2686 430 2720
rect 1516 2720 1617 2753
rect 329 2630 430 2686
rect 329 2596 364 2630
rect 398 2596 430 2630
rect 329 2540 430 2596
rect 329 2506 364 2540
rect 398 2506 430 2540
rect 329 2450 430 2506
rect 329 2416 364 2450
rect 398 2416 430 2450
rect 329 2360 430 2416
rect 329 2326 364 2360
rect 398 2326 430 2360
rect 329 2270 430 2326
rect 329 2236 364 2270
rect 398 2236 430 2270
rect 329 2180 430 2236
rect 329 2146 364 2180
rect 398 2146 430 2180
rect 329 2090 430 2146
rect 329 2056 364 2090
rect 398 2056 430 2090
rect 329 2000 430 2056
rect 329 1966 364 2000
rect 398 1966 430 2000
rect 329 1910 430 1966
rect 329 1876 364 1910
rect 398 1876 430 1910
rect 329 1820 430 1876
rect 329 1786 364 1820
rect 398 1786 430 1820
rect 329 1730 430 1786
rect 329 1696 364 1730
rect 398 1696 430 1730
rect 1516 2686 1551 2720
rect 1585 2686 1617 2720
rect 1516 2630 1617 2686
rect 1516 2596 1551 2630
rect 1585 2596 1617 2630
rect 1516 2540 1617 2596
rect 1516 2506 1551 2540
rect 1585 2506 1617 2540
rect 1516 2450 1617 2506
rect 1516 2416 1551 2450
rect 1585 2416 1617 2450
rect 1516 2360 1617 2416
rect 1516 2326 1551 2360
rect 1585 2326 1617 2360
rect 1516 2270 1617 2326
rect 1516 2236 1551 2270
rect 1585 2236 1617 2270
rect 1516 2180 1617 2236
rect 1516 2146 1551 2180
rect 1585 2146 1617 2180
rect 1516 2090 1617 2146
rect 1516 2056 1551 2090
rect 1585 2056 1617 2090
rect 1516 2000 1617 2056
rect 1516 1966 1551 2000
rect 1585 1966 1617 2000
rect 1516 1910 1617 1966
rect 1516 1876 1551 1910
rect 1585 1876 1617 1910
rect 1516 1820 1617 1876
rect 1516 1786 1551 1820
rect 1585 1786 1617 1820
rect 1516 1730 1617 1786
rect 329 1667 430 1696
rect 1516 1696 1551 1730
rect 1585 1696 1617 1730
rect 1516 1667 1617 1696
rect 329 1634 1617 1667
rect 329 1600 387 1634
rect 421 1600 477 1634
rect 511 1600 567 1634
rect 601 1600 657 1634
rect 691 1600 747 1634
rect 781 1600 837 1634
rect 871 1600 927 1634
rect 961 1600 1017 1634
rect 1051 1600 1107 1634
rect 1141 1600 1197 1634
rect 1231 1600 1287 1634
rect 1321 1600 1377 1634
rect 1411 1600 1467 1634
rect 1501 1600 1617 1634
rect 329 1566 1617 1600
rect 1717 2821 3005 2854
rect 1717 2787 1775 2821
rect 1809 2787 1865 2821
rect 1899 2787 1955 2821
rect 1989 2787 2045 2821
rect 2079 2787 2135 2821
rect 2169 2787 2225 2821
rect 2259 2787 2315 2821
rect 2349 2787 2405 2821
rect 2439 2787 2495 2821
rect 2529 2787 2585 2821
rect 2619 2787 2675 2821
rect 2709 2787 2765 2821
rect 2799 2787 2855 2821
rect 2889 2787 3005 2821
rect 1717 2753 3005 2787
rect 1717 2720 1818 2753
rect 1717 2686 1752 2720
rect 1786 2686 1818 2720
rect 2904 2720 3005 2753
rect 1717 2630 1818 2686
rect 1717 2596 1752 2630
rect 1786 2596 1818 2630
rect 1717 2540 1818 2596
rect 1717 2506 1752 2540
rect 1786 2506 1818 2540
rect 1717 2450 1818 2506
rect 1717 2416 1752 2450
rect 1786 2416 1818 2450
rect 1717 2360 1818 2416
rect 1717 2326 1752 2360
rect 1786 2326 1818 2360
rect 1717 2270 1818 2326
rect 1717 2236 1752 2270
rect 1786 2236 1818 2270
rect 1717 2180 1818 2236
rect 1717 2146 1752 2180
rect 1786 2146 1818 2180
rect 1717 2090 1818 2146
rect 1717 2056 1752 2090
rect 1786 2056 1818 2090
rect 1717 2000 1818 2056
rect 1717 1966 1752 2000
rect 1786 1966 1818 2000
rect 1717 1910 1818 1966
rect 1717 1876 1752 1910
rect 1786 1876 1818 1910
rect 1717 1820 1818 1876
rect 1717 1786 1752 1820
rect 1786 1786 1818 1820
rect 1717 1730 1818 1786
rect 1717 1696 1752 1730
rect 1786 1696 1818 1730
rect 2904 2686 2939 2720
rect 2973 2686 3005 2720
rect 2904 2630 3005 2686
rect 2904 2596 2939 2630
rect 2973 2596 3005 2630
rect 2904 2540 3005 2596
rect 2904 2506 2939 2540
rect 2973 2506 3005 2540
rect 2904 2450 3005 2506
rect 2904 2416 2939 2450
rect 2973 2416 3005 2450
rect 2904 2360 3005 2416
rect 2904 2326 2939 2360
rect 2973 2326 3005 2360
rect 2904 2270 3005 2326
rect 2904 2236 2939 2270
rect 2973 2236 3005 2270
rect 2904 2180 3005 2236
rect 2904 2146 2939 2180
rect 2973 2146 3005 2180
rect 2904 2090 3005 2146
rect 2904 2056 2939 2090
rect 2973 2056 3005 2090
rect 2904 2000 3005 2056
rect 2904 1966 2939 2000
rect 2973 1966 3005 2000
rect 2904 1910 3005 1966
rect 2904 1876 2939 1910
rect 2973 1876 3005 1910
rect 2904 1820 3005 1876
rect 2904 1786 2939 1820
rect 2973 1786 3005 1820
rect 2904 1730 3005 1786
rect 1717 1667 1818 1696
rect 2904 1696 2939 1730
rect 2973 1696 3005 1730
rect 2904 1667 3005 1696
rect 1717 1634 3005 1667
rect 1717 1600 1775 1634
rect 1809 1600 1865 1634
rect 1899 1600 1955 1634
rect 1989 1600 2045 1634
rect 2079 1600 2135 1634
rect 2169 1600 2225 1634
rect 2259 1600 2315 1634
rect 2349 1600 2405 1634
rect 2439 1600 2495 1634
rect 2529 1600 2585 1634
rect 2619 1600 2675 1634
rect 2709 1600 2765 1634
rect 2799 1600 2855 1634
rect 2889 1600 3005 1634
rect 1717 1566 3005 1600
rect 3105 2821 4393 2854
rect 3105 2787 3163 2821
rect 3197 2787 3253 2821
rect 3287 2787 3343 2821
rect 3377 2787 3433 2821
rect 3467 2787 3523 2821
rect 3557 2787 3613 2821
rect 3647 2787 3703 2821
rect 3737 2787 3793 2821
rect 3827 2787 3883 2821
rect 3917 2787 3973 2821
rect 4007 2787 4063 2821
rect 4097 2787 4153 2821
rect 4187 2787 4243 2821
rect 4277 2787 4393 2821
rect 3105 2753 4393 2787
rect 3105 2720 3206 2753
rect 3105 2686 3140 2720
rect 3174 2686 3206 2720
rect 4292 2720 4393 2753
rect 3105 2630 3206 2686
rect 3105 2596 3140 2630
rect 3174 2596 3206 2630
rect 3105 2540 3206 2596
rect 3105 2506 3140 2540
rect 3174 2506 3206 2540
rect 3105 2450 3206 2506
rect 3105 2416 3140 2450
rect 3174 2416 3206 2450
rect 3105 2360 3206 2416
rect 3105 2326 3140 2360
rect 3174 2326 3206 2360
rect 3105 2270 3206 2326
rect 3105 2236 3140 2270
rect 3174 2236 3206 2270
rect 3105 2180 3206 2236
rect 3105 2146 3140 2180
rect 3174 2146 3206 2180
rect 3105 2090 3206 2146
rect 3105 2056 3140 2090
rect 3174 2056 3206 2090
rect 3105 2000 3206 2056
rect 3105 1966 3140 2000
rect 3174 1966 3206 2000
rect 3105 1910 3206 1966
rect 3105 1876 3140 1910
rect 3174 1876 3206 1910
rect 3105 1820 3206 1876
rect 3105 1786 3140 1820
rect 3174 1786 3206 1820
rect 3105 1730 3206 1786
rect 3105 1696 3140 1730
rect 3174 1696 3206 1730
rect 4292 2686 4327 2720
rect 4361 2686 4393 2720
rect 4292 2630 4393 2686
rect 4292 2596 4327 2630
rect 4361 2596 4393 2630
rect 4292 2540 4393 2596
rect 4292 2506 4327 2540
rect 4361 2506 4393 2540
rect 4292 2450 4393 2506
rect 4292 2416 4327 2450
rect 4361 2416 4393 2450
rect 4292 2360 4393 2416
rect 4292 2326 4327 2360
rect 4361 2326 4393 2360
rect 4292 2270 4393 2326
rect 4292 2236 4327 2270
rect 4361 2236 4393 2270
rect 4292 2180 4393 2236
rect 4292 2146 4327 2180
rect 4361 2146 4393 2180
rect 4292 2090 4393 2146
rect 4292 2056 4327 2090
rect 4361 2056 4393 2090
rect 4292 2000 4393 2056
rect 4292 1966 4327 2000
rect 4361 1966 4393 2000
rect 4292 1910 4393 1966
rect 4292 1876 4327 1910
rect 4361 1876 4393 1910
rect 4292 1820 4393 1876
rect 4292 1786 4327 1820
rect 4361 1786 4393 1820
rect 4292 1730 4393 1786
rect 3105 1667 3206 1696
rect 4292 1696 4327 1730
rect 4361 1696 4393 1730
rect 4292 1667 4393 1696
rect 3105 1634 4393 1667
rect 3105 1600 3163 1634
rect 3197 1600 3253 1634
rect 3287 1600 3343 1634
rect 3377 1600 3433 1634
rect 3467 1600 3523 1634
rect 3557 1600 3613 1634
rect 3647 1600 3703 1634
rect 3737 1600 3793 1634
rect 3827 1600 3883 1634
rect 3917 1600 3973 1634
rect 4007 1600 4063 1634
rect 4097 1600 4153 1634
rect 4187 1600 4243 1634
rect 4277 1600 4393 1634
rect 3105 1566 4393 1600
rect 4493 2821 5781 2854
rect 4493 2787 4551 2821
rect 4585 2787 4641 2821
rect 4675 2787 4731 2821
rect 4765 2787 4821 2821
rect 4855 2787 4911 2821
rect 4945 2787 5001 2821
rect 5035 2787 5091 2821
rect 5125 2787 5181 2821
rect 5215 2787 5271 2821
rect 5305 2787 5361 2821
rect 5395 2787 5451 2821
rect 5485 2787 5541 2821
rect 5575 2787 5631 2821
rect 5665 2787 5781 2821
rect 4493 2753 5781 2787
rect 4493 2720 4594 2753
rect 4493 2686 4528 2720
rect 4562 2686 4594 2720
rect 5680 2720 5781 2753
rect 4493 2630 4594 2686
rect 4493 2596 4528 2630
rect 4562 2596 4594 2630
rect 4493 2540 4594 2596
rect 4493 2506 4528 2540
rect 4562 2506 4594 2540
rect 4493 2450 4594 2506
rect 4493 2416 4528 2450
rect 4562 2416 4594 2450
rect 4493 2360 4594 2416
rect 4493 2326 4528 2360
rect 4562 2326 4594 2360
rect 4493 2270 4594 2326
rect 4493 2236 4528 2270
rect 4562 2236 4594 2270
rect 4493 2180 4594 2236
rect 4493 2146 4528 2180
rect 4562 2146 4594 2180
rect 4493 2090 4594 2146
rect 4493 2056 4528 2090
rect 4562 2056 4594 2090
rect 4493 2000 4594 2056
rect 4493 1966 4528 2000
rect 4562 1966 4594 2000
rect 4493 1910 4594 1966
rect 4493 1876 4528 1910
rect 4562 1876 4594 1910
rect 4493 1820 4594 1876
rect 4493 1786 4528 1820
rect 4562 1786 4594 1820
rect 4493 1730 4594 1786
rect 4493 1696 4528 1730
rect 4562 1696 4594 1730
rect 5680 2686 5715 2720
rect 5749 2686 5781 2720
rect 5680 2630 5781 2686
rect 5680 2596 5715 2630
rect 5749 2596 5781 2630
rect 5680 2540 5781 2596
rect 5680 2506 5715 2540
rect 5749 2506 5781 2540
rect 5680 2450 5781 2506
rect 5680 2416 5715 2450
rect 5749 2416 5781 2450
rect 5680 2360 5781 2416
rect 5680 2326 5715 2360
rect 5749 2326 5781 2360
rect 5680 2270 5781 2326
rect 5680 2236 5715 2270
rect 5749 2236 5781 2270
rect 5680 2180 5781 2236
rect 5680 2146 5715 2180
rect 5749 2146 5781 2180
rect 5680 2090 5781 2146
rect 5680 2056 5715 2090
rect 5749 2056 5781 2090
rect 5680 2000 5781 2056
rect 5680 1966 5715 2000
rect 5749 1966 5781 2000
rect 5680 1910 5781 1966
rect 5680 1876 5715 1910
rect 5749 1876 5781 1910
rect 5680 1820 5781 1876
rect 5680 1786 5715 1820
rect 5749 1786 5781 1820
rect 5680 1730 5781 1786
rect 4493 1667 4594 1696
rect 5680 1696 5715 1730
rect 5749 1696 5781 1730
rect 5680 1667 5781 1696
rect 4493 1634 5781 1667
rect 4493 1600 4551 1634
rect 4585 1600 4641 1634
rect 4675 1600 4731 1634
rect 4765 1600 4821 1634
rect 4855 1600 4911 1634
rect 4945 1600 5001 1634
rect 5035 1600 5091 1634
rect 5125 1600 5181 1634
rect 5215 1600 5271 1634
rect 5305 1600 5361 1634
rect 5395 1600 5451 1634
rect 5485 1600 5541 1634
rect 5575 1600 5631 1634
rect 5665 1600 5781 1634
rect 4493 1566 5781 1600
rect 5881 2821 7169 2854
rect 5881 2787 5939 2821
rect 5973 2787 6029 2821
rect 6063 2787 6119 2821
rect 6153 2787 6209 2821
rect 6243 2787 6299 2821
rect 6333 2787 6389 2821
rect 6423 2787 6479 2821
rect 6513 2787 6569 2821
rect 6603 2787 6659 2821
rect 6693 2787 6749 2821
rect 6783 2787 6839 2821
rect 6873 2787 6929 2821
rect 6963 2787 7019 2821
rect 7053 2787 7169 2821
rect 5881 2753 7169 2787
rect 5881 2720 5982 2753
rect 5881 2686 5916 2720
rect 5950 2686 5982 2720
rect 7068 2720 7169 2753
rect 5881 2630 5982 2686
rect 5881 2596 5916 2630
rect 5950 2596 5982 2630
rect 5881 2540 5982 2596
rect 5881 2506 5916 2540
rect 5950 2506 5982 2540
rect 5881 2450 5982 2506
rect 5881 2416 5916 2450
rect 5950 2416 5982 2450
rect 5881 2360 5982 2416
rect 5881 2326 5916 2360
rect 5950 2326 5982 2360
rect 5881 2270 5982 2326
rect 5881 2236 5916 2270
rect 5950 2236 5982 2270
rect 5881 2180 5982 2236
rect 5881 2146 5916 2180
rect 5950 2146 5982 2180
rect 5881 2090 5982 2146
rect 5881 2056 5916 2090
rect 5950 2056 5982 2090
rect 5881 2000 5982 2056
rect 5881 1966 5916 2000
rect 5950 1966 5982 2000
rect 5881 1910 5982 1966
rect 5881 1876 5916 1910
rect 5950 1876 5982 1910
rect 5881 1820 5982 1876
rect 5881 1786 5916 1820
rect 5950 1786 5982 1820
rect 5881 1730 5982 1786
rect 5881 1696 5916 1730
rect 5950 1696 5982 1730
rect 7068 2686 7103 2720
rect 7137 2686 7169 2720
rect 7068 2630 7169 2686
rect 7068 2596 7103 2630
rect 7137 2596 7169 2630
rect 7068 2540 7169 2596
rect 7068 2506 7103 2540
rect 7137 2506 7169 2540
rect 7068 2450 7169 2506
rect 7068 2416 7103 2450
rect 7137 2416 7169 2450
rect 7068 2360 7169 2416
rect 7068 2326 7103 2360
rect 7137 2326 7169 2360
rect 7068 2270 7169 2326
rect 7068 2236 7103 2270
rect 7137 2236 7169 2270
rect 7068 2180 7169 2236
rect 7068 2146 7103 2180
rect 7137 2146 7169 2180
rect 7068 2090 7169 2146
rect 7068 2056 7103 2090
rect 7137 2056 7169 2090
rect 7068 2000 7169 2056
rect 7068 1966 7103 2000
rect 7137 1966 7169 2000
rect 7068 1910 7169 1966
rect 7068 1876 7103 1910
rect 7137 1876 7169 1910
rect 7068 1820 7169 1876
rect 7068 1786 7103 1820
rect 7137 1786 7169 1820
rect 7068 1730 7169 1786
rect 5881 1667 5982 1696
rect 7068 1696 7103 1730
rect 7137 1696 7169 1730
rect 7068 1667 7169 1696
rect 5881 1634 7169 1667
rect 5881 1600 5939 1634
rect 5973 1600 6029 1634
rect 6063 1600 6119 1634
rect 6153 1600 6209 1634
rect 6243 1600 6299 1634
rect 6333 1600 6389 1634
rect 6423 1600 6479 1634
rect 6513 1600 6569 1634
rect 6603 1600 6659 1634
rect 6693 1600 6749 1634
rect 6783 1600 6839 1634
rect 6873 1600 6929 1634
rect 6963 1600 7019 1634
rect 7053 1600 7169 1634
rect 5881 1566 7169 1600
<< nsubdiff >>
rect -17957 23001 9221 23021
rect -17957 22967 -17877 23001
rect 9141 22967 9221 23001
rect -17957 22947 9221 22967
rect -17957 22941 -17883 22947
rect -17957 -375 -17937 22941
rect -17903 -375 -17883 22941
rect 9147 22941 9221 22947
rect -16699 17607 -16606 17641
rect -7986 17607 -7901 17641
rect -16699 17581 -16665 17607
rect -7935 17581 -7901 17607
rect -16699 15698 -16665 15724
rect -7935 15698 -7901 15724
rect -16699 15664 -16606 15698
rect -7986 15664 -7901 15698
rect -7670 17518 -7585 17552
rect -3081 17518 -2996 17552
rect -7670 17492 -7636 17518
rect -3030 17492 -2996 17518
rect -7670 15692 -7636 15718
rect -3030 15692 -2996 15718
rect -7670 15658 -7585 15692
rect -3081 15658 -2996 15692
rect -12483 15558 -12423 15592
rect -7986 15558 -7926 15592
rect -12483 15532 -12449 15558
rect -7960 15532 -7926 15558
rect -12483 14696 -12449 14722
rect -7562 15543 -7502 15577
rect -3096 15543 -3036 15577
rect -7562 15517 -7528 15543
rect -3070 15517 -3036 15543
rect -7562 14759 -7528 14785
rect -3070 14759 -3036 14785
rect -7562 14725 -7502 14759
rect -3096 14725 -3036 14759
rect -7960 14696 -7926 14722
rect -12483 14662 -12423 14696
rect -7986 14662 -7926 14696
rect 287 12589 6421 12609
rect 287 12555 367 12589
rect 6341 12555 6421 12589
rect 287 12535 6421 12555
rect 287 12529 361 12535
rect 287 10033 307 12529
rect 341 10033 361 12529
rect 6347 12529 6421 12535
rect 4836 11878 4896 11912
rect 6076 11878 6136 11912
rect 4836 11852 4870 11878
rect 6102 11852 6136 11878
rect 4836 10620 4870 10646
rect 6102 10620 6136 10646
rect 4836 10586 4896 10620
rect 6076 10586 6136 10620
rect 287 10027 361 10033
rect 6347 10033 6367 12529
rect 6401 10033 6421 12529
rect 6347 10027 6421 10033
rect 287 10007 6421 10027
rect 287 9973 367 10007
rect 6341 9973 6421 10007
rect 287 9953 6421 9973
rect 492 8224 1454 8243
rect 492 8190 587 8224
rect 621 8190 677 8224
rect 711 8190 767 8224
rect 801 8190 857 8224
rect 891 8190 947 8224
rect 981 8190 1037 8224
rect 1071 8190 1127 8224
rect 1161 8190 1217 8224
rect 1251 8190 1307 8224
rect 1341 8190 1454 8224
rect 492 8171 1454 8190
rect 492 8166 564 8171
rect 492 8132 511 8166
rect 545 8132 564 8166
rect 492 8076 564 8132
rect 1382 8132 1454 8171
rect 492 8042 511 8076
rect 545 8042 564 8076
rect 492 7986 564 8042
rect 492 7952 511 7986
rect 545 7952 564 7986
rect 492 7896 564 7952
rect 492 7862 511 7896
rect 545 7862 564 7896
rect 492 7806 564 7862
rect 492 7772 511 7806
rect 545 7772 564 7806
rect 492 7716 564 7772
rect 492 7682 511 7716
rect 545 7682 564 7716
rect 492 7626 564 7682
rect 492 7592 511 7626
rect 545 7592 564 7626
rect 492 7536 564 7592
rect 492 7502 511 7536
rect 545 7502 564 7536
rect 492 7446 564 7502
rect 492 7412 511 7446
rect 545 7412 564 7446
rect 1382 8098 1401 8132
rect 1435 8098 1454 8132
rect 1382 8042 1454 8098
rect 1382 8008 1401 8042
rect 1435 8008 1454 8042
rect 1382 7952 1454 8008
rect 1382 7918 1401 7952
rect 1435 7918 1454 7952
rect 1382 7862 1454 7918
rect 1382 7828 1401 7862
rect 1435 7828 1454 7862
rect 1382 7772 1454 7828
rect 1382 7738 1401 7772
rect 1435 7738 1454 7772
rect 1382 7682 1454 7738
rect 1382 7648 1401 7682
rect 1435 7648 1454 7682
rect 1382 7592 1454 7648
rect 1382 7558 1401 7592
rect 1435 7558 1454 7592
rect 1382 7502 1454 7558
rect 1382 7468 1401 7502
rect 1435 7468 1454 7502
rect 492 7353 564 7412
rect 1382 7412 1454 7468
rect 1382 7378 1401 7412
rect 1435 7378 1454 7412
rect 1382 7353 1454 7378
rect 492 7334 1454 7353
rect 492 7300 568 7334
rect 602 7300 658 7334
rect 692 7300 748 7334
rect 782 7300 838 7334
rect 872 7300 928 7334
rect 962 7300 1018 7334
rect 1052 7300 1108 7334
rect 1142 7300 1198 7334
rect 1232 7300 1288 7334
rect 1322 7300 1454 7334
rect 492 7281 1454 7300
rect 1880 8224 2842 8243
rect 1880 8190 1975 8224
rect 2009 8190 2065 8224
rect 2099 8190 2155 8224
rect 2189 8190 2245 8224
rect 2279 8190 2335 8224
rect 2369 8190 2425 8224
rect 2459 8190 2515 8224
rect 2549 8190 2605 8224
rect 2639 8190 2695 8224
rect 2729 8190 2842 8224
rect 1880 8171 2842 8190
rect 1880 8166 1952 8171
rect 1880 8132 1899 8166
rect 1933 8132 1952 8166
rect 1880 8076 1952 8132
rect 2770 8132 2842 8171
rect 1880 8042 1899 8076
rect 1933 8042 1952 8076
rect 1880 7986 1952 8042
rect 1880 7952 1899 7986
rect 1933 7952 1952 7986
rect 1880 7896 1952 7952
rect 1880 7862 1899 7896
rect 1933 7862 1952 7896
rect 1880 7806 1952 7862
rect 1880 7772 1899 7806
rect 1933 7772 1952 7806
rect 1880 7716 1952 7772
rect 1880 7682 1899 7716
rect 1933 7682 1952 7716
rect 1880 7626 1952 7682
rect 1880 7592 1899 7626
rect 1933 7592 1952 7626
rect 1880 7536 1952 7592
rect 1880 7502 1899 7536
rect 1933 7502 1952 7536
rect 1880 7446 1952 7502
rect 1880 7412 1899 7446
rect 1933 7412 1952 7446
rect 2770 8098 2789 8132
rect 2823 8098 2842 8132
rect 2770 8042 2842 8098
rect 2770 8008 2789 8042
rect 2823 8008 2842 8042
rect 2770 7952 2842 8008
rect 2770 7918 2789 7952
rect 2823 7918 2842 7952
rect 2770 7862 2842 7918
rect 2770 7828 2789 7862
rect 2823 7828 2842 7862
rect 2770 7772 2842 7828
rect 2770 7738 2789 7772
rect 2823 7738 2842 7772
rect 2770 7682 2842 7738
rect 2770 7648 2789 7682
rect 2823 7648 2842 7682
rect 2770 7592 2842 7648
rect 2770 7558 2789 7592
rect 2823 7558 2842 7592
rect 2770 7502 2842 7558
rect 2770 7468 2789 7502
rect 2823 7468 2842 7502
rect 1880 7353 1952 7412
rect 2770 7412 2842 7468
rect 2770 7378 2789 7412
rect 2823 7378 2842 7412
rect 2770 7353 2842 7378
rect 1880 7334 2842 7353
rect 1880 7300 1956 7334
rect 1990 7300 2046 7334
rect 2080 7300 2136 7334
rect 2170 7300 2226 7334
rect 2260 7300 2316 7334
rect 2350 7300 2406 7334
rect 2440 7300 2496 7334
rect 2530 7300 2586 7334
rect 2620 7300 2676 7334
rect 2710 7300 2842 7334
rect 1880 7281 2842 7300
rect 3268 8224 4230 8243
rect 3268 8190 3363 8224
rect 3397 8190 3453 8224
rect 3487 8190 3543 8224
rect 3577 8190 3633 8224
rect 3667 8190 3723 8224
rect 3757 8190 3813 8224
rect 3847 8190 3903 8224
rect 3937 8190 3993 8224
rect 4027 8190 4083 8224
rect 4117 8190 4230 8224
rect 3268 8171 4230 8190
rect 3268 8166 3340 8171
rect 3268 8132 3287 8166
rect 3321 8132 3340 8166
rect 3268 8076 3340 8132
rect 4158 8132 4230 8171
rect 3268 8042 3287 8076
rect 3321 8042 3340 8076
rect 3268 7986 3340 8042
rect 3268 7952 3287 7986
rect 3321 7952 3340 7986
rect 3268 7896 3340 7952
rect 3268 7862 3287 7896
rect 3321 7862 3340 7896
rect 3268 7806 3340 7862
rect 3268 7772 3287 7806
rect 3321 7772 3340 7806
rect 3268 7716 3340 7772
rect 3268 7682 3287 7716
rect 3321 7682 3340 7716
rect 3268 7626 3340 7682
rect 3268 7592 3287 7626
rect 3321 7592 3340 7626
rect 3268 7536 3340 7592
rect 3268 7502 3287 7536
rect 3321 7502 3340 7536
rect 3268 7446 3340 7502
rect 3268 7412 3287 7446
rect 3321 7412 3340 7446
rect 4158 8098 4177 8132
rect 4211 8098 4230 8132
rect 4158 8042 4230 8098
rect 4158 8008 4177 8042
rect 4211 8008 4230 8042
rect 4158 7952 4230 8008
rect 4158 7918 4177 7952
rect 4211 7918 4230 7952
rect 4158 7862 4230 7918
rect 4158 7828 4177 7862
rect 4211 7828 4230 7862
rect 4158 7772 4230 7828
rect 4158 7738 4177 7772
rect 4211 7738 4230 7772
rect 4158 7682 4230 7738
rect 4158 7648 4177 7682
rect 4211 7648 4230 7682
rect 4158 7592 4230 7648
rect 4158 7558 4177 7592
rect 4211 7558 4230 7592
rect 4158 7502 4230 7558
rect 4158 7468 4177 7502
rect 4211 7468 4230 7502
rect 3268 7353 3340 7412
rect 4158 7412 4230 7468
rect 4158 7378 4177 7412
rect 4211 7378 4230 7412
rect 4158 7353 4230 7378
rect 3268 7334 4230 7353
rect 3268 7300 3344 7334
rect 3378 7300 3434 7334
rect 3468 7300 3524 7334
rect 3558 7300 3614 7334
rect 3648 7300 3704 7334
rect 3738 7300 3794 7334
rect 3828 7300 3884 7334
rect 3918 7300 3974 7334
rect 4008 7300 4064 7334
rect 4098 7300 4230 7334
rect 3268 7281 4230 7300
rect 4656 8224 5618 8243
rect 4656 8190 4751 8224
rect 4785 8190 4841 8224
rect 4875 8190 4931 8224
rect 4965 8190 5021 8224
rect 5055 8190 5111 8224
rect 5145 8190 5201 8224
rect 5235 8190 5291 8224
rect 5325 8190 5381 8224
rect 5415 8190 5471 8224
rect 5505 8190 5618 8224
rect 4656 8171 5618 8190
rect 4656 8166 4728 8171
rect 4656 8132 4675 8166
rect 4709 8132 4728 8166
rect 4656 8076 4728 8132
rect 5546 8132 5618 8171
rect 4656 8042 4675 8076
rect 4709 8042 4728 8076
rect 4656 7986 4728 8042
rect 4656 7952 4675 7986
rect 4709 7952 4728 7986
rect 4656 7896 4728 7952
rect 4656 7862 4675 7896
rect 4709 7862 4728 7896
rect 4656 7806 4728 7862
rect 4656 7772 4675 7806
rect 4709 7772 4728 7806
rect 4656 7716 4728 7772
rect 4656 7682 4675 7716
rect 4709 7682 4728 7716
rect 4656 7626 4728 7682
rect 4656 7592 4675 7626
rect 4709 7592 4728 7626
rect 4656 7536 4728 7592
rect 4656 7502 4675 7536
rect 4709 7502 4728 7536
rect 4656 7446 4728 7502
rect 4656 7412 4675 7446
rect 4709 7412 4728 7446
rect 5546 8098 5565 8132
rect 5599 8098 5618 8132
rect 5546 8042 5618 8098
rect 5546 8008 5565 8042
rect 5599 8008 5618 8042
rect 5546 7952 5618 8008
rect 5546 7918 5565 7952
rect 5599 7918 5618 7952
rect 5546 7862 5618 7918
rect 5546 7828 5565 7862
rect 5599 7828 5618 7862
rect 5546 7772 5618 7828
rect 5546 7738 5565 7772
rect 5599 7738 5618 7772
rect 5546 7682 5618 7738
rect 5546 7648 5565 7682
rect 5599 7648 5618 7682
rect 5546 7592 5618 7648
rect 5546 7558 5565 7592
rect 5599 7558 5618 7592
rect 5546 7502 5618 7558
rect 5546 7468 5565 7502
rect 5599 7468 5618 7502
rect 4656 7353 4728 7412
rect 5546 7412 5618 7468
rect 5546 7378 5565 7412
rect 5599 7378 5618 7412
rect 5546 7353 5618 7378
rect 4656 7334 5618 7353
rect 4656 7300 4732 7334
rect 4766 7300 4822 7334
rect 4856 7300 4912 7334
rect 4946 7300 5002 7334
rect 5036 7300 5092 7334
rect 5126 7300 5182 7334
rect 5216 7300 5272 7334
rect 5306 7300 5362 7334
rect 5396 7300 5452 7334
rect 5486 7300 5618 7334
rect 4656 7281 5618 7300
rect 6044 8224 7006 8243
rect 6044 8190 6139 8224
rect 6173 8190 6229 8224
rect 6263 8190 6319 8224
rect 6353 8190 6409 8224
rect 6443 8190 6499 8224
rect 6533 8190 6589 8224
rect 6623 8190 6679 8224
rect 6713 8190 6769 8224
rect 6803 8190 6859 8224
rect 6893 8190 7006 8224
rect 6044 8171 7006 8190
rect 6044 8166 6116 8171
rect 6044 8132 6063 8166
rect 6097 8132 6116 8166
rect 6044 8076 6116 8132
rect 6934 8132 7006 8171
rect 6044 8042 6063 8076
rect 6097 8042 6116 8076
rect 6044 7986 6116 8042
rect 6044 7952 6063 7986
rect 6097 7952 6116 7986
rect 6044 7896 6116 7952
rect 6044 7862 6063 7896
rect 6097 7862 6116 7896
rect 6044 7806 6116 7862
rect 6044 7772 6063 7806
rect 6097 7772 6116 7806
rect 6044 7716 6116 7772
rect 6044 7682 6063 7716
rect 6097 7682 6116 7716
rect 6044 7626 6116 7682
rect 6044 7592 6063 7626
rect 6097 7592 6116 7626
rect 6044 7536 6116 7592
rect 6044 7502 6063 7536
rect 6097 7502 6116 7536
rect 6044 7446 6116 7502
rect 6044 7412 6063 7446
rect 6097 7412 6116 7446
rect 6934 8098 6953 8132
rect 6987 8098 7006 8132
rect 6934 8042 7006 8098
rect 6934 8008 6953 8042
rect 6987 8008 7006 8042
rect 6934 7952 7006 8008
rect 6934 7918 6953 7952
rect 6987 7918 7006 7952
rect 6934 7862 7006 7918
rect 6934 7828 6953 7862
rect 6987 7828 7006 7862
rect 6934 7772 7006 7828
rect 6934 7738 6953 7772
rect 6987 7738 7006 7772
rect 6934 7682 7006 7738
rect 6934 7648 6953 7682
rect 6987 7648 7006 7682
rect 6934 7592 7006 7648
rect 6934 7558 6953 7592
rect 6987 7558 7006 7592
rect 6934 7502 7006 7558
rect 6934 7468 6953 7502
rect 6987 7468 7006 7502
rect 6044 7353 6116 7412
rect 6934 7412 7006 7468
rect 6934 7378 6953 7412
rect 6987 7378 7006 7412
rect 6934 7353 7006 7378
rect 6044 7334 7006 7353
rect 6044 7300 6120 7334
rect 6154 7300 6210 7334
rect 6244 7300 6300 7334
rect 6334 7300 6390 7334
rect 6424 7300 6480 7334
rect 6514 7300 6570 7334
rect 6604 7300 6660 7334
rect 6694 7300 6750 7334
rect 6784 7300 6840 7334
rect 6874 7300 7006 7334
rect 6044 7281 7006 7300
rect 492 6836 1454 6855
rect 492 6802 587 6836
rect 621 6802 677 6836
rect 711 6802 767 6836
rect 801 6802 857 6836
rect 891 6802 947 6836
rect 981 6802 1037 6836
rect 1071 6802 1127 6836
rect 1161 6802 1217 6836
rect 1251 6802 1307 6836
rect 1341 6802 1454 6836
rect 492 6783 1454 6802
rect 492 6778 564 6783
rect 492 6744 511 6778
rect 545 6744 564 6778
rect 492 6688 564 6744
rect 1382 6744 1454 6783
rect 492 6654 511 6688
rect 545 6654 564 6688
rect 492 6598 564 6654
rect 492 6564 511 6598
rect 545 6564 564 6598
rect 492 6508 564 6564
rect 492 6474 511 6508
rect 545 6474 564 6508
rect 492 6418 564 6474
rect 492 6384 511 6418
rect 545 6384 564 6418
rect 492 6328 564 6384
rect 492 6294 511 6328
rect 545 6294 564 6328
rect 492 6238 564 6294
rect 492 6204 511 6238
rect 545 6204 564 6238
rect 492 6148 564 6204
rect 492 6114 511 6148
rect 545 6114 564 6148
rect 492 6058 564 6114
rect 492 6024 511 6058
rect 545 6024 564 6058
rect 1382 6710 1401 6744
rect 1435 6710 1454 6744
rect 1382 6654 1454 6710
rect 1382 6620 1401 6654
rect 1435 6620 1454 6654
rect 1382 6564 1454 6620
rect 1382 6530 1401 6564
rect 1435 6530 1454 6564
rect 1382 6474 1454 6530
rect 1382 6440 1401 6474
rect 1435 6440 1454 6474
rect 1382 6384 1454 6440
rect 1382 6350 1401 6384
rect 1435 6350 1454 6384
rect 1382 6294 1454 6350
rect 1382 6260 1401 6294
rect 1435 6260 1454 6294
rect 1382 6204 1454 6260
rect 1382 6170 1401 6204
rect 1435 6170 1454 6204
rect 1382 6114 1454 6170
rect 1382 6080 1401 6114
rect 1435 6080 1454 6114
rect 492 5965 564 6024
rect 1382 6024 1454 6080
rect 1382 5990 1401 6024
rect 1435 5990 1454 6024
rect 1382 5965 1454 5990
rect 492 5946 1454 5965
rect 492 5912 568 5946
rect 602 5912 658 5946
rect 692 5912 748 5946
rect 782 5912 838 5946
rect 872 5912 928 5946
rect 962 5912 1018 5946
rect 1052 5912 1108 5946
rect 1142 5912 1198 5946
rect 1232 5912 1288 5946
rect 1322 5912 1454 5946
rect 492 5893 1454 5912
rect 1880 6836 2842 6855
rect 1880 6802 1975 6836
rect 2009 6802 2065 6836
rect 2099 6802 2155 6836
rect 2189 6802 2245 6836
rect 2279 6802 2335 6836
rect 2369 6802 2425 6836
rect 2459 6802 2515 6836
rect 2549 6802 2605 6836
rect 2639 6802 2695 6836
rect 2729 6802 2842 6836
rect 1880 6783 2842 6802
rect 1880 6778 1952 6783
rect 1880 6744 1899 6778
rect 1933 6744 1952 6778
rect 1880 6688 1952 6744
rect 2770 6744 2842 6783
rect 1880 6654 1899 6688
rect 1933 6654 1952 6688
rect 1880 6598 1952 6654
rect 1880 6564 1899 6598
rect 1933 6564 1952 6598
rect 1880 6508 1952 6564
rect 1880 6474 1899 6508
rect 1933 6474 1952 6508
rect 1880 6418 1952 6474
rect 1880 6384 1899 6418
rect 1933 6384 1952 6418
rect 1880 6328 1952 6384
rect 1880 6294 1899 6328
rect 1933 6294 1952 6328
rect 1880 6238 1952 6294
rect 1880 6204 1899 6238
rect 1933 6204 1952 6238
rect 1880 6148 1952 6204
rect 1880 6114 1899 6148
rect 1933 6114 1952 6148
rect 1880 6058 1952 6114
rect 1880 6024 1899 6058
rect 1933 6024 1952 6058
rect 2770 6710 2789 6744
rect 2823 6710 2842 6744
rect 2770 6654 2842 6710
rect 2770 6620 2789 6654
rect 2823 6620 2842 6654
rect 2770 6564 2842 6620
rect 2770 6530 2789 6564
rect 2823 6530 2842 6564
rect 2770 6474 2842 6530
rect 2770 6440 2789 6474
rect 2823 6440 2842 6474
rect 2770 6384 2842 6440
rect 2770 6350 2789 6384
rect 2823 6350 2842 6384
rect 2770 6294 2842 6350
rect 2770 6260 2789 6294
rect 2823 6260 2842 6294
rect 2770 6204 2842 6260
rect 2770 6170 2789 6204
rect 2823 6170 2842 6204
rect 2770 6114 2842 6170
rect 2770 6080 2789 6114
rect 2823 6080 2842 6114
rect 1880 5965 1952 6024
rect 2770 6024 2842 6080
rect 2770 5990 2789 6024
rect 2823 5990 2842 6024
rect 2770 5965 2842 5990
rect 1880 5946 2842 5965
rect 1880 5912 1956 5946
rect 1990 5912 2046 5946
rect 2080 5912 2136 5946
rect 2170 5912 2226 5946
rect 2260 5912 2316 5946
rect 2350 5912 2406 5946
rect 2440 5912 2496 5946
rect 2530 5912 2586 5946
rect 2620 5912 2676 5946
rect 2710 5912 2842 5946
rect 1880 5893 2842 5912
rect 3268 6836 4230 6855
rect 3268 6802 3363 6836
rect 3397 6802 3453 6836
rect 3487 6802 3543 6836
rect 3577 6802 3633 6836
rect 3667 6802 3723 6836
rect 3757 6802 3813 6836
rect 3847 6802 3903 6836
rect 3937 6802 3993 6836
rect 4027 6802 4083 6836
rect 4117 6802 4230 6836
rect 3268 6783 4230 6802
rect 3268 6778 3340 6783
rect 3268 6744 3287 6778
rect 3321 6744 3340 6778
rect 3268 6688 3340 6744
rect 4158 6744 4230 6783
rect 3268 6654 3287 6688
rect 3321 6654 3340 6688
rect 3268 6598 3340 6654
rect 3268 6564 3287 6598
rect 3321 6564 3340 6598
rect 3268 6508 3340 6564
rect 3268 6474 3287 6508
rect 3321 6474 3340 6508
rect 3268 6418 3340 6474
rect 3268 6384 3287 6418
rect 3321 6384 3340 6418
rect 3268 6328 3340 6384
rect 3268 6294 3287 6328
rect 3321 6294 3340 6328
rect 3268 6238 3340 6294
rect 3268 6204 3287 6238
rect 3321 6204 3340 6238
rect 3268 6148 3340 6204
rect 3268 6114 3287 6148
rect 3321 6114 3340 6148
rect 3268 6058 3340 6114
rect 3268 6024 3287 6058
rect 3321 6024 3340 6058
rect 4158 6710 4177 6744
rect 4211 6710 4230 6744
rect 4158 6654 4230 6710
rect 4158 6620 4177 6654
rect 4211 6620 4230 6654
rect 4158 6564 4230 6620
rect 4158 6530 4177 6564
rect 4211 6530 4230 6564
rect 4158 6474 4230 6530
rect 4158 6440 4177 6474
rect 4211 6440 4230 6474
rect 4158 6384 4230 6440
rect 4158 6350 4177 6384
rect 4211 6350 4230 6384
rect 4158 6294 4230 6350
rect 4158 6260 4177 6294
rect 4211 6260 4230 6294
rect 4158 6204 4230 6260
rect 4158 6170 4177 6204
rect 4211 6170 4230 6204
rect 4158 6114 4230 6170
rect 4158 6080 4177 6114
rect 4211 6080 4230 6114
rect 3268 5965 3340 6024
rect 4158 6024 4230 6080
rect 4158 5990 4177 6024
rect 4211 5990 4230 6024
rect 4158 5965 4230 5990
rect 3268 5946 4230 5965
rect 3268 5912 3344 5946
rect 3378 5912 3434 5946
rect 3468 5912 3524 5946
rect 3558 5912 3614 5946
rect 3648 5912 3704 5946
rect 3738 5912 3794 5946
rect 3828 5912 3884 5946
rect 3918 5912 3974 5946
rect 4008 5912 4064 5946
rect 4098 5912 4230 5946
rect 3268 5893 4230 5912
rect 4656 6836 5618 6855
rect 4656 6802 4751 6836
rect 4785 6802 4841 6836
rect 4875 6802 4931 6836
rect 4965 6802 5021 6836
rect 5055 6802 5111 6836
rect 5145 6802 5201 6836
rect 5235 6802 5291 6836
rect 5325 6802 5381 6836
rect 5415 6802 5471 6836
rect 5505 6802 5618 6836
rect 4656 6783 5618 6802
rect 4656 6778 4728 6783
rect 4656 6744 4675 6778
rect 4709 6744 4728 6778
rect 4656 6688 4728 6744
rect 5546 6744 5618 6783
rect 4656 6654 4675 6688
rect 4709 6654 4728 6688
rect 4656 6598 4728 6654
rect 4656 6564 4675 6598
rect 4709 6564 4728 6598
rect 4656 6508 4728 6564
rect 4656 6474 4675 6508
rect 4709 6474 4728 6508
rect 4656 6418 4728 6474
rect 4656 6384 4675 6418
rect 4709 6384 4728 6418
rect 4656 6328 4728 6384
rect 4656 6294 4675 6328
rect 4709 6294 4728 6328
rect 4656 6238 4728 6294
rect 4656 6204 4675 6238
rect 4709 6204 4728 6238
rect 4656 6148 4728 6204
rect 4656 6114 4675 6148
rect 4709 6114 4728 6148
rect 4656 6058 4728 6114
rect 4656 6024 4675 6058
rect 4709 6024 4728 6058
rect 5546 6710 5565 6744
rect 5599 6710 5618 6744
rect 5546 6654 5618 6710
rect 5546 6620 5565 6654
rect 5599 6620 5618 6654
rect 5546 6564 5618 6620
rect 5546 6530 5565 6564
rect 5599 6530 5618 6564
rect 5546 6474 5618 6530
rect 5546 6440 5565 6474
rect 5599 6440 5618 6474
rect 5546 6384 5618 6440
rect 5546 6350 5565 6384
rect 5599 6350 5618 6384
rect 5546 6294 5618 6350
rect 5546 6260 5565 6294
rect 5599 6260 5618 6294
rect 5546 6204 5618 6260
rect 5546 6170 5565 6204
rect 5599 6170 5618 6204
rect 5546 6114 5618 6170
rect 5546 6080 5565 6114
rect 5599 6080 5618 6114
rect 4656 5965 4728 6024
rect 5546 6024 5618 6080
rect 5546 5990 5565 6024
rect 5599 5990 5618 6024
rect 5546 5965 5618 5990
rect 4656 5946 5618 5965
rect 4656 5912 4732 5946
rect 4766 5912 4822 5946
rect 4856 5912 4912 5946
rect 4946 5912 5002 5946
rect 5036 5912 5092 5946
rect 5126 5912 5182 5946
rect 5216 5912 5272 5946
rect 5306 5912 5362 5946
rect 5396 5912 5452 5946
rect 5486 5912 5618 5946
rect 4656 5893 5618 5912
rect 6044 6836 7006 6855
rect 6044 6802 6139 6836
rect 6173 6802 6229 6836
rect 6263 6802 6319 6836
rect 6353 6802 6409 6836
rect 6443 6802 6499 6836
rect 6533 6802 6589 6836
rect 6623 6802 6679 6836
rect 6713 6802 6769 6836
rect 6803 6802 6859 6836
rect 6893 6802 7006 6836
rect 6044 6783 7006 6802
rect 6044 6778 6116 6783
rect 6044 6744 6063 6778
rect 6097 6744 6116 6778
rect 6044 6688 6116 6744
rect 6934 6744 7006 6783
rect 6044 6654 6063 6688
rect 6097 6654 6116 6688
rect 6044 6598 6116 6654
rect 6044 6564 6063 6598
rect 6097 6564 6116 6598
rect 6044 6508 6116 6564
rect 6044 6474 6063 6508
rect 6097 6474 6116 6508
rect 6044 6418 6116 6474
rect 6044 6384 6063 6418
rect 6097 6384 6116 6418
rect 6044 6328 6116 6384
rect 6044 6294 6063 6328
rect 6097 6294 6116 6328
rect 6044 6238 6116 6294
rect 6044 6204 6063 6238
rect 6097 6204 6116 6238
rect 6044 6148 6116 6204
rect 6044 6114 6063 6148
rect 6097 6114 6116 6148
rect 6044 6058 6116 6114
rect 6044 6024 6063 6058
rect 6097 6024 6116 6058
rect 6934 6710 6953 6744
rect 6987 6710 7006 6744
rect 6934 6654 7006 6710
rect 6934 6620 6953 6654
rect 6987 6620 7006 6654
rect 6934 6564 7006 6620
rect 6934 6530 6953 6564
rect 6987 6530 7006 6564
rect 6934 6474 7006 6530
rect 6934 6440 6953 6474
rect 6987 6440 7006 6474
rect 6934 6384 7006 6440
rect 6934 6350 6953 6384
rect 6987 6350 7006 6384
rect 6934 6294 7006 6350
rect 6934 6260 6953 6294
rect 6987 6260 7006 6294
rect 6934 6204 7006 6260
rect 6934 6170 6953 6204
rect 6987 6170 7006 6204
rect 6934 6114 7006 6170
rect 6934 6080 6953 6114
rect 6987 6080 7006 6114
rect 6044 5965 6116 6024
rect 6934 6024 7006 6080
rect 6934 5990 6953 6024
rect 6987 5990 7006 6024
rect 6934 5965 7006 5990
rect 6044 5946 7006 5965
rect 6044 5912 6120 5946
rect 6154 5912 6210 5946
rect 6244 5912 6300 5946
rect 6334 5912 6390 5946
rect 6424 5912 6480 5946
rect 6514 5912 6570 5946
rect 6604 5912 6660 5946
rect 6694 5912 6750 5946
rect 6784 5912 6840 5946
rect 6874 5912 7006 5946
rect 6044 5893 7006 5912
rect 492 5448 1454 5467
rect 492 5414 587 5448
rect 621 5414 677 5448
rect 711 5414 767 5448
rect 801 5414 857 5448
rect 891 5414 947 5448
rect 981 5414 1037 5448
rect 1071 5414 1127 5448
rect 1161 5414 1217 5448
rect 1251 5414 1307 5448
rect 1341 5414 1454 5448
rect 492 5395 1454 5414
rect 492 5390 564 5395
rect 492 5356 511 5390
rect 545 5356 564 5390
rect 492 5300 564 5356
rect 1382 5356 1454 5395
rect 492 5266 511 5300
rect 545 5266 564 5300
rect 492 5210 564 5266
rect 492 5176 511 5210
rect 545 5176 564 5210
rect 492 5120 564 5176
rect 492 5086 511 5120
rect 545 5086 564 5120
rect 492 5030 564 5086
rect 492 4996 511 5030
rect 545 4996 564 5030
rect 492 4940 564 4996
rect 492 4906 511 4940
rect 545 4906 564 4940
rect 492 4850 564 4906
rect 492 4816 511 4850
rect 545 4816 564 4850
rect 492 4760 564 4816
rect 492 4726 511 4760
rect 545 4726 564 4760
rect 492 4670 564 4726
rect 492 4636 511 4670
rect 545 4636 564 4670
rect 1382 5322 1401 5356
rect 1435 5322 1454 5356
rect 1382 5266 1454 5322
rect 1382 5232 1401 5266
rect 1435 5232 1454 5266
rect 1382 5176 1454 5232
rect 1382 5142 1401 5176
rect 1435 5142 1454 5176
rect 1382 5086 1454 5142
rect 1382 5052 1401 5086
rect 1435 5052 1454 5086
rect 1382 4996 1454 5052
rect 1382 4962 1401 4996
rect 1435 4962 1454 4996
rect 1382 4906 1454 4962
rect 1382 4872 1401 4906
rect 1435 4872 1454 4906
rect 1382 4816 1454 4872
rect 1382 4782 1401 4816
rect 1435 4782 1454 4816
rect 1382 4726 1454 4782
rect 1382 4692 1401 4726
rect 1435 4692 1454 4726
rect 492 4577 564 4636
rect 1382 4636 1454 4692
rect 1382 4602 1401 4636
rect 1435 4602 1454 4636
rect 1382 4577 1454 4602
rect 492 4558 1454 4577
rect 492 4524 568 4558
rect 602 4524 658 4558
rect 692 4524 748 4558
rect 782 4524 838 4558
rect 872 4524 928 4558
rect 962 4524 1018 4558
rect 1052 4524 1108 4558
rect 1142 4524 1198 4558
rect 1232 4524 1288 4558
rect 1322 4524 1454 4558
rect 492 4505 1454 4524
rect 1880 5448 2842 5467
rect 1880 5414 1975 5448
rect 2009 5414 2065 5448
rect 2099 5414 2155 5448
rect 2189 5414 2245 5448
rect 2279 5414 2335 5448
rect 2369 5414 2425 5448
rect 2459 5414 2515 5448
rect 2549 5414 2605 5448
rect 2639 5414 2695 5448
rect 2729 5414 2842 5448
rect 1880 5395 2842 5414
rect 1880 5390 1952 5395
rect 1880 5356 1899 5390
rect 1933 5356 1952 5390
rect 1880 5300 1952 5356
rect 2770 5356 2842 5395
rect 1880 5266 1899 5300
rect 1933 5266 1952 5300
rect 1880 5210 1952 5266
rect 1880 5176 1899 5210
rect 1933 5176 1952 5210
rect 1880 5120 1952 5176
rect 1880 5086 1899 5120
rect 1933 5086 1952 5120
rect 1880 5030 1952 5086
rect 1880 4996 1899 5030
rect 1933 4996 1952 5030
rect 1880 4940 1952 4996
rect 1880 4906 1899 4940
rect 1933 4906 1952 4940
rect 1880 4850 1952 4906
rect 1880 4816 1899 4850
rect 1933 4816 1952 4850
rect 1880 4760 1952 4816
rect 1880 4726 1899 4760
rect 1933 4726 1952 4760
rect 1880 4670 1952 4726
rect 1880 4636 1899 4670
rect 1933 4636 1952 4670
rect 2770 5322 2789 5356
rect 2823 5322 2842 5356
rect 2770 5266 2842 5322
rect 2770 5232 2789 5266
rect 2823 5232 2842 5266
rect 2770 5176 2842 5232
rect 2770 5142 2789 5176
rect 2823 5142 2842 5176
rect 2770 5086 2842 5142
rect 2770 5052 2789 5086
rect 2823 5052 2842 5086
rect 2770 4996 2842 5052
rect 2770 4962 2789 4996
rect 2823 4962 2842 4996
rect 2770 4906 2842 4962
rect 2770 4872 2789 4906
rect 2823 4872 2842 4906
rect 2770 4816 2842 4872
rect 2770 4782 2789 4816
rect 2823 4782 2842 4816
rect 2770 4726 2842 4782
rect 2770 4692 2789 4726
rect 2823 4692 2842 4726
rect 1880 4577 1952 4636
rect 2770 4636 2842 4692
rect 2770 4602 2789 4636
rect 2823 4602 2842 4636
rect 2770 4577 2842 4602
rect 1880 4558 2842 4577
rect 1880 4524 1956 4558
rect 1990 4524 2046 4558
rect 2080 4524 2136 4558
rect 2170 4524 2226 4558
rect 2260 4524 2316 4558
rect 2350 4524 2406 4558
rect 2440 4524 2496 4558
rect 2530 4524 2586 4558
rect 2620 4524 2676 4558
rect 2710 4524 2842 4558
rect 1880 4505 2842 4524
rect 3268 5448 4230 5467
rect 3268 5414 3363 5448
rect 3397 5414 3453 5448
rect 3487 5414 3543 5448
rect 3577 5414 3633 5448
rect 3667 5414 3723 5448
rect 3757 5414 3813 5448
rect 3847 5414 3903 5448
rect 3937 5414 3993 5448
rect 4027 5414 4083 5448
rect 4117 5414 4230 5448
rect 3268 5395 4230 5414
rect 3268 5390 3340 5395
rect 3268 5356 3287 5390
rect 3321 5356 3340 5390
rect 3268 5300 3340 5356
rect 4158 5356 4230 5395
rect 3268 5266 3287 5300
rect 3321 5266 3340 5300
rect 3268 5210 3340 5266
rect 3268 5176 3287 5210
rect 3321 5176 3340 5210
rect 3268 5120 3340 5176
rect 3268 5086 3287 5120
rect 3321 5086 3340 5120
rect 3268 5030 3340 5086
rect 3268 4996 3287 5030
rect 3321 4996 3340 5030
rect 3268 4940 3340 4996
rect 3268 4906 3287 4940
rect 3321 4906 3340 4940
rect 3268 4850 3340 4906
rect 3268 4816 3287 4850
rect 3321 4816 3340 4850
rect 3268 4760 3340 4816
rect 3268 4726 3287 4760
rect 3321 4726 3340 4760
rect 3268 4670 3340 4726
rect 3268 4636 3287 4670
rect 3321 4636 3340 4670
rect 4158 5322 4177 5356
rect 4211 5322 4230 5356
rect 4158 5266 4230 5322
rect 4158 5232 4177 5266
rect 4211 5232 4230 5266
rect 4158 5176 4230 5232
rect 4158 5142 4177 5176
rect 4211 5142 4230 5176
rect 4158 5086 4230 5142
rect 4158 5052 4177 5086
rect 4211 5052 4230 5086
rect 4158 4996 4230 5052
rect 4158 4962 4177 4996
rect 4211 4962 4230 4996
rect 4158 4906 4230 4962
rect 4158 4872 4177 4906
rect 4211 4872 4230 4906
rect 4158 4816 4230 4872
rect 4158 4782 4177 4816
rect 4211 4782 4230 4816
rect 4158 4726 4230 4782
rect 4158 4692 4177 4726
rect 4211 4692 4230 4726
rect 3268 4577 3340 4636
rect 4158 4636 4230 4692
rect 4158 4602 4177 4636
rect 4211 4602 4230 4636
rect 4158 4577 4230 4602
rect 3268 4558 4230 4577
rect 3268 4524 3344 4558
rect 3378 4524 3434 4558
rect 3468 4524 3524 4558
rect 3558 4524 3614 4558
rect 3648 4524 3704 4558
rect 3738 4524 3794 4558
rect 3828 4524 3884 4558
rect 3918 4524 3974 4558
rect 4008 4524 4064 4558
rect 4098 4524 4230 4558
rect 3268 4505 4230 4524
rect 4656 5448 5618 5467
rect 4656 5414 4751 5448
rect 4785 5414 4841 5448
rect 4875 5414 4931 5448
rect 4965 5414 5021 5448
rect 5055 5414 5111 5448
rect 5145 5414 5201 5448
rect 5235 5414 5291 5448
rect 5325 5414 5381 5448
rect 5415 5414 5471 5448
rect 5505 5414 5618 5448
rect 4656 5395 5618 5414
rect 4656 5390 4728 5395
rect 4656 5356 4675 5390
rect 4709 5356 4728 5390
rect 4656 5300 4728 5356
rect 5546 5356 5618 5395
rect 4656 5266 4675 5300
rect 4709 5266 4728 5300
rect 4656 5210 4728 5266
rect 4656 5176 4675 5210
rect 4709 5176 4728 5210
rect 4656 5120 4728 5176
rect 4656 5086 4675 5120
rect 4709 5086 4728 5120
rect 4656 5030 4728 5086
rect 4656 4996 4675 5030
rect 4709 4996 4728 5030
rect 4656 4940 4728 4996
rect 4656 4906 4675 4940
rect 4709 4906 4728 4940
rect 4656 4850 4728 4906
rect 4656 4816 4675 4850
rect 4709 4816 4728 4850
rect 4656 4760 4728 4816
rect 4656 4726 4675 4760
rect 4709 4726 4728 4760
rect 4656 4670 4728 4726
rect 4656 4636 4675 4670
rect 4709 4636 4728 4670
rect 5546 5322 5565 5356
rect 5599 5322 5618 5356
rect 5546 5266 5618 5322
rect 5546 5232 5565 5266
rect 5599 5232 5618 5266
rect 5546 5176 5618 5232
rect 5546 5142 5565 5176
rect 5599 5142 5618 5176
rect 5546 5086 5618 5142
rect 5546 5052 5565 5086
rect 5599 5052 5618 5086
rect 5546 4996 5618 5052
rect 5546 4962 5565 4996
rect 5599 4962 5618 4996
rect 5546 4906 5618 4962
rect 5546 4872 5565 4906
rect 5599 4872 5618 4906
rect 5546 4816 5618 4872
rect 5546 4782 5565 4816
rect 5599 4782 5618 4816
rect 5546 4726 5618 4782
rect 5546 4692 5565 4726
rect 5599 4692 5618 4726
rect 4656 4577 4728 4636
rect 5546 4636 5618 4692
rect 5546 4602 5565 4636
rect 5599 4602 5618 4636
rect 5546 4577 5618 4602
rect 4656 4558 5618 4577
rect 4656 4524 4732 4558
rect 4766 4524 4822 4558
rect 4856 4524 4912 4558
rect 4946 4524 5002 4558
rect 5036 4524 5092 4558
rect 5126 4524 5182 4558
rect 5216 4524 5272 4558
rect 5306 4524 5362 4558
rect 5396 4524 5452 4558
rect 5486 4524 5618 4558
rect 4656 4505 5618 4524
rect 6044 5448 7006 5467
rect 6044 5414 6139 5448
rect 6173 5414 6229 5448
rect 6263 5414 6319 5448
rect 6353 5414 6409 5448
rect 6443 5414 6499 5448
rect 6533 5414 6589 5448
rect 6623 5414 6679 5448
rect 6713 5414 6769 5448
rect 6803 5414 6859 5448
rect 6893 5414 7006 5448
rect 6044 5395 7006 5414
rect 6044 5390 6116 5395
rect 6044 5356 6063 5390
rect 6097 5356 6116 5390
rect 6044 5300 6116 5356
rect 6934 5356 7006 5395
rect 6044 5266 6063 5300
rect 6097 5266 6116 5300
rect 6044 5210 6116 5266
rect 6044 5176 6063 5210
rect 6097 5176 6116 5210
rect 6044 5120 6116 5176
rect 6044 5086 6063 5120
rect 6097 5086 6116 5120
rect 6044 5030 6116 5086
rect 6044 4996 6063 5030
rect 6097 4996 6116 5030
rect 6044 4940 6116 4996
rect 6044 4906 6063 4940
rect 6097 4906 6116 4940
rect 6044 4850 6116 4906
rect 6044 4816 6063 4850
rect 6097 4816 6116 4850
rect 6044 4760 6116 4816
rect 6044 4726 6063 4760
rect 6097 4726 6116 4760
rect 6044 4670 6116 4726
rect 6044 4636 6063 4670
rect 6097 4636 6116 4670
rect 6934 5322 6953 5356
rect 6987 5322 7006 5356
rect 6934 5266 7006 5322
rect 6934 5232 6953 5266
rect 6987 5232 7006 5266
rect 6934 5176 7006 5232
rect 6934 5142 6953 5176
rect 6987 5142 7006 5176
rect 6934 5086 7006 5142
rect 6934 5052 6953 5086
rect 6987 5052 7006 5086
rect 6934 4996 7006 5052
rect 6934 4962 6953 4996
rect 6987 4962 7006 4996
rect 6934 4906 7006 4962
rect 6934 4872 6953 4906
rect 6987 4872 7006 4906
rect 6934 4816 7006 4872
rect 6934 4782 6953 4816
rect 6987 4782 7006 4816
rect 6934 4726 7006 4782
rect 6934 4692 6953 4726
rect 6987 4692 7006 4726
rect 6044 4577 6116 4636
rect 6934 4636 7006 4692
rect 6934 4602 6953 4636
rect 6987 4602 7006 4636
rect 6934 4577 7006 4602
rect 6044 4558 7006 4577
rect 6044 4524 6120 4558
rect 6154 4524 6210 4558
rect 6244 4524 6300 4558
rect 6334 4524 6390 4558
rect 6424 4524 6480 4558
rect 6514 4524 6570 4558
rect 6604 4524 6660 4558
rect 6694 4524 6750 4558
rect 6784 4524 6840 4558
rect 6874 4524 7006 4558
rect 6044 4505 7006 4524
rect 492 4060 1454 4079
rect 492 4026 587 4060
rect 621 4026 677 4060
rect 711 4026 767 4060
rect 801 4026 857 4060
rect 891 4026 947 4060
rect 981 4026 1037 4060
rect 1071 4026 1127 4060
rect 1161 4026 1217 4060
rect 1251 4026 1307 4060
rect 1341 4026 1454 4060
rect 492 4007 1454 4026
rect 492 4002 564 4007
rect 492 3968 511 4002
rect 545 3968 564 4002
rect 492 3912 564 3968
rect 1382 3968 1454 4007
rect 492 3878 511 3912
rect 545 3878 564 3912
rect 492 3822 564 3878
rect 492 3788 511 3822
rect 545 3788 564 3822
rect 492 3732 564 3788
rect 492 3698 511 3732
rect 545 3698 564 3732
rect 492 3642 564 3698
rect 492 3608 511 3642
rect 545 3608 564 3642
rect 492 3552 564 3608
rect 492 3518 511 3552
rect 545 3518 564 3552
rect 492 3462 564 3518
rect 492 3428 511 3462
rect 545 3428 564 3462
rect 492 3372 564 3428
rect 492 3338 511 3372
rect 545 3338 564 3372
rect 492 3282 564 3338
rect 492 3248 511 3282
rect 545 3248 564 3282
rect 1382 3934 1401 3968
rect 1435 3934 1454 3968
rect 1382 3878 1454 3934
rect 1382 3844 1401 3878
rect 1435 3844 1454 3878
rect 1382 3788 1454 3844
rect 1382 3754 1401 3788
rect 1435 3754 1454 3788
rect 1382 3698 1454 3754
rect 1382 3664 1401 3698
rect 1435 3664 1454 3698
rect 1382 3608 1454 3664
rect 1382 3574 1401 3608
rect 1435 3574 1454 3608
rect 1382 3518 1454 3574
rect 1382 3484 1401 3518
rect 1435 3484 1454 3518
rect 1382 3428 1454 3484
rect 1382 3394 1401 3428
rect 1435 3394 1454 3428
rect 1382 3338 1454 3394
rect 1382 3304 1401 3338
rect 1435 3304 1454 3338
rect 492 3189 564 3248
rect 1382 3248 1454 3304
rect 1382 3214 1401 3248
rect 1435 3214 1454 3248
rect 1382 3189 1454 3214
rect 492 3170 1454 3189
rect 492 3136 568 3170
rect 602 3136 658 3170
rect 692 3136 748 3170
rect 782 3136 838 3170
rect 872 3136 928 3170
rect 962 3136 1018 3170
rect 1052 3136 1108 3170
rect 1142 3136 1198 3170
rect 1232 3136 1288 3170
rect 1322 3136 1454 3170
rect 492 3117 1454 3136
rect 1880 4060 2842 4079
rect 1880 4026 1975 4060
rect 2009 4026 2065 4060
rect 2099 4026 2155 4060
rect 2189 4026 2245 4060
rect 2279 4026 2335 4060
rect 2369 4026 2425 4060
rect 2459 4026 2515 4060
rect 2549 4026 2605 4060
rect 2639 4026 2695 4060
rect 2729 4026 2842 4060
rect 1880 4007 2842 4026
rect 1880 4002 1952 4007
rect 1880 3968 1899 4002
rect 1933 3968 1952 4002
rect 1880 3912 1952 3968
rect 2770 3968 2842 4007
rect 1880 3878 1899 3912
rect 1933 3878 1952 3912
rect 1880 3822 1952 3878
rect 1880 3788 1899 3822
rect 1933 3788 1952 3822
rect 1880 3732 1952 3788
rect 1880 3698 1899 3732
rect 1933 3698 1952 3732
rect 1880 3642 1952 3698
rect 1880 3608 1899 3642
rect 1933 3608 1952 3642
rect 1880 3552 1952 3608
rect 1880 3518 1899 3552
rect 1933 3518 1952 3552
rect 1880 3462 1952 3518
rect 1880 3428 1899 3462
rect 1933 3428 1952 3462
rect 1880 3372 1952 3428
rect 1880 3338 1899 3372
rect 1933 3338 1952 3372
rect 1880 3282 1952 3338
rect 1880 3248 1899 3282
rect 1933 3248 1952 3282
rect 2770 3934 2789 3968
rect 2823 3934 2842 3968
rect 2770 3878 2842 3934
rect 2770 3844 2789 3878
rect 2823 3844 2842 3878
rect 2770 3788 2842 3844
rect 2770 3754 2789 3788
rect 2823 3754 2842 3788
rect 2770 3698 2842 3754
rect 2770 3664 2789 3698
rect 2823 3664 2842 3698
rect 2770 3608 2842 3664
rect 2770 3574 2789 3608
rect 2823 3574 2842 3608
rect 2770 3518 2842 3574
rect 2770 3484 2789 3518
rect 2823 3484 2842 3518
rect 2770 3428 2842 3484
rect 2770 3394 2789 3428
rect 2823 3394 2842 3428
rect 2770 3338 2842 3394
rect 2770 3304 2789 3338
rect 2823 3304 2842 3338
rect 1880 3189 1952 3248
rect 2770 3248 2842 3304
rect 2770 3214 2789 3248
rect 2823 3214 2842 3248
rect 2770 3189 2842 3214
rect 1880 3170 2842 3189
rect 1880 3136 1956 3170
rect 1990 3136 2046 3170
rect 2080 3136 2136 3170
rect 2170 3136 2226 3170
rect 2260 3136 2316 3170
rect 2350 3136 2406 3170
rect 2440 3136 2496 3170
rect 2530 3136 2586 3170
rect 2620 3136 2676 3170
rect 2710 3136 2842 3170
rect 1880 3117 2842 3136
rect 3268 4060 4230 4079
rect 3268 4026 3363 4060
rect 3397 4026 3453 4060
rect 3487 4026 3543 4060
rect 3577 4026 3633 4060
rect 3667 4026 3723 4060
rect 3757 4026 3813 4060
rect 3847 4026 3903 4060
rect 3937 4026 3993 4060
rect 4027 4026 4083 4060
rect 4117 4026 4230 4060
rect 3268 4007 4230 4026
rect 3268 4002 3340 4007
rect 3268 3968 3287 4002
rect 3321 3968 3340 4002
rect 3268 3912 3340 3968
rect 4158 3968 4230 4007
rect 3268 3878 3287 3912
rect 3321 3878 3340 3912
rect 3268 3822 3340 3878
rect 3268 3788 3287 3822
rect 3321 3788 3340 3822
rect 3268 3732 3340 3788
rect 3268 3698 3287 3732
rect 3321 3698 3340 3732
rect 3268 3642 3340 3698
rect 3268 3608 3287 3642
rect 3321 3608 3340 3642
rect 3268 3552 3340 3608
rect 3268 3518 3287 3552
rect 3321 3518 3340 3552
rect 3268 3462 3340 3518
rect 3268 3428 3287 3462
rect 3321 3428 3340 3462
rect 3268 3372 3340 3428
rect 3268 3338 3287 3372
rect 3321 3338 3340 3372
rect 3268 3282 3340 3338
rect 3268 3248 3287 3282
rect 3321 3248 3340 3282
rect 4158 3934 4177 3968
rect 4211 3934 4230 3968
rect 4158 3878 4230 3934
rect 4158 3844 4177 3878
rect 4211 3844 4230 3878
rect 4158 3788 4230 3844
rect 4158 3754 4177 3788
rect 4211 3754 4230 3788
rect 4158 3698 4230 3754
rect 4158 3664 4177 3698
rect 4211 3664 4230 3698
rect 4158 3608 4230 3664
rect 4158 3574 4177 3608
rect 4211 3574 4230 3608
rect 4158 3518 4230 3574
rect 4158 3484 4177 3518
rect 4211 3484 4230 3518
rect 4158 3428 4230 3484
rect 4158 3394 4177 3428
rect 4211 3394 4230 3428
rect 4158 3338 4230 3394
rect 4158 3304 4177 3338
rect 4211 3304 4230 3338
rect 3268 3189 3340 3248
rect 4158 3248 4230 3304
rect 4158 3214 4177 3248
rect 4211 3214 4230 3248
rect 4158 3189 4230 3214
rect 3268 3170 4230 3189
rect 3268 3136 3344 3170
rect 3378 3136 3434 3170
rect 3468 3136 3524 3170
rect 3558 3136 3614 3170
rect 3648 3136 3704 3170
rect 3738 3136 3794 3170
rect 3828 3136 3884 3170
rect 3918 3136 3974 3170
rect 4008 3136 4064 3170
rect 4098 3136 4230 3170
rect 3268 3117 4230 3136
rect 4656 4060 5618 4079
rect 4656 4026 4751 4060
rect 4785 4026 4841 4060
rect 4875 4026 4931 4060
rect 4965 4026 5021 4060
rect 5055 4026 5111 4060
rect 5145 4026 5201 4060
rect 5235 4026 5291 4060
rect 5325 4026 5381 4060
rect 5415 4026 5471 4060
rect 5505 4026 5618 4060
rect 4656 4007 5618 4026
rect 4656 4002 4728 4007
rect 4656 3968 4675 4002
rect 4709 3968 4728 4002
rect 4656 3912 4728 3968
rect 5546 3968 5618 4007
rect 4656 3878 4675 3912
rect 4709 3878 4728 3912
rect 4656 3822 4728 3878
rect 4656 3788 4675 3822
rect 4709 3788 4728 3822
rect 4656 3732 4728 3788
rect 4656 3698 4675 3732
rect 4709 3698 4728 3732
rect 4656 3642 4728 3698
rect 4656 3608 4675 3642
rect 4709 3608 4728 3642
rect 4656 3552 4728 3608
rect 4656 3518 4675 3552
rect 4709 3518 4728 3552
rect 4656 3462 4728 3518
rect 4656 3428 4675 3462
rect 4709 3428 4728 3462
rect 4656 3372 4728 3428
rect 4656 3338 4675 3372
rect 4709 3338 4728 3372
rect 4656 3282 4728 3338
rect 4656 3248 4675 3282
rect 4709 3248 4728 3282
rect 5546 3934 5565 3968
rect 5599 3934 5618 3968
rect 5546 3878 5618 3934
rect 5546 3844 5565 3878
rect 5599 3844 5618 3878
rect 5546 3788 5618 3844
rect 5546 3754 5565 3788
rect 5599 3754 5618 3788
rect 5546 3698 5618 3754
rect 5546 3664 5565 3698
rect 5599 3664 5618 3698
rect 5546 3608 5618 3664
rect 5546 3574 5565 3608
rect 5599 3574 5618 3608
rect 5546 3518 5618 3574
rect 5546 3484 5565 3518
rect 5599 3484 5618 3518
rect 5546 3428 5618 3484
rect 5546 3394 5565 3428
rect 5599 3394 5618 3428
rect 5546 3338 5618 3394
rect 5546 3304 5565 3338
rect 5599 3304 5618 3338
rect 4656 3189 4728 3248
rect 5546 3248 5618 3304
rect 5546 3214 5565 3248
rect 5599 3214 5618 3248
rect 5546 3189 5618 3214
rect 4656 3170 5618 3189
rect 4656 3136 4732 3170
rect 4766 3136 4822 3170
rect 4856 3136 4912 3170
rect 4946 3136 5002 3170
rect 5036 3136 5092 3170
rect 5126 3136 5182 3170
rect 5216 3136 5272 3170
rect 5306 3136 5362 3170
rect 5396 3136 5452 3170
rect 5486 3136 5618 3170
rect 4656 3117 5618 3136
rect 6044 4060 7006 4079
rect 6044 4026 6139 4060
rect 6173 4026 6229 4060
rect 6263 4026 6319 4060
rect 6353 4026 6409 4060
rect 6443 4026 6499 4060
rect 6533 4026 6589 4060
rect 6623 4026 6679 4060
rect 6713 4026 6769 4060
rect 6803 4026 6859 4060
rect 6893 4026 7006 4060
rect 6044 4007 7006 4026
rect 6044 4002 6116 4007
rect 6044 3968 6063 4002
rect 6097 3968 6116 4002
rect 6044 3912 6116 3968
rect 6934 3968 7006 4007
rect 6044 3878 6063 3912
rect 6097 3878 6116 3912
rect 6044 3822 6116 3878
rect 6044 3788 6063 3822
rect 6097 3788 6116 3822
rect 6044 3732 6116 3788
rect 6044 3698 6063 3732
rect 6097 3698 6116 3732
rect 6044 3642 6116 3698
rect 6044 3608 6063 3642
rect 6097 3608 6116 3642
rect 6044 3552 6116 3608
rect 6044 3518 6063 3552
rect 6097 3518 6116 3552
rect 6044 3462 6116 3518
rect 6044 3428 6063 3462
rect 6097 3428 6116 3462
rect 6044 3372 6116 3428
rect 6044 3338 6063 3372
rect 6097 3338 6116 3372
rect 6044 3282 6116 3338
rect 6044 3248 6063 3282
rect 6097 3248 6116 3282
rect 6934 3934 6953 3968
rect 6987 3934 7006 3968
rect 6934 3878 7006 3934
rect 6934 3844 6953 3878
rect 6987 3844 7006 3878
rect 6934 3788 7006 3844
rect 6934 3754 6953 3788
rect 6987 3754 7006 3788
rect 6934 3698 7006 3754
rect 6934 3664 6953 3698
rect 6987 3664 7006 3698
rect 6934 3608 7006 3664
rect 6934 3574 6953 3608
rect 6987 3574 7006 3608
rect 6934 3518 7006 3574
rect 6934 3484 6953 3518
rect 6987 3484 7006 3518
rect 6934 3428 7006 3484
rect 6934 3394 6953 3428
rect 6987 3394 7006 3428
rect 6934 3338 7006 3394
rect 6934 3304 6953 3338
rect 6987 3304 7006 3338
rect 6044 3189 6116 3248
rect 6934 3248 7006 3304
rect 6934 3214 6953 3248
rect 6987 3214 7006 3248
rect 6934 3189 7006 3214
rect 6044 3170 7006 3189
rect 6044 3136 6120 3170
rect 6154 3136 6210 3170
rect 6244 3136 6300 3170
rect 6334 3136 6390 3170
rect 6424 3136 6480 3170
rect 6514 3136 6570 3170
rect 6604 3136 6660 3170
rect 6694 3136 6750 3170
rect 6784 3136 6840 3170
rect 6874 3136 7006 3170
rect 6044 3117 7006 3136
rect 492 2672 1454 2691
rect 492 2638 587 2672
rect 621 2638 677 2672
rect 711 2638 767 2672
rect 801 2638 857 2672
rect 891 2638 947 2672
rect 981 2638 1037 2672
rect 1071 2638 1127 2672
rect 1161 2638 1217 2672
rect 1251 2638 1307 2672
rect 1341 2638 1454 2672
rect 492 2619 1454 2638
rect 492 2614 564 2619
rect 492 2580 511 2614
rect 545 2580 564 2614
rect 492 2524 564 2580
rect 1382 2580 1454 2619
rect 492 2490 511 2524
rect 545 2490 564 2524
rect 492 2434 564 2490
rect 492 2400 511 2434
rect 545 2400 564 2434
rect 492 2344 564 2400
rect 492 2310 511 2344
rect 545 2310 564 2344
rect 492 2254 564 2310
rect 492 2220 511 2254
rect 545 2220 564 2254
rect 492 2164 564 2220
rect 492 2130 511 2164
rect 545 2130 564 2164
rect 492 2074 564 2130
rect 492 2040 511 2074
rect 545 2040 564 2074
rect 492 1984 564 2040
rect 492 1950 511 1984
rect 545 1950 564 1984
rect 492 1894 564 1950
rect 492 1860 511 1894
rect 545 1860 564 1894
rect 1382 2546 1401 2580
rect 1435 2546 1454 2580
rect 1382 2490 1454 2546
rect 1382 2456 1401 2490
rect 1435 2456 1454 2490
rect 1382 2400 1454 2456
rect 1382 2366 1401 2400
rect 1435 2366 1454 2400
rect 1382 2310 1454 2366
rect 1382 2276 1401 2310
rect 1435 2276 1454 2310
rect 1382 2220 1454 2276
rect 1382 2186 1401 2220
rect 1435 2186 1454 2220
rect 1382 2130 1454 2186
rect 1382 2096 1401 2130
rect 1435 2096 1454 2130
rect 1382 2040 1454 2096
rect 1382 2006 1401 2040
rect 1435 2006 1454 2040
rect 1382 1950 1454 2006
rect 1382 1916 1401 1950
rect 1435 1916 1454 1950
rect 492 1801 564 1860
rect 1382 1860 1454 1916
rect 1382 1826 1401 1860
rect 1435 1826 1454 1860
rect 1382 1801 1454 1826
rect 492 1782 1454 1801
rect 492 1748 568 1782
rect 602 1748 658 1782
rect 692 1748 748 1782
rect 782 1748 838 1782
rect 872 1748 928 1782
rect 962 1748 1018 1782
rect 1052 1748 1108 1782
rect 1142 1748 1198 1782
rect 1232 1748 1288 1782
rect 1322 1748 1454 1782
rect 492 1729 1454 1748
rect 1880 2672 2842 2691
rect 1880 2638 1975 2672
rect 2009 2638 2065 2672
rect 2099 2638 2155 2672
rect 2189 2638 2245 2672
rect 2279 2638 2335 2672
rect 2369 2638 2425 2672
rect 2459 2638 2515 2672
rect 2549 2638 2605 2672
rect 2639 2638 2695 2672
rect 2729 2638 2842 2672
rect 1880 2619 2842 2638
rect 1880 2614 1952 2619
rect 1880 2580 1899 2614
rect 1933 2580 1952 2614
rect 1880 2524 1952 2580
rect 2770 2580 2842 2619
rect 1880 2490 1899 2524
rect 1933 2490 1952 2524
rect 1880 2434 1952 2490
rect 1880 2400 1899 2434
rect 1933 2400 1952 2434
rect 1880 2344 1952 2400
rect 1880 2310 1899 2344
rect 1933 2310 1952 2344
rect 1880 2254 1952 2310
rect 1880 2220 1899 2254
rect 1933 2220 1952 2254
rect 1880 2164 1952 2220
rect 1880 2130 1899 2164
rect 1933 2130 1952 2164
rect 1880 2074 1952 2130
rect 1880 2040 1899 2074
rect 1933 2040 1952 2074
rect 1880 1984 1952 2040
rect 1880 1950 1899 1984
rect 1933 1950 1952 1984
rect 1880 1894 1952 1950
rect 1880 1860 1899 1894
rect 1933 1860 1952 1894
rect 2770 2546 2789 2580
rect 2823 2546 2842 2580
rect 2770 2490 2842 2546
rect 2770 2456 2789 2490
rect 2823 2456 2842 2490
rect 2770 2400 2842 2456
rect 2770 2366 2789 2400
rect 2823 2366 2842 2400
rect 2770 2310 2842 2366
rect 2770 2276 2789 2310
rect 2823 2276 2842 2310
rect 2770 2220 2842 2276
rect 2770 2186 2789 2220
rect 2823 2186 2842 2220
rect 2770 2130 2842 2186
rect 2770 2096 2789 2130
rect 2823 2096 2842 2130
rect 2770 2040 2842 2096
rect 2770 2006 2789 2040
rect 2823 2006 2842 2040
rect 2770 1950 2842 2006
rect 2770 1916 2789 1950
rect 2823 1916 2842 1950
rect 1880 1801 1952 1860
rect 2770 1860 2842 1916
rect 2770 1826 2789 1860
rect 2823 1826 2842 1860
rect 2770 1801 2842 1826
rect 1880 1782 2842 1801
rect 1880 1748 1956 1782
rect 1990 1748 2046 1782
rect 2080 1748 2136 1782
rect 2170 1748 2226 1782
rect 2260 1748 2316 1782
rect 2350 1748 2406 1782
rect 2440 1748 2496 1782
rect 2530 1748 2586 1782
rect 2620 1748 2676 1782
rect 2710 1748 2842 1782
rect 1880 1729 2842 1748
rect 3268 2672 4230 2691
rect 3268 2638 3363 2672
rect 3397 2638 3453 2672
rect 3487 2638 3543 2672
rect 3577 2638 3633 2672
rect 3667 2638 3723 2672
rect 3757 2638 3813 2672
rect 3847 2638 3903 2672
rect 3937 2638 3993 2672
rect 4027 2638 4083 2672
rect 4117 2638 4230 2672
rect 3268 2619 4230 2638
rect 3268 2614 3340 2619
rect 3268 2580 3287 2614
rect 3321 2580 3340 2614
rect 3268 2524 3340 2580
rect 4158 2580 4230 2619
rect 3268 2490 3287 2524
rect 3321 2490 3340 2524
rect 3268 2434 3340 2490
rect 3268 2400 3287 2434
rect 3321 2400 3340 2434
rect 3268 2344 3340 2400
rect 3268 2310 3287 2344
rect 3321 2310 3340 2344
rect 3268 2254 3340 2310
rect 3268 2220 3287 2254
rect 3321 2220 3340 2254
rect 3268 2164 3340 2220
rect 3268 2130 3287 2164
rect 3321 2130 3340 2164
rect 3268 2074 3340 2130
rect 3268 2040 3287 2074
rect 3321 2040 3340 2074
rect 3268 1984 3340 2040
rect 3268 1950 3287 1984
rect 3321 1950 3340 1984
rect 3268 1894 3340 1950
rect 3268 1860 3287 1894
rect 3321 1860 3340 1894
rect 4158 2546 4177 2580
rect 4211 2546 4230 2580
rect 4158 2490 4230 2546
rect 4158 2456 4177 2490
rect 4211 2456 4230 2490
rect 4158 2400 4230 2456
rect 4158 2366 4177 2400
rect 4211 2366 4230 2400
rect 4158 2310 4230 2366
rect 4158 2276 4177 2310
rect 4211 2276 4230 2310
rect 4158 2220 4230 2276
rect 4158 2186 4177 2220
rect 4211 2186 4230 2220
rect 4158 2130 4230 2186
rect 4158 2096 4177 2130
rect 4211 2096 4230 2130
rect 4158 2040 4230 2096
rect 4158 2006 4177 2040
rect 4211 2006 4230 2040
rect 4158 1950 4230 2006
rect 4158 1916 4177 1950
rect 4211 1916 4230 1950
rect 3268 1801 3340 1860
rect 4158 1860 4230 1916
rect 4158 1826 4177 1860
rect 4211 1826 4230 1860
rect 4158 1801 4230 1826
rect 3268 1782 4230 1801
rect 3268 1748 3344 1782
rect 3378 1748 3434 1782
rect 3468 1748 3524 1782
rect 3558 1748 3614 1782
rect 3648 1748 3704 1782
rect 3738 1748 3794 1782
rect 3828 1748 3884 1782
rect 3918 1748 3974 1782
rect 4008 1748 4064 1782
rect 4098 1748 4230 1782
rect 3268 1729 4230 1748
rect 4656 2672 5618 2691
rect 4656 2638 4751 2672
rect 4785 2638 4841 2672
rect 4875 2638 4931 2672
rect 4965 2638 5021 2672
rect 5055 2638 5111 2672
rect 5145 2638 5201 2672
rect 5235 2638 5291 2672
rect 5325 2638 5381 2672
rect 5415 2638 5471 2672
rect 5505 2638 5618 2672
rect 4656 2619 5618 2638
rect 4656 2614 4728 2619
rect 4656 2580 4675 2614
rect 4709 2580 4728 2614
rect 4656 2524 4728 2580
rect 5546 2580 5618 2619
rect 4656 2490 4675 2524
rect 4709 2490 4728 2524
rect 4656 2434 4728 2490
rect 4656 2400 4675 2434
rect 4709 2400 4728 2434
rect 4656 2344 4728 2400
rect 4656 2310 4675 2344
rect 4709 2310 4728 2344
rect 4656 2254 4728 2310
rect 4656 2220 4675 2254
rect 4709 2220 4728 2254
rect 4656 2164 4728 2220
rect 4656 2130 4675 2164
rect 4709 2130 4728 2164
rect 4656 2074 4728 2130
rect 4656 2040 4675 2074
rect 4709 2040 4728 2074
rect 4656 1984 4728 2040
rect 4656 1950 4675 1984
rect 4709 1950 4728 1984
rect 4656 1894 4728 1950
rect 4656 1860 4675 1894
rect 4709 1860 4728 1894
rect 5546 2546 5565 2580
rect 5599 2546 5618 2580
rect 5546 2490 5618 2546
rect 5546 2456 5565 2490
rect 5599 2456 5618 2490
rect 5546 2400 5618 2456
rect 5546 2366 5565 2400
rect 5599 2366 5618 2400
rect 5546 2310 5618 2366
rect 5546 2276 5565 2310
rect 5599 2276 5618 2310
rect 5546 2220 5618 2276
rect 5546 2186 5565 2220
rect 5599 2186 5618 2220
rect 5546 2130 5618 2186
rect 5546 2096 5565 2130
rect 5599 2096 5618 2130
rect 5546 2040 5618 2096
rect 5546 2006 5565 2040
rect 5599 2006 5618 2040
rect 5546 1950 5618 2006
rect 5546 1916 5565 1950
rect 5599 1916 5618 1950
rect 4656 1801 4728 1860
rect 5546 1860 5618 1916
rect 5546 1826 5565 1860
rect 5599 1826 5618 1860
rect 5546 1801 5618 1826
rect 4656 1782 5618 1801
rect 4656 1748 4732 1782
rect 4766 1748 4822 1782
rect 4856 1748 4912 1782
rect 4946 1748 5002 1782
rect 5036 1748 5092 1782
rect 5126 1748 5182 1782
rect 5216 1748 5272 1782
rect 5306 1748 5362 1782
rect 5396 1748 5452 1782
rect 5486 1748 5618 1782
rect 4656 1729 5618 1748
rect 6044 2672 7006 2691
rect 6044 2638 6139 2672
rect 6173 2638 6229 2672
rect 6263 2638 6319 2672
rect 6353 2638 6409 2672
rect 6443 2638 6499 2672
rect 6533 2638 6589 2672
rect 6623 2638 6679 2672
rect 6713 2638 6769 2672
rect 6803 2638 6859 2672
rect 6893 2638 7006 2672
rect 6044 2619 7006 2638
rect 6044 2614 6116 2619
rect 6044 2580 6063 2614
rect 6097 2580 6116 2614
rect 6044 2524 6116 2580
rect 6934 2580 7006 2619
rect 6044 2490 6063 2524
rect 6097 2490 6116 2524
rect 6044 2434 6116 2490
rect 6044 2400 6063 2434
rect 6097 2400 6116 2434
rect 6044 2344 6116 2400
rect 6044 2310 6063 2344
rect 6097 2310 6116 2344
rect 6044 2254 6116 2310
rect 6044 2220 6063 2254
rect 6097 2220 6116 2254
rect 6044 2164 6116 2220
rect 6044 2130 6063 2164
rect 6097 2130 6116 2164
rect 6044 2074 6116 2130
rect 6044 2040 6063 2074
rect 6097 2040 6116 2074
rect 6044 1984 6116 2040
rect 6044 1950 6063 1984
rect 6097 1950 6116 1984
rect 6044 1894 6116 1950
rect 6044 1860 6063 1894
rect 6097 1860 6116 1894
rect 6934 2546 6953 2580
rect 6987 2546 7006 2580
rect 6934 2490 7006 2546
rect 6934 2456 6953 2490
rect 6987 2456 7006 2490
rect 6934 2400 7006 2456
rect 6934 2366 6953 2400
rect 6987 2366 7006 2400
rect 6934 2310 7006 2366
rect 6934 2276 6953 2310
rect 6987 2276 7006 2310
rect 6934 2220 7006 2276
rect 6934 2186 6953 2220
rect 6987 2186 7006 2220
rect 6934 2130 7006 2186
rect 6934 2096 6953 2130
rect 6987 2096 7006 2130
rect 6934 2040 7006 2096
rect 6934 2006 6953 2040
rect 6987 2006 7006 2040
rect 6934 1950 7006 2006
rect 6934 1916 6953 1950
rect 6987 1916 7006 1950
rect 6044 1801 6116 1860
rect 6934 1860 7006 1916
rect 6934 1826 6953 1860
rect 6987 1826 7006 1860
rect 6934 1801 7006 1826
rect 6044 1782 7006 1801
rect 6044 1748 6120 1782
rect 6154 1748 6210 1782
rect 6244 1748 6300 1782
rect 6334 1748 6390 1782
rect 6424 1748 6480 1782
rect 6514 1748 6570 1782
rect 6604 1748 6660 1782
rect 6694 1748 6750 1782
rect 6784 1748 6840 1782
rect 6874 1748 7006 1782
rect 6044 1729 7006 1748
rect -17957 -381 -17883 -375
rect 9147 -375 9167 22941
rect 9201 -375 9221 22941
rect 9147 -381 9221 -375
rect -17957 -401 9221 -381
rect -17957 -435 -17877 -401
rect 9141 -435 9221 -401
rect -17957 -455 9221 -435
<< psubdiffcont >>
rect -17440 22657 8642 22691
rect -17500 20912 -17466 22631
rect 8668 20912 8702 22631
rect -17440 20852 8642 20886
rect -13053 20761 8591 20795
rect -13149 19399 -13115 20699
rect 8653 19399 8687 20699
rect -13053 19303 8591 19337
rect -7069 19197 8591 19231
rect -7165 17835 -7131 19135
rect 8653 17835 8687 19135
rect -7069 17739 8591 17773
rect -1210 17574 -404 17608
rect -1270 16854 -1236 17541
rect -378 16843 -344 17541
rect -1210 16786 -404 16820
rect -149 17587 8627 17621
rect -209 15985 -175 17539
rect 8653 15985 8687 17539
rect -149 15925 8627 15959
rect -1160 15829 2568 15863
rect -1220 14763 -1186 15803
rect 2594 14763 2628 15803
rect 2927 15744 8625 15778
rect 2865 14861 2899 15703
rect 8653 14861 8687 15703
rect 2927 14786 8625 14820
rect -1160 14703 2568 14737
rect 664 12297 1470 12331
rect 1556 12297 2362 12331
rect 2448 12297 3254 12331
rect 3340 12297 4146 12331
rect 604 10291 638 12271
rect 1496 10291 1530 12271
rect 2388 10291 2422 12271
rect 3280 10291 3314 12271
rect 4172 10291 4206 12271
rect 4320 12267 4712 12301
rect 4260 11435 4294 12241
rect 4738 11435 4772 12241
rect 4320 11375 4712 11409
rect 664 10231 1470 10265
rect 1556 10231 2362 10265
rect 2448 10231 3254 10265
rect 3340 10231 4146 10265
rect 4320 11153 4712 11187
rect 4260 10321 4294 11127
rect 4738 10321 4772 11127
rect 4320 10261 4712 10295
rect 387 8339 421 8373
rect 477 8339 511 8373
rect 567 8339 601 8373
rect 657 8339 691 8373
rect 747 8339 781 8373
rect 837 8339 871 8373
rect 927 8339 961 8373
rect 1017 8339 1051 8373
rect 1107 8339 1141 8373
rect 1197 8339 1231 8373
rect 1287 8339 1321 8373
rect 1377 8339 1411 8373
rect 1467 8339 1501 8373
rect 364 8238 398 8272
rect 364 8148 398 8182
rect 364 8058 398 8092
rect 364 7968 398 8002
rect 364 7878 398 7912
rect 364 7788 398 7822
rect 364 7698 398 7732
rect 364 7608 398 7642
rect 364 7518 398 7552
rect 364 7428 398 7462
rect 364 7338 398 7372
rect 364 7248 398 7282
rect 1551 8238 1585 8272
rect 1551 8148 1585 8182
rect 1551 8058 1585 8092
rect 1551 7968 1585 8002
rect 1551 7878 1585 7912
rect 1551 7788 1585 7822
rect 1551 7698 1585 7732
rect 1551 7608 1585 7642
rect 1551 7518 1585 7552
rect 1551 7428 1585 7462
rect 1551 7338 1585 7372
rect 1551 7248 1585 7282
rect 387 7152 421 7186
rect 477 7152 511 7186
rect 567 7152 601 7186
rect 657 7152 691 7186
rect 747 7152 781 7186
rect 837 7152 871 7186
rect 927 7152 961 7186
rect 1017 7152 1051 7186
rect 1107 7152 1141 7186
rect 1197 7152 1231 7186
rect 1287 7152 1321 7186
rect 1377 7152 1411 7186
rect 1467 7152 1501 7186
rect 1775 8339 1809 8373
rect 1865 8339 1899 8373
rect 1955 8339 1989 8373
rect 2045 8339 2079 8373
rect 2135 8339 2169 8373
rect 2225 8339 2259 8373
rect 2315 8339 2349 8373
rect 2405 8339 2439 8373
rect 2495 8339 2529 8373
rect 2585 8339 2619 8373
rect 2675 8339 2709 8373
rect 2765 8339 2799 8373
rect 2855 8339 2889 8373
rect 1752 8238 1786 8272
rect 1752 8148 1786 8182
rect 1752 8058 1786 8092
rect 1752 7968 1786 8002
rect 1752 7878 1786 7912
rect 1752 7788 1786 7822
rect 1752 7698 1786 7732
rect 1752 7608 1786 7642
rect 1752 7518 1786 7552
rect 1752 7428 1786 7462
rect 1752 7338 1786 7372
rect 1752 7248 1786 7282
rect 2939 8238 2973 8272
rect 2939 8148 2973 8182
rect 2939 8058 2973 8092
rect 2939 7968 2973 8002
rect 2939 7878 2973 7912
rect 2939 7788 2973 7822
rect 2939 7698 2973 7732
rect 2939 7608 2973 7642
rect 2939 7518 2973 7552
rect 2939 7428 2973 7462
rect 2939 7338 2973 7372
rect 2939 7248 2973 7282
rect 1775 7152 1809 7186
rect 1865 7152 1899 7186
rect 1955 7152 1989 7186
rect 2045 7152 2079 7186
rect 2135 7152 2169 7186
rect 2225 7152 2259 7186
rect 2315 7152 2349 7186
rect 2405 7152 2439 7186
rect 2495 7152 2529 7186
rect 2585 7152 2619 7186
rect 2675 7152 2709 7186
rect 2765 7152 2799 7186
rect 2855 7152 2889 7186
rect 3163 8339 3197 8373
rect 3253 8339 3287 8373
rect 3343 8339 3377 8373
rect 3433 8339 3467 8373
rect 3523 8339 3557 8373
rect 3613 8339 3647 8373
rect 3703 8339 3737 8373
rect 3793 8339 3827 8373
rect 3883 8339 3917 8373
rect 3973 8339 4007 8373
rect 4063 8339 4097 8373
rect 4153 8339 4187 8373
rect 4243 8339 4277 8373
rect 3140 8238 3174 8272
rect 3140 8148 3174 8182
rect 3140 8058 3174 8092
rect 3140 7968 3174 8002
rect 3140 7878 3174 7912
rect 3140 7788 3174 7822
rect 3140 7698 3174 7732
rect 3140 7608 3174 7642
rect 3140 7518 3174 7552
rect 3140 7428 3174 7462
rect 3140 7338 3174 7372
rect 3140 7248 3174 7282
rect 4327 8238 4361 8272
rect 4327 8148 4361 8182
rect 4327 8058 4361 8092
rect 4327 7968 4361 8002
rect 4327 7878 4361 7912
rect 4327 7788 4361 7822
rect 4327 7698 4361 7732
rect 4327 7608 4361 7642
rect 4327 7518 4361 7552
rect 4327 7428 4361 7462
rect 4327 7338 4361 7372
rect 4327 7248 4361 7282
rect 3163 7152 3197 7186
rect 3253 7152 3287 7186
rect 3343 7152 3377 7186
rect 3433 7152 3467 7186
rect 3523 7152 3557 7186
rect 3613 7152 3647 7186
rect 3703 7152 3737 7186
rect 3793 7152 3827 7186
rect 3883 7152 3917 7186
rect 3973 7152 4007 7186
rect 4063 7152 4097 7186
rect 4153 7152 4187 7186
rect 4243 7152 4277 7186
rect 4551 8339 4585 8373
rect 4641 8339 4675 8373
rect 4731 8339 4765 8373
rect 4821 8339 4855 8373
rect 4911 8339 4945 8373
rect 5001 8339 5035 8373
rect 5091 8339 5125 8373
rect 5181 8339 5215 8373
rect 5271 8339 5305 8373
rect 5361 8339 5395 8373
rect 5451 8339 5485 8373
rect 5541 8339 5575 8373
rect 5631 8339 5665 8373
rect 4528 8238 4562 8272
rect 4528 8148 4562 8182
rect 4528 8058 4562 8092
rect 4528 7968 4562 8002
rect 4528 7878 4562 7912
rect 4528 7788 4562 7822
rect 4528 7698 4562 7732
rect 4528 7608 4562 7642
rect 4528 7518 4562 7552
rect 4528 7428 4562 7462
rect 4528 7338 4562 7372
rect 4528 7248 4562 7282
rect 5715 8238 5749 8272
rect 5715 8148 5749 8182
rect 5715 8058 5749 8092
rect 5715 7968 5749 8002
rect 5715 7878 5749 7912
rect 5715 7788 5749 7822
rect 5715 7698 5749 7732
rect 5715 7608 5749 7642
rect 5715 7518 5749 7552
rect 5715 7428 5749 7462
rect 5715 7338 5749 7372
rect 5715 7248 5749 7282
rect 4551 7152 4585 7186
rect 4641 7152 4675 7186
rect 4731 7152 4765 7186
rect 4821 7152 4855 7186
rect 4911 7152 4945 7186
rect 5001 7152 5035 7186
rect 5091 7152 5125 7186
rect 5181 7152 5215 7186
rect 5271 7152 5305 7186
rect 5361 7152 5395 7186
rect 5451 7152 5485 7186
rect 5541 7152 5575 7186
rect 5631 7152 5665 7186
rect 5939 8339 5973 8373
rect 6029 8339 6063 8373
rect 6119 8339 6153 8373
rect 6209 8339 6243 8373
rect 6299 8339 6333 8373
rect 6389 8339 6423 8373
rect 6479 8339 6513 8373
rect 6569 8339 6603 8373
rect 6659 8339 6693 8373
rect 6749 8339 6783 8373
rect 6839 8339 6873 8373
rect 6929 8339 6963 8373
rect 7019 8339 7053 8373
rect 5916 8238 5950 8272
rect 5916 8148 5950 8182
rect 5916 8058 5950 8092
rect 5916 7968 5950 8002
rect 5916 7878 5950 7912
rect 5916 7788 5950 7822
rect 5916 7698 5950 7732
rect 5916 7608 5950 7642
rect 5916 7518 5950 7552
rect 5916 7428 5950 7462
rect 5916 7338 5950 7372
rect 5916 7248 5950 7282
rect 7103 8238 7137 8272
rect 7103 8148 7137 8182
rect 7103 8058 7137 8092
rect 7103 7968 7137 8002
rect 7103 7878 7137 7912
rect 7103 7788 7137 7822
rect 7103 7698 7137 7732
rect 7103 7608 7137 7642
rect 7103 7518 7137 7552
rect 7103 7428 7137 7462
rect 7103 7338 7137 7372
rect 7103 7248 7137 7282
rect 5939 7152 5973 7186
rect 6029 7152 6063 7186
rect 6119 7152 6153 7186
rect 6209 7152 6243 7186
rect 6299 7152 6333 7186
rect 6389 7152 6423 7186
rect 6479 7152 6513 7186
rect 6569 7152 6603 7186
rect 6659 7152 6693 7186
rect 6749 7152 6783 7186
rect 6839 7152 6873 7186
rect 6929 7152 6963 7186
rect 7019 7152 7053 7186
rect 387 6951 421 6985
rect 477 6951 511 6985
rect 567 6951 601 6985
rect 657 6951 691 6985
rect 747 6951 781 6985
rect 837 6951 871 6985
rect 927 6951 961 6985
rect 1017 6951 1051 6985
rect 1107 6951 1141 6985
rect 1197 6951 1231 6985
rect 1287 6951 1321 6985
rect 1377 6951 1411 6985
rect 1467 6951 1501 6985
rect 364 6850 398 6884
rect 364 6760 398 6794
rect 364 6670 398 6704
rect 364 6580 398 6614
rect 364 6490 398 6524
rect 364 6400 398 6434
rect 364 6310 398 6344
rect 364 6220 398 6254
rect 364 6130 398 6164
rect 364 6040 398 6074
rect 364 5950 398 5984
rect 364 5860 398 5894
rect 1551 6850 1585 6884
rect 1551 6760 1585 6794
rect 1551 6670 1585 6704
rect 1551 6580 1585 6614
rect 1551 6490 1585 6524
rect 1551 6400 1585 6434
rect 1551 6310 1585 6344
rect 1551 6220 1585 6254
rect 1551 6130 1585 6164
rect 1551 6040 1585 6074
rect 1551 5950 1585 5984
rect 1551 5860 1585 5894
rect 387 5764 421 5798
rect 477 5764 511 5798
rect 567 5764 601 5798
rect 657 5764 691 5798
rect 747 5764 781 5798
rect 837 5764 871 5798
rect 927 5764 961 5798
rect 1017 5764 1051 5798
rect 1107 5764 1141 5798
rect 1197 5764 1231 5798
rect 1287 5764 1321 5798
rect 1377 5764 1411 5798
rect 1467 5764 1501 5798
rect 1775 6951 1809 6985
rect 1865 6951 1899 6985
rect 1955 6951 1989 6985
rect 2045 6951 2079 6985
rect 2135 6951 2169 6985
rect 2225 6951 2259 6985
rect 2315 6951 2349 6985
rect 2405 6951 2439 6985
rect 2495 6951 2529 6985
rect 2585 6951 2619 6985
rect 2675 6951 2709 6985
rect 2765 6951 2799 6985
rect 2855 6951 2889 6985
rect 1752 6850 1786 6884
rect 1752 6760 1786 6794
rect 1752 6670 1786 6704
rect 1752 6580 1786 6614
rect 1752 6490 1786 6524
rect 1752 6400 1786 6434
rect 1752 6310 1786 6344
rect 1752 6220 1786 6254
rect 1752 6130 1786 6164
rect 1752 6040 1786 6074
rect 1752 5950 1786 5984
rect 1752 5860 1786 5894
rect 2939 6850 2973 6884
rect 2939 6760 2973 6794
rect 2939 6670 2973 6704
rect 2939 6580 2973 6614
rect 2939 6490 2973 6524
rect 2939 6400 2973 6434
rect 2939 6310 2973 6344
rect 2939 6220 2973 6254
rect 2939 6130 2973 6164
rect 2939 6040 2973 6074
rect 2939 5950 2973 5984
rect 2939 5860 2973 5894
rect 1775 5764 1809 5798
rect 1865 5764 1899 5798
rect 1955 5764 1989 5798
rect 2045 5764 2079 5798
rect 2135 5764 2169 5798
rect 2225 5764 2259 5798
rect 2315 5764 2349 5798
rect 2405 5764 2439 5798
rect 2495 5764 2529 5798
rect 2585 5764 2619 5798
rect 2675 5764 2709 5798
rect 2765 5764 2799 5798
rect 2855 5764 2889 5798
rect 3163 6951 3197 6985
rect 3253 6951 3287 6985
rect 3343 6951 3377 6985
rect 3433 6951 3467 6985
rect 3523 6951 3557 6985
rect 3613 6951 3647 6985
rect 3703 6951 3737 6985
rect 3793 6951 3827 6985
rect 3883 6951 3917 6985
rect 3973 6951 4007 6985
rect 4063 6951 4097 6985
rect 4153 6951 4187 6985
rect 4243 6951 4277 6985
rect 3140 6850 3174 6884
rect 3140 6760 3174 6794
rect 3140 6670 3174 6704
rect 3140 6580 3174 6614
rect 3140 6490 3174 6524
rect 3140 6400 3174 6434
rect 3140 6310 3174 6344
rect 3140 6220 3174 6254
rect 3140 6130 3174 6164
rect 3140 6040 3174 6074
rect 3140 5950 3174 5984
rect 3140 5860 3174 5894
rect 4327 6850 4361 6884
rect 4327 6760 4361 6794
rect 4327 6670 4361 6704
rect 4327 6580 4361 6614
rect 4327 6490 4361 6524
rect 4327 6400 4361 6434
rect 4327 6310 4361 6344
rect 4327 6220 4361 6254
rect 4327 6130 4361 6164
rect 4327 6040 4361 6074
rect 4327 5950 4361 5984
rect 4327 5860 4361 5894
rect 3163 5764 3197 5798
rect 3253 5764 3287 5798
rect 3343 5764 3377 5798
rect 3433 5764 3467 5798
rect 3523 5764 3557 5798
rect 3613 5764 3647 5798
rect 3703 5764 3737 5798
rect 3793 5764 3827 5798
rect 3883 5764 3917 5798
rect 3973 5764 4007 5798
rect 4063 5764 4097 5798
rect 4153 5764 4187 5798
rect 4243 5764 4277 5798
rect 4551 6951 4585 6985
rect 4641 6951 4675 6985
rect 4731 6951 4765 6985
rect 4821 6951 4855 6985
rect 4911 6951 4945 6985
rect 5001 6951 5035 6985
rect 5091 6951 5125 6985
rect 5181 6951 5215 6985
rect 5271 6951 5305 6985
rect 5361 6951 5395 6985
rect 5451 6951 5485 6985
rect 5541 6951 5575 6985
rect 5631 6951 5665 6985
rect 4528 6850 4562 6884
rect 4528 6760 4562 6794
rect 4528 6670 4562 6704
rect 4528 6580 4562 6614
rect 4528 6490 4562 6524
rect 4528 6400 4562 6434
rect 4528 6310 4562 6344
rect 4528 6220 4562 6254
rect 4528 6130 4562 6164
rect 4528 6040 4562 6074
rect 4528 5950 4562 5984
rect 4528 5860 4562 5894
rect 5715 6850 5749 6884
rect 5715 6760 5749 6794
rect 5715 6670 5749 6704
rect 5715 6580 5749 6614
rect 5715 6490 5749 6524
rect 5715 6400 5749 6434
rect 5715 6310 5749 6344
rect 5715 6220 5749 6254
rect 5715 6130 5749 6164
rect 5715 6040 5749 6074
rect 5715 5950 5749 5984
rect 5715 5860 5749 5894
rect 4551 5764 4585 5798
rect 4641 5764 4675 5798
rect 4731 5764 4765 5798
rect 4821 5764 4855 5798
rect 4911 5764 4945 5798
rect 5001 5764 5035 5798
rect 5091 5764 5125 5798
rect 5181 5764 5215 5798
rect 5271 5764 5305 5798
rect 5361 5764 5395 5798
rect 5451 5764 5485 5798
rect 5541 5764 5575 5798
rect 5631 5764 5665 5798
rect 5939 6951 5973 6985
rect 6029 6951 6063 6985
rect 6119 6951 6153 6985
rect 6209 6951 6243 6985
rect 6299 6951 6333 6985
rect 6389 6951 6423 6985
rect 6479 6951 6513 6985
rect 6569 6951 6603 6985
rect 6659 6951 6693 6985
rect 6749 6951 6783 6985
rect 6839 6951 6873 6985
rect 6929 6951 6963 6985
rect 7019 6951 7053 6985
rect 5916 6850 5950 6884
rect 5916 6760 5950 6794
rect 5916 6670 5950 6704
rect 5916 6580 5950 6614
rect 5916 6490 5950 6524
rect 5916 6400 5950 6434
rect 5916 6310 5950 6344
rect 5916 6220 5950 6254
rect 5916 6130 5950 6164
rect 5916 6040 5950 6074
rect 5916 5950 5950 5984
rect 5916 5860 5950 5894
rect 7103 6850 7137 6884
rect 7103 6760 7137 6794
rect 7103 6670 7137 6704
rect 7103 6580 7137 6614
rect 7103 6490 7137 6524
rect 7103 6400 7137 6434
rect 7103 6310 7137 6344
rect 7103 6220 7137 6254
rect 7103 6130 7137 6164
rect 7103 6040 7137 6074
rect 7103 5950 7137 5984
rect 7103 5860 7137 5894
rect 5939 5764 5973 5798
rect 6029 5764 6063 5798
rect 6119 5764 6153 5798
rect 6209 5764 6243 5798
rect 6299 5764 6333 5798
rect 6389 5764 6423 5798
rect 6479 5764 6513 5798
rect 6569 5764 6603 5798
rect 6659 5764 6693 5798
rect 6749 5764 6783 5798
rect 6839 5764 6873 5798
rect 6929 5764 6963 5798
rect 7019 5764 7053 5798
rect 387 5563 421 5597
rect 477 5563 511 5597
rect 567 5563 601 5597
rect 657 5563 691 5597
rect 747 5563 781 5597
rect 837 5563 871 5597
rect 927 5563 961 5597
rect 1017 5563 1051 5597
rect 1107 5563 1141 5597
rect 1197 5563 1231 5597
rect 1287 5563 1321 5597
rect 1377 5563 1411 5597
rect 1467 5563 1501 5597
rect 364 5462 398 5496
rect 364 5372 398 5406
rect 364 5282 398 5316
rect 364 5192 398 5226
rect 364 5102 398 5136
rect 364 5012 398 5046
rect 364 4922 398 4956
rect 364 4832 398 4866
rect 364 4742 398 4776
rect 364 4652 398 4686
rect 364 4562 398 4596
rect 364 4472 398 4506
rect 1551 5462 1585 5496
rect 1551 5372 1585 5406
rect 1551 5282 1585 5316
rect 1551 5192 1585 5226
rect 1551 5102 1585 5136
rect 1551 5012 1585 5046
rect 1551 4922 1585 4956
rect 1551 4832 1585 4866
rect 1551 4742 1585 4776
rect 1551 4652 1585 4686
rect 1551 4562 1585 4596
rect 1551 4472 1585 4506
rect 387 4376 421 4410
rect 477 4376 511 4410
rect 567 4376 601 4410
rect 657 4376 691 4410
rect 747 4376 781 4410
rect 837 4376 871 4410
rect 927 4376 961 4410
rect 1017 4376 1051 4410
rect 1107 4376 1141 4410
rect 1197 4376 1231 4410
rect 1287 4376 1321 4410
rect 1377 4376 1411 4410
rect 1467 4376 1501 4410
rect 1775 5563 1809 5597
rect 1865 5563 1899 5597
rect 1955 5563 1989 5597
rect 2045 5563 2079 5597
rect 2135 5563 2169 5597
rect 2225 5563 2259 5597
rect 2315 5563 2349 5597
rect 2405 5563 2439 5597
rect 2495 5563 2529 5597
rect 2585 5563 2619 5597
rect 2675 5563 2709 5597
rect 2765 5563 2799 5597
rect 2855 5563 2889 5597
rect 1752 5462 1786 5496
rect 1752 5372 1786 5406
rect 1752 5282 1786 5316
rect 1752 5192 1786 5226
rect 1752 5102 1786 5136
rect 1752 5012 1786 5046
rect 1752 4922 1786 4956
rect 1752 4832 1786 4866
rect 1752 4742 1786 4776
rect 1752 4652 1786 4686
rect 1752 4562 1786 4596
rect 1752 4472 1786 4506
rect 2939 5462 2973 5496
rect 2939 5372 2973 5406
rect 2939 5282 2973 5316
rect 2939 5192 2973 5226
rect 2939 5102 2973 5136
rect 2939 5012 2973 5046
rect 2939 4922 2973 4956
rect 2939 4832 2973 4866
rect 2939 4742 2973 4776
rect 2939 4652 2973 4686
rect 2939 4562 2973 4596
rect 2939 4472 2973 4506
rect 1775 4376 1809 4410
rect 1865 4376 1899 4410
rect 1955 4376 1989 4410
rect 2045 4376 2079 4410
rect 2135 4376 2169 4410
rect 2225 4376 2259 4410
rect 2315 4376 2349 4410
rect 2405 4376 2439 4410
rect 2495 4376 2529 4410
rect 2585 4376 2619 4410
rect 2675 4376 2709 4410
rect 2765 4376 2799 4410
rect 2855 4376 2889 4410
rect 3163 5563 3197 5597
rect 3253 5563 3287 5597
rect 3343 5563 3377 5597
rect 3433 5563 3467 5597
rect 3523 5563 3557 5597
rect 3613 5563 3647 5597
rect 3703 5563 3737 5597
rect 3793 5563 3827 5597
rect 3883 5563 3917 5597
rect 3973 5563 4007 5597
rect 4063 5563 4097 5597
rect 4153 5563 4187 5597
rect 4243 5563 4277 5597
rect 3140 5462 3174 5496
rect 3140 5372 3174 5406
rect 3140 5282 3174 5316
rect 3140 5192 3174 5226
rect 3140 5102 3174 5136
rect 3140 5012 3174 5046
rect 3140 4922 3174 4956
rect 3140 4832 3174 4866
rect 3140 4742 3174 4776
rect 3140 4652 3174 4686
rect 3140 4562 3174 4596
rect 3140 4472 3174 4506
rect 4327 5462 4361 5496
rect 4327 5372 4361 5406
rect 4327 5282 4361 5316
rect 4327 5192 4361 5226
rect 4327 5102 4361 5136
rect 4327 5012 4361 5046
rect 4327 4922 4361 4956
rect 4327 4832 4361 4866
rect 4327 4742 4361 4776
rect 4327 4652 4361 4686
rect 4327 4562 4361 4596
rect 4327 4472 4361 4506
rect 3163 4376 3197 4410
rect 3253 4376 3287 4410
rect 3343 4376 3377 4410
rect 3433 4376 3467 4410
rect 3523 4376 3557 4410
rect 3613 4376 3647 4410
rect 3703 4376 3737 4410
rect 3793 4376 3827 4410
rect 3883 4376 3917 4410
rect 3973 4376 4007 4410
rect 4063 4376 4097 4410
rect 4153 4376 4187 4410
rect 4243 4376 4277 4410
rect 4551 5563 4585 5597
rect 4641 5563 4675 5597
rect 4731 5563 4765 5597
rect 4821 5563 4855 5597
rect 4911 5563 4945 5597
rect 5001 5563 5035 5597
rect 5091 5563 5125 5597
rect 5181 5563 5215 5597
rect 5271 5563 5305 5597
rect 5361 5563 5395 5597
rect 5451 5563 5485 5597
rect 5541 5563 5575 5597
rect 5631 5563 5665 5597
rect 4528 5462 4562 5496
rect 4528 5372 4562 5406
rect 4528 5282 4562 5316
rect 4528 5192 4562 5226
rect 4528 5102 4562 5136
rect 4528 5012 4562 5046
rect 4528 4922 4562 4956
rect 4528 4832 4562 4866
rect 4528 4742 4562 4776
rect 4528 4652 4562 4686
rect 4528 4562 4562 4596
rect 4528 4472 4562 4506
rect 5715 5462 5749 5496
rect 5715 5372 5749 5406
rect 5715 5282 5749 5316
rect 5715 5192 5749 5226
rect 5715 5102 5749 5136
rect 5715 5012 5749 5046
rect 5715 4922 5749 4956
rect 5715 4832 5749 4866
rect 5715 4742 5749 4776
rect 5715 4652 5749 4686
rect 5715 4562 5749 4596
rect 5715 4472 5749 4506
rect 4551 4376 4585 4410
rect 4641 4376 4675 4410
rect 4731 4376 4765 4410
rect 4821 4376 4855 4410
rect 4911 4376 4945 4410
rect 5001 4376 5035 4410
rect 5091 4376 5125 4410
rect 5181 4376 5215 4410
rect 5271 4376 5305 4410
rect 5361 4376 5395 4410
rect 5451 4376 5485 4410
rect 5541 4376 5575 4410
rect 5631 4376 5665 4410
rect 5939 5563 5973 5597
rect 6029 5563 6063 5597
rect 6119 5563 6153 5597
rect 6209 5563 6243 5597
rect 6299 5563 6333 5597
rect 6389 5563 6423 5597
rect 6479 5563 6513 5597
rect 6569 5563 6603 5597
rect 6659 5563 6693 5597
rect 6749 5563 6783 5597
rect 6839 5563 6873 5597
rect 6929 5563 6963 5597
rect 7019 5563 7053 5597
rect 5916 5462 5950 5496
rect 5916 5372 5950 5406
rect 5916 5282 5950 5316
rect 5916 5192 5950 5226
rect 5916 5102 5950 5136
rect 5916 5012 5950 5046
rect 5916 4922 5950 4956
rect 5916 4832 5950 4866
rect 5916 4742 5950 4776
rect 5916 4652 5950 4686
rect 5916 4562 5950 4596
rect 5916 4472 5950 4506
rect 7103 5462 7137 5496
rect 7103 5372 7137 5406
rect 7103 5282 7137 5316
rect 7103 5192 7137 5226
rect 7103 5102 7137 5136
rect 7103 5012 7137 5046
rect 7103 4922 7137 4956
rect 7103 4832 7137 4866
rect 7103 4742 7137 4776
rect 7103 4652 7137 4686
rect 7103 4562 7137 4596
rect 7103 4472 7137 4506
rect 5939 4376 5973 4410
rect 6029 4376 6063 4410
rect 6119 4376 6153 4410
rect 6209 4376 6243 4410
rect 6299 4376 6333 4410
rect 6389 4376 6423 4410
rect 6479 4376 6513 4410
rect 6569 4376 6603 4410
rect 6659 4376 6693 4410
rect 6749 4376 6783 4410
rect 6839 4376 6873 4410
rect 6929 4376 6963 4410
rect 7019 4376 7053 4410
rect 387 4175 421 4209
rect 477 4175 511 4209
rect 567 4175 601 4209
rect 657 4175 691 4209
rect 747 4175 781 4209
rect 837 4175 871 4209
rect 927 4175 961 4209
rect 1017 4175 1051 4209
rect 1107 4175 1141 4209
rect 1197 4175 1231 4209
rect 1287 4175 1321 4209
rect 1377 4175 1411 4209
rect 1467 4175 1501 4209
rect 364 4074 398 4108
rect 364 3984 398 4018
rect 364 3894 398 3928
rect 364 3804 398 3838
rect 364 3714 398 3748
rect 364 3624 398 3658
rect 364 3534 398 3568
rect 364 3444 398 3478
rect 364 3354 398 3388
rect 364 3264 398 3298
rect 364 3174 398 3208
rect 364 3084 398 3118
rect 1551 4074 1585 4108
rect 1551 3984 1585 4018
rect 1551 3894 1585 3928
rect 1551 3804 1585 3838
rect 1551 3714 1585 3748
rect 1551 3624 1585 3658
rect 1551 3534 1585 3568
rect 1551 3444 1585 3478
rect 1551 3354 1585 3388
rect 1551 3264 1585 3298
rect 1551 3174 1585 3208
rect 1551 3084 1585 3118
rect 387 2988 421 3022
rect 477 2988 511 3022
rect 567 2988 601 3022
rect 657 2988 691 3022
rect 747 2988 781 3022
rect 837 2988 871 3022
rect 927 2988 961 3022
rect 1017 2988 1051 3022
rect 1107 2988 1141 3022
rect 1197 2988 1231 3022
rect 1287 2988 1321 3022
rect 1377 2988 1411 3022
rect 1467 2988 1501 3022
rect 1775 4175 1809 4209
rect 1865 4175 1899 4209
rect 1955 4175 1989 4209
rect 2045 4175 2079 4209
rect 2135 4175 2169 4209
rect 2225 4175 2259 4209
rect 2315 4175 2349 4209
rect 2405 4175 2439 4209
rect 2495 4175 2529 4209
rect 2585 4175 2619 4209
rect 2675 4175 2709 4209
rect 2765 4175 2799 4209
rect 2855 4175 2889 4209
rect 1752 4074 1786 4108
rect 1752 3984 1786 4018
rect 1752 3894 1786 3928
rect 1752 3804 1786 3838
rect 1752 3714 1786 3748
rect 1752 3624 1786 3658
rect 1752 3534 1786 3568
rect 1752 3444 1786 3478
rect 1752 3354 1786 3388
rect 1752 3264 1786 3298
rect 1752 3174 1786 3208
rect 1752 3084 1786 3118
rect 2939 4074 2973 4108
rect 2939 3984 2973 4018
rect 2939 3894 2973 3928
rect 2939 3804 2973 3838
rect 2939 3714 2973 3748
rect 2939 3624 2973 3658
rect 2939 3534 2973 3568
rect 2939 3444 2973 3478
rect 2939 3354 2973 3388
rect 2939 3264 2973 3298
rect 2939 3174 2973 3208
rect 2939 3084 2973 3118
rect 1775 2988 1809 3022
rect 1865 2988 1899 3022
rect 1955 2988 1989 3022
rect 2045 2988 2079 3022
rect 2135 2988 2169 3022
rect 2225 2988 2259 3022
rect 2315 2988 2349 3022
rect 2405 2988 2439 3022
rect 2495 2988 2529 3022
rect 2585 2988 2619 3022
rect 2675 2988 2709 3022
rect 2765 2988 2799 3022
rect 2855 2988 2889 3022
rect 3163 4175 3197 4209
rect 3253 4175 3287 4209
rect 3343 4175 3377 4209
rect 3433 4175 3467 4209
rect 3523 4175 3557 4209
rect 3613 4175 3647 4209
rect 3703 4175 3737 4209
rect 3793 4175 3827 4209
rect 3883 4175 3917 4209
rect 3973 4175 4007 4209
rect 4063 4175 4097 4209
rect 4153 4175 4187 4209
rect 4243 4175 4277 4209
rect 3140 4074 3174 4108
rect 3140 3984 3174 4018
rect 3140 3894 3174 3928
rect 3140 3804 3174 3838
rect 3140 3714 3174 3748
rect 3140 3624 3174 3658
rect 3140 3534 3174 3568
rect 3140 3444 3174 3478
rect 3140 3354 3174 3388
rect 3140 3264 3174 3298
rect 3140 3174 3174 3208
rect 3140 3084 3174 3118
rect 4327 4074 4361 4108
rect 4327 3984 4361 4018
rect 4327 3894 4361 3928
rect 4327 3804 4361 3838
rect 4327 3714 4361 3748
rect 4327 3624 4361 3658
rect 4327 3534 4361 3568
rect 4327 3444 4361 3478
rect 4327 3354 4361 3388
rect 4327 3264 4361 3298
rect 4327 3174 4361 3208
rect 4327 3084 4361 3118
rect 3163 2988 3197 3022
rect 3253 2988 3287 3022
rect 3343 2988 3377 3022
rect 3433 2988 3467 3022
rect 3523 2988 3557 3022
rect 3613 2988 3647 3022
rect 3703 2988 3737 3022
rect 3793 2988 3827 3022
rect 3883 2988 3917 3022
rect 3973 2988 4007 3022
rect 4063 2988 4097 3022
rect 4153 2988 4187 3022
rect 4243 2988 4277 3022
rect 4551 4175 4585 4209
rect 4641 4175 4675 4209
rect 4731 4175 4765 4209
rect 4821 4175 4855 4209
rect 4911 4175 4945 4209
rect 5001 4175 5035 4209
rect 5091 4175 5125 4209
rect 5181 4175 5215 4209
rect 5271 4175 5305 4209
rect 5361 4175 5395 4209
rect 5451 4175 5485 4209
rect 5541 4175 5575 4209
rect 5631 4175 5665 4209
rect 4528 4074 4562 4108
rect 4528 3984 4562 4018
rect 4528 3894 4562 3928
rect 4528 3804 4562 3838
rect 4528 3714 4562 3748
rect 4528 3624 4562 3658
rect 4528 3534 4562 3568
rect 4528 3444 4562 3478
rect 4528 3354 4562 3388
rect 4528 3264 4562 3298
rect 4528 3174 4562 3208
rect 4528 3084 4562 3118
rect 5715 4074 5749 4108
rect 5715 3984 5749 4018
rect 5715 3894 5749 3928
rect 5715 3804 5749 3838
rect 5715 3714 5749 3748
rect 5715 3624 5749 3658
rect 5715 3534 5749 3568
rect 5715 3444 5749 3478
rect 5715 3354 5749 3388
rect 5715 3264 5749 3298
rect 5715 3174 5749 3208
rect 5715 3084 5749 3118
rect 4551 2988 4585 3022
rect 4641 2988 4675 3022
rect 4731 2988 4765 3022
rect 4821 2988 4855 3022
rect 4911 2988 4945 3022
rect 5001 2988 5035 3022
rect 5091 2988 5125 3022
rect 5181 2988 5215 3022
rect 5271 2988 5305 3022
rect 5361 2988 5395 3022
rect 5451 2988 5485 3022
rect 5541 2988 5575 3022
rect 5631 2988 5665 3022
rect 5939 4175 5973 4209
rect 6029 4175 6063 4209
rect 6119 4175 6153 4209
rect 6209 4175 6243 4209
rect 6299 4175 6333 4209
rect 6389 4175 6423 4209
rect 6479 4175 6513 4209
rect 6569 4175 6603 4209
rect 6659 4175 6693 4209
rect 6749 4175 6783 4209
rect 6839 4175 6873 4209
rect 6929 4175 6963 4209
rect 7019 4175 7053 4209
rect 5916 4074 5950 4108
rect 5916 3984 5950 4018
rect 5916 3894 5950 3928
rect 5916 3804 5950 3838
rect 5916 3714 5950 3748
rect 5916 3624 5950 3658
rect 5916 3534 5950 3568
rect 5916 3444 5950 3478
rect 5916 3354 5950 3388
rect 5916 3264 5950 3298
rect 5916 3174 5950 3208
rect 5916 3084 5950 3118
rect 7103 4074 7137 4108
rect 7103 3984 7137 4018
rect 7103 3894 7137 3928
rect 7103 3804 7137 3838
rect 7103 3714 7137 3748
rect 7103 3624 7137 3658
rect 7103 3534 7137 3568
rect 7103 3444 7137 3478
rect 7103 3354 7137 3388
rect 7103 3264 7137 3298
rect 7103 3174 7137 3208
rect 7103 3084 7137 3118
rect 5939 2988 5973 3022
rect 6029 2988 6063 3022
rect 6119 2988 6153 3022
rect 6209 2988 6243 3022
rect 6299 2988 6333 3022
rect 6389 2988 6423 3022
rect 6479 2988 6513 3022
rect 6569 2988 6603 3022
rect 6659 2988 6693 3022
rect 6749 2988 6783 3022
rect 6839 2988 6873 3022
rect 6929 2988 6963 3022
rect 7019 2988 7053 3022
rect 387 2787 421 2821
rect 477 2787 511 2821
rect 567 2787 601 2821
rect 657 2787 691 2821
rect 747 2787 781 2821
rect 837 2787 871 2821
rect 927 2787 961 2821
rect 1017 2787 1051 2821
rect 1107 2787 1141 2821
rect 1197 2787 1231 2821
rect 1287 2787 1321 2821
rect 1377 2787 1411 2821
rect 1467 2787 1501 2821
rect 364 2686 398 2720
rect 364 2596 398 2630
rect 364 2506 398 2540
rect 364 2416 398 2450
rect 364 2326 398 2360
rect 364 2236 398 2270
rect 364 2146 398 2180
rect 364 2056 398 2090
rect 364 1966 398 2000
rect 364 1876 398 1910
rect 364 1786 398 1820
rect 364 1696 398 1730
rect 1551 2686 1585 2720
rect 1551 2596 1585 2630
rect 1551 2506 1585 2540
rect 1551 2416 1585 2450
rect 1551 2326 1585 2360
rect 1551 2236 1585 2270
rect 1551 2146 1585 2180
rect 1551 2056 1585 2090
rect 1551 1966 1585 2000
rect 1551 1876 1585 1910
rect 1551 1786 1585 1820
rect 1551 1696 1585 1730
rect 387 1600 421 1634
rect 477 1600 511 1634
rect 567 1600 601 1634
rect 657 1600 691 1634
rect 747 1600 781 1634
rect 837 1600 871 1634
rect 927 1600 961 1634
rect 1017 1600 1051 1634
rect 1107 1600 1141 1634
rect 1197 1600 1231 1634
rect 1287 1600 1321 1634
rect 1377 1600 1411 1634
rect 1467 1600 1501 1634
rect 1775 2787 1809 2821
rect 1865 2787 1899 2821
rect 1955 2787 1989 2821
rect 2045 2787 2079 2821
rect 2135 2787 2169 2821
rect 2225 2787 2259 2821
rect 2315 2787 2349 2821
rect 2405 2787 2439 2821
rect 2495 2787 2529 2821
rect 2585 2787 2619 2821
rect 2675 2787 2709 2821
rect 2765 2787 2799 2821
rect 2855 2787 2889 2821
rect 1752 2686 1786 2720
rect 1752 2596 1786 2630
rect 1752 2506 1786 2540
rect 1752 2416 1786 2450
rect 1752 2326 1786 2360
rect 1752 2236 1786 2270
rect 1752 2146 1786 2180
rect 1752 2056 1786 2090
rect 1752 1966 1786 2000
rect 1752 1876 1786 1910
rect 1752 1786 1786 1820
rect 1752 1696 1786 1730
rect 2939 2686 2973 2720
rect 2939 2596 2973 2630
rect 2939 2506 2973 2540
rect 2939 2416 2973 2450
rect 2939 2326 2973 2360
rect 2939 2236 2973 2270
rect 2939 2146 2973 2180
rect 2939 2056 2973 2090
rect 2939 1966 2973 2000
rect 2939 1876 2973 1910
rect 2939 1786 2973 1820
rect 2939 1696 2973 1730
rect 1775 1600 1809 1634
rect 1865 1600 1899 1634
rect 1955 1600 1989 1634
rect 2045 1600 2079 1634
rect 2135 1600 2169 1634
rect 2225 1600 2259 1634
rect 2315 1600 2349 1634
rect 2405 1600 2439 1634
rect 2495 1600 2529 1634
rect 2585 1600 2619 1634
rect 2675 1600 2709 1634
rect 2765 1600 2799 1634
rect 2855 1600 2889 1634
rect 3163 2787 3197 2821
rect 3253 2787 3287 2821
rect 3343 2787 3377 2821
rect 3433 2787 3467 2821
rect 3523 2787 3557 2821
rect 3613 2787 3647 2821
rect 3703 2787 3737 2821
rect 3793 2787 3827 2821
rect 3883 2787 3917 2821
rect 3973 2787 4007 2821
rect 4063 2787 4097 2821
rect 4153 2787 4187 2821
rect 4243 2787 4277 2821
rect 3140 2686 3174 2720
rect 3140 2596 3174 2630
rect 3140 2506 3174 2540
rect 3140 2416 3174 2450
rect 3140 2326 3174 2360
rect 3140 2236 3174 2270
rect 3140 2146 3174 2180
rect 3140 2056 3174 2090
rect 3140 1966 3174 2000
rect 3140 1876 3174 1910
rect 3140 1786 3174 1820
rect 3140 1696 3174 1730
rect 4327 2686 4361 2720
rect 4327 2596 4361 2630
rect 4327 2506 4361 2540
rect 4327 2416 4361 2450
rect 4327 2326 4361 2360
rect 4327 2236 4361 2270
rect 4327 2146 4361 2180
rect 4327 2056 4361 2090
rect 4327 1966 4361 2000
rect 4327 1876 4361 1910
rect 4327 1786 4361 1820
rect 4327 1696 4361 1730
rect 3163 1600 3197 1634
rect 3253 1600 3287 1634
rect 3343 1600 3377 1634
rect 3433 1600 3467 1634
rect 3523 1600 3557 1634
rect 3613 1600 3647 1634
rect 3703 1600 3737 1634
rect 3793 1600 3827 1634
rect 3883 1600 3917 1634
rect 3973 1600 4007 1634
rect 4063 1600 4097 1634
rect 4153 1600 4187 1634
rect 4243 1600 4277 1634
rect 4551 2787 4585 2821
rect 4641 2787 4675 2821
rect 4731 2787 4765 2821
rect 4821 2787 4855 2821
rect 4911 2787 4945 2821
rect 5001 2787 5035 2821
rect 5091 2787 5125 2821
rect 5181 2787 5215 2821
rect 5271 2787 5305 2821
rect 5361 2787 5395 2821
rect 5451 2787 5485 2821
rect 5541 2787 5575 2821
rect 5631 2787 5665 2821
rect 4528 2686 4562 2720
rect 4528 2596 4562 2630
rect 4528 2506 4562 2540
rect 4528 2416 4562 2450
rect 4528 2326 4562 2360
rect 4528 2236 4562 2270
rect 4528 2146 4562 2180
rect 4528 2056 4562 2090
rect 4528 1966 4562 2000
rect 4528 1876 4562 1910
rect 4528 1786 4562 1820
rect 4528 1696 4562 1730
rect 5715 2686 5749 2720
rect 5715 2596 5749 2630
rect 5715 2506 5749 2540
rect 5715 2416 5749 2450
rect 5715 2326 5749 2360
rect 5715 2236 5749 2270
rect 5715 2146 5749 2180
rect 5715 2056 5749 2090
rect 5715 1966 5749 2000
rect 5715 1876 5749 1910
rect 5715 1786 5749 1820
rect 5715 1696 5749 1730
rect 4551 1600 4585 1634
rect 4641 1600 4675 1634
rect 4731 1600 4765 1634
rect 4821 1600 4855 1634
rect 4911 1600 4945 1634
rect 5001 1600 5035 1634
rect 5091 1600 5125 1634
rect 5181 1600 5215 1634
rect 5271 1600 5305 1634
rect 5361 1600 5395 1634
rect 5451 1600 5485 1634
rect 5541 1600 5575 1634
rect 5631 1600 5665 1634
rect 5939 2787 5973 2821
rect 6029 2787 6063 2821
rect 6119 2787 6153 2821
rect 6209 2787 6243 2821
rect 6299 2787 6333 2821
rect 6389 2787 6423 2821
rect 6479 2787 6513 2821
rect 6569 2787 6603 2821
rect 6659 2787 6693 2821
rect 6749 2787 6783 2821
rect 6839 2787 6873 2821
rect 6929 2787 6963 2821
rect 7019 2787 7053 2821
rect 5916 2686 5950 2720
rect 5916 2596 5950 2630
rect 5916 2506 5950 2540
rect 5916 2416 5950 2450
rect 5916 2326 5950 2360
rect 5916 2236 5950 2270
rect 5916 2146 5950 2180
rect 5916 2056 5950 2090
rect 5916 1966 5950 2000
rect 5916 1876 5950 1910
rect 5916 1786 5950 1820
rect 5916 1696 5950 1730
rect 7103 2686 7137 2720
rect 7103 2596 7137 2630
rect 7103 2506 7137 2540
rect 7103 2416 7137 2450
rect 7103 2326 7137 2360
rect 7103 2236 7137 2270
rect 7103 2146 7137 2180
rect 7103 2056 7137 2090
rect 7103 1966 7137 2000
rect 7103 1876 7137 1910
rect 7103 1786 7137 1820
rect 7103 1696 7137 1730
rect 5939 1600 5973 1634
rect 6029 1600 6063 1634
rect 6119 1600 6153 1634
rect 6209 1600 6243 1634
rect 6299 1600 6333 1634
rect 6389 1600 6423 1634
rect 6479 1600 6513 1634
rect 6569 1600 6603 1634
rect 6659 1600 6693 1634
rect 6749 1600 6783 1634
rect 6839 1600 6873 1634
rect 6929 1600 6963 1634
rect 7019 1600 7053 1634
<< nsubdiffcont >>
rect -17877 22967 9141 23001
rect -17937 -375 -17903 22941
rect -16606 17607 -7986 17641
rect -16699 15724 -16665 17581
rect -7935 15724 -7901 17581
rect -16606 15664 -7986 15698
rect -7585 17518 -3081 17552
rect -7670 15718 -7636 17492
rect -3030 15718 -2996 17492
rect -7585 15658 -3081 15692
rect -12423 15558 -7986 15592
rect -12483 14722 -12449 15532
rect -7960 14722 -7926 15532
rect -7502 15543 -3096 15577
rect -7562 14785 -7528 15517
rect -3070 14785 -3036 15517
rect -7502 14725 -3096 14759
rect -12423 14662 -7986 14696
rect 367 12555 6341 12589
rect 307 10033 341 12529
rect 4896 11878 6076 11912
rect 4836 10646 4870 11852
rect 6102 10646 6136 11852
rect 4896 10586 6076 10620
rect 6367 10033 6401 12529
rect 367 9973 6341 10007
rect 587 8190 621 8224
rect 677 8190 711 8224
rect 767 8190 801 8224
rect 857 8190 891 8224
rect 947 8190 981 8224
rect 1037 8190 1071 8224
rect 1127 8190 1161 8224
rect 1217 8190 1251 8224
rect 1307 8190 1341 8224
rect 511 8132 545 8166
rect 511 8042 545 8076
rect 511 7952 545 7986
rect 511 7862 545 7896
rect 511 7772 545 7806
rect 511 7682 545 7716
rect 511 7592 545 7626
rect 511 7502 545 7536
rect 511 7412 545 7446
rect 1401 8098 1435 8132
rect 1401 8008 1435 8042
rect 1401 7918 1435 7952
rect 1401 7828 1435 7862
rect 1401 7738 1435 7772
rect 1401 7648 1435 7682
rect 1401 7558 1435 7592
rect 1401 7468 1435 7502
rect 1401 7378 1435 7412
rect 568 7300 602 7334
rect 658 7300 692 7334
rect 748 7300 782 7334
rect 838 7300 872 7334
rect 928 7300 962 7334
rect 1018 7300 1052 7334
rect 1108 7300 1142 7334
rect 1198 7300 1232 7334
rect 1288 7300 1322 7334
rect 1975 8190 2009 8224
rect 2065 8190 2099 8224
rect 2155 8190 2189 8224
rect 2245 8190 2279 8224
rect 2335 8190 2369 8224
rect 2425 8190 2459 8224
rect 2515 8190 2549 8224
rect 2605 8190 2639 8224
rect 2695 8190 2729 8224
rect 1899 8132 1933 8166
rect 1899 8042 1933 8076
rect 1899 7952 1933 7986
rect 1899 7862 1933 7896
rect 1899 7772 1933 7806
rect 1899 7682 1933 7716
rect 1899 7592 1933 7626
rect 1899 7502 1933 7536
rect 1899 7412 1933 7446
rect 2789 8098 2823 8132
rect 2789 8008 2823 8042
rect 2789 7918 2823 7952
rect 2789 7828 2823 7862
rect 2789 7738 2823 7772
rect 2789 7648 2823 7682
rect 2789 7558 2823 7592
rect 2789 7468 2823 7502
rect 2789 7378 2823 7412
rect 1956 7300 1990 7334
rect 2046 7300 2080 7334
rect 2136 7300 2170 7334
rect 2226 7300 2260 7334
rect 2316 7300 2350 7334
rect 2406 7300 2440 7334
rect 2496 7300 2530 7334
rect 2586 7300 2620 7334
rect 2676 7300 2710 7334
rect 3363 8190 3397 8224
rect 3453 8190 3487 8224
rect 3543 8190 3577 8224
rect 3633 8190 3667 8224
rect 3723 8190 3757 8224
rect 3813 8190 3847 8224
rect 3903 8190 3937 8224
rect 3993 8190 4027 8224
rect 4083 8190 4117 8224
rect 3287 8132 3321 8166
rect 3287 8042 3321 8076
rect 3287 7952 3321 7986
rect 3287 7862 3321 7896
rect 3287 7772 3321 7806
rect 3287 7682 3321 7716
rect 3287 7592 3321 7626
rect 3287 7502 3321 7536
rect 3287 7412 3321 7446
rect 4177 8098 4211 8132
rect 4177 8008 4211 8042
rect 4177 7918 4211 7952
rect 4177 7828 4211 7862
rect 4177 7738 4211 7772
rect 4177 7648 4211 7682
rect 4177 7558 4211 7592
rect 4177 7468 4211 7502
rect 4177 7378 4211 7412
rect 3344 7300 3378 7334
rect 3434 7300 3468 7334
rect 3524 7300 3558 7334
rect 3614 7300 3648 7334
rect 3704 7300 3738 7334
rect 3794 7300 3828 7334
rect 3884 7300 3918 7334
rect 3974 7300 4008 7334
rect 4064 7300 4098 7334
rect 4751 8190 4785 8224
rect 4841 8190 4875 8224
rect 4931 8190 4965 8224
rect 5021 8190 5055 8224
rect 5111 8190 5145 8224
rect 5201 8190 5235 8224
rect 5291 8190 5325 8224
rect 5381 8190 5415 8224
rect 5471 8190 5505 8224
rect 4675 8132 4709 8166
rect 4675 8042 4709 8076
rect 4675 7952 4709 7986
rect 4675 7862 4709 7896
rect 4675 7772 4709 7806
rect 4675 7682 4709 7716
rect 4675 7592 4709 7626
rect 4675 7502 4709 7536
rect 4675 7412 4709 7446
rect 5565 8098 5599 8132
rect 5565 8008 5599 8042
rect 5565 7918 5599 7952
rect 5565 7828 5599 7862
rect 5565 7738 5599 7772
rect 5565 7648 5599 7682
rect 5565 7558 5599 7592
rect 5565 7468 5599 7502
rect 5565 7378 5599 7412
rect 4732 7300 4766 7334
rect 4822 7300 4856 7334
rect 4912 7300 4946 7334
rect 5002 7300 5036 7334
rect 5092 7300 5126 7334
rect 5182 7300 5216 7334
rect 5272 7300 5306 7334
rect 5362 7300 5396 7334
rect 5452 7300 5486 7334
rect 6139 8190 6173 8224
rect 6229 8190 6263 8224
rect 6319 8190 6353 8224
rect 6409 8190 6443 8224
rect 6499 8190 6533 8224
rect 6589 8190 6623 8224
rect 6679 8190 6713 8224
rect 6769 8190 6803 8224
rect 6859 8190 6893 8224
rect 6063 8132 6097 8166
rect 6063 8042 6097 8076
rect 6063 7952 6097 7986
rect 6063 7862 6097 7896
rect 6063 7772 6097 7806
rect 6063 7682 6097 7716
rect 6063 7592 6097 7626
rect 6063 7502 6097 7536
rect 6063 7412 6097 7446
rect 6953 8098 6987 8132
rect 6953 8008 6987 8042
rect 6953 7918 6987 7952
rect 6953 7828 6987 7862
rect 6953 7738 6987 7772
rect 6953 7648 6987 7682
rect 6953 7558 6987 7592
rect 6953 7468 6987 7502
rect 6953 7378 6987 7412
rect 6120 7300 6154 7334
rect 6210 7300 6244 7334
rect 6300 7300 6334 7334
rect 6390 7300 6424 7334
rect 6480 7300 6514 7334
rect 6570 7300 6604 7334
rect 6660 7300 6694 7334
rect 6750 7300 6784 7334
rect 6840 7300 6874 7334
rect 587 6802 621 6836
rect 677 6802 711 6836
rect 767 6802 801 6836
rect 857 6802 891 6836
rect 947 6802 981 6836
rect 1037 6802 1071 6836
rect 1127 6802 1161 6836
rect 1217 6802 1251 6836
rect 1307 6802 1341 6836
rect 511 6744 545 6778
rect 511 6654 545 6688
rect 511 6564 545 6598
rect 511 6474 545 6508
rect 511 6384 545 6418
rect 511 6294 545 6328
rect 511 6204 545 6238
rect 511 6114 545 6148
rect 511 6024 545 6058
rect 1401 6710 1435 6744
rect 1401 6620 1435 6654
rect 1401 6530 1435 6564
rect 1401 6440 1435 6474
rect 1401 6350 1435 6384
rect 1401 6260 1435 6294
rect 1401 6170 1435 6204
rect 1401 6080 1435 6114
rect 1401 5990 1435 6024
rect 568 5912 602 5946
rect 658 5912 692 5946
rect 748 5912 782 5946
rect 838 5912 872 5946
rect 928 5912 962 5946
rect 1018 5912 1052 5946
rect 1108 5912 1142 5946
rect 1198 5912 1232 5946
rect 1288 5912 1322 5946
rect 1975 6802 2009 6836
rect 2065 6802 2099 6836
rect 2155 6802 2189 6836
rect 2245 6802 2279 6836
rect 2335 6802 2369 6836
rect 2425 6802 2459 6836
rect 2515 6802 2549 6836
rect 2605 6802 2639 6836
rect 2695 6802 2729 6836
rect 1899 6744 1933 6778
rect 1899 6654 1933 6688
rect 1899 6564 1933 6598
rect 1899 6474 1933 6508
rect 1899 6384 1933 6418
rect 1899 6294 1933 6328
rect 1899 6204 1933 6238
rect 1899 6114 1933 6148
rect 1899 6024 1933 6058
rect 2789 6710 2823 6744
rect 2789 6620 2823 6654
rect 2789 6530 2823 6564
rect 2789 6440 2823 6474
rect 2789 6350 2823 6384
rect 2789 6260 2823 6294
rect 2789 6170 2823 6204
rect 2789 6080 2823 6114
rect 2789 5990 2823 6024
rect 1956 5912 1990 5946
rect 2046 5912 2080 5946
rect 2136 5912 2170 5946
rect 2226 5912 2260 5946
rect 2316 5912 2350 5946
rect 2406 5912 2440 5946
rect 2496 5912 2530 5946
rect 2586 5912 2620 5946
rect 2676 5912 2710 5946
rect 3363 6802 3397 6836
rect 3453 6802 3487 6836
rect 3543 6802 3577 6836
rect 3633 6802 3667 6836
rect 3723 6802 3757 6836
rect 3813 6802 3847 6836
rect 3903 6802 3937 6836
rect 3993 6802 4027 6836
rect 4083 6802 4117 6836
rect 3287 6744 3321 6778
rect 3287 6654 3321 6688
rect 3287 6564 3321 6598
rect 3287 6474 3321 6508
rect 3287 6384 3321 6418
rect 3287 6294 3321 6328
rect 3287 6204 3321 6238
rect 3287 6114 3321 6148
rect 3287 6024 3321 6058
rect 4177 6710 4211 6744
rect 4177 6620 4211 6654
rect 4177 6530 4211 6564
rect 4177 6440 4211 6474
rect 4177 6350 4211 6384
rect 4177 6260 4211 6294
rect 4177 6170 4211 6204
rect 4177 6080 4211 6114
rect 4177 5990 4211 6024
rect 3344 5912 3378 5946
rect 3434 5912 3468 5946
rect 3524 5912 3558 5946
rect 3614 5912 3648 5946
rect 3704 5912 3738 5946
rect 3794 5912 3828 5946
rect 3884 5912 3918 5946
rect 3974 5912 4008 5946
rect 4064 5912 4098 5946
rect 4751 6802 4785 6836
rect 4841 6802 4875 6836
rect 4931 6802 4965 6836
rect 5021 6802 5055 6836
rect 5111 6802 5145 6836
rect 5201 6802 5235 6836
rect 5291 6802 5325 6836
rect 5381 6802 5415 6836
rect 5471 6802 5505 6836
rect 4675 6744 4709 6778
rect 4675 6654 4709 6688
rect 4675 6564 4709 6598
rect 4675 6474 4709 6508
rect 4675 6384 4709 6418
rect 4675 6294 4709 6328
rect 4675 6204 4709 6238
rect 4675 6114 4709 6148
rect 4675 6024 4709 6058
rect 5565 6710 5599 6744
rect 5565 6620 5599 6654
rect 5565 6530 5599 6564
rect 5565 6440 5599 6474
rect 5565 6350 5599 6384
rect 5565 6260 5599 6294
rect 5565 6170 5599 6204
rect 5565 6080 5599 6114
rect 5565 5990 5599 6024
rect 4732 5912 4766 5946
rect 4822 5912 4856 5946
rect 4912 5912 4946 5946
rect 5002 5912 5036 5946
rect 5092 5912 5126 5946
rect 5182 5912 5216 5946
rect 5272 5912 5306 5946
rect 5362 5912 5396 5946
rect 5452 5912 5486 5946
rect 6139 6802 6173 6836
rect 6229 6802 6263 6836
rect 6319 6802 6353 6836
rect 6409 6802 6443 6836
rect 6499 6802 6533 6836
rect 6589 6802 6623 6836
rect 6679 6802 6713 6836
rect 6769 6802 6803 6836
rect 6859 6802 6893 6836
rect 6063 6744 6097 6778
rect 6063 6654 6097 6688
rect 6063 6564 6097 6598
rect 6063 6474 6097 6508
rect 6063 6384 6097 6418
rect 6063 6294 6097 6328
rect 6063 6204 6097 6238
rect 6063 6114 6097 6148
rect 6063 6024 6097 6058
rect 6953 6710 6987 6744
rect 6953 6620 6987 6654
rect 6953 6530 6987 6564
rect 6953 6440 6987 6474
rect 6953 6350 6987 6384
rect 6953 6260 6987 6294
rect 6953 6170 6987 6204
rect 6953 6080 6987 6114
rect 6953 5990 6987 6024
rect 6120 5912 6154 5946
rect 6210 5912 6244 5946
rect 6300 5912 6334 5946
rect 6390 5912 6424 5946
rect 6480 5912 6514 5946
rect 6570 5912 6604 5946
rect 6660 5912 6694 5946
rect 6750 5912 6784 5946
rect 6840 5912 6874 5946
rect 587 5414 621 5448
rect 677 5414 711 5448
rect 767 5414 801 5448
rect 857 5414 891 5448
rect 947 5414 981 5448
rect 1037 5414 1071 5448
rect 1127 5414 1161 5448
rect 1217 5414 1251 5448
rect 1307 5414 1341 5448
rect 511 5356 545 5390
rect 511 5266 545 5300
rect 511 5176 545 5210
rect 511 5086 545 5120
rect 511 4996 545 5030
rect 511 4906 545 4940
rect 511 4816 545 4850
rect 511 4726 545 4760
rect 511 4636 545 4670
rect 1401 5322 1435 5356
rect 1401 5232 1435 5266
rect 1401 5142 1435 5176
rect 1401 5052 1435 5086
rect 1401 4962 1435 4996
rect 1401 4872 1435 4906
rect 1401 4782 1435 4816
rect 1401 4692 1435 4726
rect 1401 4602 1435 4636
rect 568 4524 602 4558
rect 658 4524 692 4558
rect 748 4524 782 4558
rect 838 4524 872 4558
rect 928 4524 962 4558
rect 1018 4524 1052 4558
rect 1108 4524 1142 4558
rect 1198 4524 1232 4558
rect 1288 4524 1322 4558
rect 1975 5414 2009 5448
rect 2065 5414 2099 5448
rect 2155 5414 2189 5448
rect 2245 5414 2279 5448
rect 2335 5414 2369 5448
rect 2425 5414 2459 5448
rect 2515 5414 2549 5448
rect 2605 5414 2639 5448
rect 2695 5414 2729 5448
rect 1899 5356 1933 5390
rect 1899 5266 1933 5300
rect 1899 5176 1933 5210
rect 1899 5086 1933 5120
rect 1899 4996 1933 5030
rect 1899 4906 1933 4940
rect 1899 4816 1933 4850
rect 1899 4726 1933 4760
rect 1899 4636 1933 4670
rect 2789 5322 2823 5356
rect 2789 5232 2823 5266
rect 2789 5142 2823 5176
rect 2789 5052 2823 5086
rect 2789 4962 2823 4996
rect 2789 4872 2823 4906
rect 2789 4782 2823 4816
rect 2789 4692 2823 4726
rect 2789 4602 2823 4636
rect 1956 4524 1990 4558
rect 2046 4524 2080 4558
rect 2136 4524 2170 4558
rect 2226 4524 2260 4558
rect 2316 4524 2350 4558
rect 2406 4524 2440 4558
rect 2496 4524 2530 4558
rect 2586 4524 2620 4558
rect 2676 4524 2710 4558
rect 3363 5414 3397 5448
rect 3453 5414 3487 5448
rect 3543 5414 3577 5448
rect 3633 5414 3667 5448
rect 3723 5414 3757 5448
rect 3813 5414 3847 5448
rect 3903 5414 3937 5448
rect 3993 5414 4027 5448
rect 4083 5414 4117 5448
rect 3287 5356 3321 5390
rect 3287 5266 3321 5300
rect 3287 5176 3321 5210
rect 3287 5086 3321 5120
rect 3287 4996 3321 5030
rect 3287 4906 3321 4940
rect 3287 4816 3321 4850
rect 3287 4726 3321 4760
rect 3287 4636 3321 4670
rect 4177 5322 4211 5356
rect 4177 5232 4211 5266
rect 4177 5142 4211 5176
rect 4177 5052 4211 5086
rect 4177 4962 4211 4996
rect 4177 4872 4211 4906
rect 4177 4782 4211 4816
rect 4177 4692 4211 4726
rect 4177 4602 4211 4636
rect 3344 4524 3378 4558
rect 3434 4524 3468 4558
rect 3524 4524 3558 4558
rect 3614 4524 3648 4558
rect 3704 4524 3738 4558
rect 3794 4524 3828 4558
rect 3884 4524 3918 4558
rect 3974 4524 4008 4558
rect 4064 4524 4098 4558
rect 4751 5414 4785 5448
rect 4841 5414 4875 5448
rect 4931 5414 4965 5448
rect 5021 5414 5055 5448
rect 5111 5414 5145 5448
rect 5201 5414 5235 5448
rect 5291 5414 5325 5448
rect 5381 5414 5415 5448
rect 5471 5414 5505 5448
rect 4675 5356 4709 5390
rect 4675 5266 4709 5300
rect 4675 5176 4709 5210
rect 4675 5086 4709 5120
rect 4675 4996 4709 5030
rect 4675 4906 4709 4940
rect 4675 4816 4709 4850
rect 4675 4726 4709 4760
rect 4675 4636 4709 4670
rect 5565 5322 5599 5356
rect 5565 5232 5599 5266
rect 5565 5142 5599 5176
rect 5565 5052 5599 5086
rect 5565 4962 5599 4996
rect 5565 4872 5599 4906
rect 5565 4782 5599 4816
rect 5565 4692 5599 4726
rect 5565 4602 5599 4636
rect 4732 4524 4766 4558
rect 4822 4524 4856 4558
rect 4912 4524 4946 4558
rect 5002 4524 5036 4558
rect 5092 4524 5126 4558
rect 5182 4524 5216 4558
rect 5272 4524 5306 4558
rect 5362 4524 5396 4558
rect 5452 4524 5486 4558
rect 6139 5414 6173 5448
rect 6229 5414 6263 5448
rect 6319 5414 6353 5448
rect 6409 5414 6443 5448
rect 6499 5414 6533 5448
rect 6589 5414 6623 5448
rect 6679 5414 6713 5448
rect 6769 5414 6803 5448
rect 6859 5414 6893 5448
rect 6063 5356 6097 5390
rect 6063 5266 6097 5300
rect 6063 5176 6097 5210
rect 6063 5086 6097 5120
rect 6063 4996 6097 5030
rect 6063 4906 6097 4940
rect 6063 4816 6097 4850
rect 6063 4726 6097 4760
rect 6063 4636 6097 4670
rect 6953 5322 6987 5356
rect 6953 5232 6987 5266
rect 6953 5142 6987 5176
rect 6953 5052 6987 5086
rect 6953 4962 6987 4996
rect 6953 4872 6987 4906
rect 6953 4782 6987 4816
rect 6953 4692 6987 4726
rect 6953 4602 6987 4636
rect 6120 4524 6154 4558
rect 6210 4524 6244 4558
rect 6300 4524 6334 4558
rect 6390 4524 6424 4558
rect 6480 4524 6514 4558
rect 6570 4524 6604 4558
rect 6660 4524 6694 4558
rect 6750 4524 6784 4558
rect 6840 4524 6874 4558
rect 587 4026 621 4060
rect 677 4026 711 4060
rect 767 4026 801 4060
rect 857 4026 891 4060
rect 947 4026 981 4060
rect 1037 4026 1071 4060
rect 1127 4026 1161 4060
rect 1217 4026 1251 4060
rect 1307 4026 1341 4060
rect 511 3968 545 4002
rect 511 3878 545 3912
rect 511 3788 545 3822
rect 511 3698 545 3732
rect 511 3608 545 3642
rect 511 3518 545 3552
rect 511 3428 545 3462
rect 511 3338 545 3372
rect 511 3248 545 3282
rect 1401 3934 1435 3968
rect 1401 3844 1435 3878
rect 1401 3754 1435 3788
rect 1401 3664 1435 3698
rect 1401 3574 1435 3608
rect 1401 3484 1435 3518
rect 1401 3394 1435 3428
rect 1401 3304 1435 3338
rect 1401 3214 1435 3248
rect 568 3136 602 3170
rect 658 3136 692 3170
rect 748 3136 782 3170
rect 838 3136 872 3170
rect 928 3136 962 3170
rect 1018 3136 1052 3170
rect 1108 3136 1142 3170
rect 1198 3136 1232 3170
rect 1288 3136 1322 3170
rect 1975 4026 2009 4060
rect 2065 4026 2099 4060
rect 2155 4026 2189 4060
rect 2245 4026 2279 4060
rect 2335 4026 2369 4060
rect 2425 4026 2459 4060
rect 2515 4026 2549 4060
rect 2605 4026 2639 4060
rect 2695 4026 2729 4060
rect 1899 3968 1933 4002
rect 1899 3878 1933 3912
rect 1899 3788 1933 3822
rect 1899 3698 1933 3732
rect 1899 3608 1933 3642
rect 1899 3518 1933 3552
rect 1899 3428 1933 3462
rect 1899 3338 1933 3372
rect 1899 3248 1933 3282
rect 2789 3934 2823 3968
rect 2789 3844 2823 3878
rect 2789 3754 2823 3788
rect 2789 3664 2823 3698
rect 2789 3574 2823 3608
rect 2789 3484 2823 3518
rect 2789 3394 2823 3428
rect 2789 3304 2823 3338
rect 2789 3214 2823 3248
rect 1956 3136 1990 3170
rect 2046 3136 2080 3170
rect 2136 3136 2170 3170
rect 2226 3136 2260 3170
rect 2316 3136 2350 3170
rect 2406 3136 2440 3170
rect 2496 3136 2530 3170
rect 2586 3136 2620 3170
rect 2676 3136 2710 3170
rect 3363 4026 3397 4060
rect 3453 4026 3487 4060
rect 3543 4026 3577 4060
rect 3633 4026 3667 4060
rect 3723 4026 3757 4060
rect 3813 4026 3847 4060
rect 3903 4026 3937 4060
rect 3993 4026 4027 4060
rect 4083 4026 4117 4060
rect 3287 3968 3321 4002
rect 3287 3878 3321 3912
rect 3287 3788 3321 3822
rect 3287 3698 3321 3732
rect 3287 3608 3321 3642
rect 3287 3518 3321 3552
rect 3287 3428 3321 3462
rect 3287 3338 3321 3372
rect 3287 3248 3321 3282
rect 4177 3934 4211 3968
rect 4177 3844 4211 3878
rect 4177 3754 4211 3788
rect 4177 3664 4211 3698
rect 4177 3574 4211 3608
rect 4177 3484 4211 3518
rect 4177 3394 4211 3428
rect 4177 3304 4211 3338
rect 4177 3214 4211 3248
rect 3344 3136 3378 3170
rect 3434 3136 3468 3170
rect 3524 3136 3558 3170
rect 3614 3136 3648 3170
rect 3704 3136 3738 3170
rect 3794 3136 3828 3170
rect 3884 3136 3918 3170
rect 3974 3136 4008 3170
rect 4064 3136 4098 3170
rect 4751 4026 4785 4060
rect 4841 4026 4875 4060
rect 4931 4026 4965 4060
rect 5021 4026 5055 4060
rect 5111 4026 5145 4060
rect 5201 4026 5235 4060
rect 5291 4026 5325 4060
rect 5381 4026 5415 4060
rect 5471 4026 5505 4060
rect 4675 3968 4709 4002
rect 4675 3878 4709 3912
rect 4675 3788 4709 3822
rect 4675 3698 4709 3732
rect 4675 3608 4709 3642
rect 4675 3518 4709 3552
rect 4675 3428 4709 3462
rect 4675 3338 4709 3372
rect 4675 3248 4709 3282
rect 5565 3934 5599 3968
rect 5565 3844 5599 3878
rect 5565 3754 5599 3788
rect 5565 3664 5599 3698
rect 5565 3574 5599 3608
rect 5565 3484 5599 3518
rect 5565 3394 5599 3428
rect 5565 3304 5599 3338
rect 5565 3214 5599 3248
rect 4732 3136 4766 3170
rect 4822 3136 4856 3170
rect 4912 3136 4946 3170
rect 5002 3136 5036 3170
rect 5092 3136 5126 3170
rect 5182 3136 5216 3170
rect 5272 3136 5306 3170
rect 5362 3136 5396 3170
rect 5452 3136 5486 3170
rect 6139 4026 6173 4060
rect 6229 4026 6263 4060
rect 6319 4026 6353 4060
rect 6409 4026 6443 4060
rect 6499 4026 6533 4060
rect 6589 4026 6623 4060
rect 6679 4026 6713 4060
rect 6769 4026 6803 4060
rect 6859 4026 6893 4060
rect 6063 3968 6097 4002
rect 6063 3878 6097 3912
rect 6063 3788 6097 3822
rect 6063 3698 6097 3732
rect 6063 3608 6097 3642
rect 6063 3518 6097 3552
rect 6063 3428 6097 3462
rect 6063 3338 6097 3372
rect 6063 3248 6097 3282
rect 6953 3934 6987 3968
rect 6953 3844 6987 3878
rect 6953 3754 6987 3788
rect 6953 3664 6987 3698
rect 6953 3574 6987 3608
rect 6953 3484 6987 3518
rect 6953 3394 6987 3428
rect 6953 3304 6987 3338
rect 6953 3214 6987 3248
rect 6120 3136 6154 3170
rect 6210 3136 6244 3170
rect 6300 3136 6334 3170
rect 6390 3136 6424 3170
rect 6480 3136 6514 3170
rect 6570 3136 6604 3170
rect 6660 3136 6694 3170
rect 6750 3136 6784 3170
rect 6840 3136 6874 3170
rect 587 2638 621 2672
rect 677 2638 711 2672
rect 767 2638 801 2672
rect 857 2638 891 2672
rect 947 2638 981 2672
rect 1037 2638 1071 2672
rect 1127 2638 1161 2672
rect 1217 2638 1251 2672
rect 1307 2638 1341 2672
rect 511 2580 545 2614
rect 511 2490 545 2524
rect 511 2400 545 2434
rect 511 2310 545 2344
rect 511 2220 545 2254
rect 511 2130 545 2164
rect 511 2040 545 2074
rect 511 1950 545 1984
rect 511 1860 545 1894
rect 1401 2546 1435 2580
rect 1401 2456 1435 2490
rect 1401 2366 1435 2400
rect 1401 2276 1435 2310
rect 1401 2186 1435 2220
rect 1401 2096 1435 2130
rect 1401 2006 1435 2040
rect 1401 1916 1435 1950
rect 1401 1826 1435 1860
rect 568 1748 602 1782
rect 658 1748 692 1782
rect 748 1748 782 1782
rect 838 1748 872 1782
rect 928 1748 962 1782
rect 1018 1748 1052 1782
rect 1108 1748 1142 1782
rect 1198 1748 1232 1782
rect 1288 1748 1322 1782
rect 1975 2638 2009 2672
rect 2065 2638 2099 2672
rect 2155 2638 2189 2672
rect 2245 2638 2279 2672
rect 2335 2638 2369 2672
rect 2425 2638 2459 2672
rect 2515 2638 2549 2672
rect 2605 2638 2639 2672
rect 2695 2638 2729 2672
rect 1899 2580 1933 2614
rect 1899 2490 1933 2524
rect 1899 2400 1933 2434
rect 1899 2310 1933 2344
rect 1899 2220 1933 2254
rect 1899 2130 1933 2164
rect 1899 2040 1933 2074
rect 1899 1950 1933 1984
rect 1899 1860 1933 1894
rect 2789 2546 2823 2580
rect 2789 2456 2823 2490
rect 2789 2366 2823 2400
rect 2789 2276 2823 2310
rect 2789 2186 2823 2220
rect 2789 2096 2823 2130
rect 2789 2006 2823 2040
rect 2789 1916 2823 1950
rect 2789 1826 2823 1860
rect 1956 1748 1990 1782
rect 2046 1748 2080 1782
rect 2136 1748 2170 1782
rect 2226 1748 2260 1782
rect 2316 1748 2350 1782
rect 2406 1748 2440 1782
rect 2496 1748 2530 1782
rect 2586 1748 2620 1782
rect 2676 1748 2710 1782
rect 3363 2638 3397 2672
rect 3453 2638 3487 2672
rect 3543 2638 3577 2672
rect 3633 2638 3667 2672
rect 3723 2638 3757 2672
rect 3813 2638 3847 2672
rect 3903 2638 3937 2672
rect 3993 2638 4027 2672
rect 4083 2638 4117 2672
rect 3287 2580 3321 2614
rect 3287 2490 3321 2524
rect 3287 2400 3321 2434
rect 3287 2310 3321 2344
rect 3287 2220 3321 2254
rect 3287 2130 3321 2164
rect 3287 2040 3321 2074
rect 3287 1950 3321 1984
rect 3287 1860 3321 1894
rect 4177 2546 4211 2580
rect 4177 2456 4211 2490
rect 4177 2366 4211 2400
rect 4177 2276 4211 2310
rect 4177 2186 4211 2220
rect 4177 2096 4211 2130
rect 4177 2006 4211 2040
rect 4177 1916 4211 1950
rect 4177 1826 4211 1860
rect 3344 1748 3378 1782
rect 3434 1748 3468 1782
rect 3524 1748 3558 1782
rect 3614 1748 3648 1782
rect 3704 1748 3738 1782
rect 3794 1748 3828 1782
rect 3884 1748 3918 1782
rect 3974 1748 4008 1782
rect 4064 1748 4098 1782
rect 4751 2638 4785 2672
rect 4841 2638 4875 2672
rect 4931 2638 4965 2672
rect 5021 2638 5055 2672
rect 5111 2638 5145 2672
rect 5201 2638 5235 2672
rect 5291 2638 5325 2672
rect 5381 2638 5415 2672
rect 5471 2638 5505 2672
rect 4675 2580 4709 2614
rect 4675 2490 4709 2524
rect 4675 2400 4709 2434
rect 4675 2310 4709 2344
rect 4675 2220 4709 2254
rect 4675 2130 4709 2164
rect 4675 2040 4709 2074
rect 4675 1950 4709 1984
rect 4675 1860 4709 1894
rect 5565 2546 5599 2580
rect 5565 2456 5599 2490
rect 5565 2366 5599 2400
rect 5565 2276 5599 2310
rect 5565 2186 5599 2220
rect 5565 2096 5599 2130
rect 5565 2006 5599 2040
rect 5565 1916 5599 1950
rect 5565 1826 5599 1860
rect 4732 1748 4766 1782
rect 4822 1748 4856 1782
rect 4912 1748 4946 1782
rect 5002 1748 5036 1782
rect 5092 1748 5126 1782
rect 5182 1748 5216 1782
rect 5272 1748 5306 1782
rect 5362 1748 5396 1782
rect 5452 1748 5486 1782
rect 6139 2638 6173 2672
rect 6229 2638 6263 2672
rect 6319 2638 6353 2672
rect 6409 2638 6443 2672
rect 6499 2638 6533 2672
rect 6589 2638 6623 2672
rect 6679 2638 6713 2672
rect 6769 2638 6803 2672
rect 6859 2638 6893 2672
rect 6063 2580 6097 2614
rect 6063 2490 6097 2524
rect 6063 2400 6097 2434
rect 6063 2310 6097 2344
rect 6063 2220 6097 2254
rect 6063 2130 6097 2164
rect 6063 2040 6097 2074
rect 6063 1950 6097 1984
rect 6063 1860 6097 1894
rect 6953 2546 6987 2580
rect 6953 2456 6987 2490
rect 6953 2366 6987 2400
rect 6953 2276 6987 2310
rect 6953 2186 6987 2220
rect 6953 2096 6987 2130
rect 6953 2006 6987 2040
rect 6953 1916 6987 1950
rect 6953 1826 6987 1860
rect 6120 1748 6154 1782
rect 6210 1748 6244 1782
rect 6300 1748 6334 1782
rect 6390 1748 6424 1782
rect 6480 1748 6514 1782
rect 6570 1748 6604 1782
rect 6660 1748 6694 1782
rect 6750 1748 6784 1782
rect 6840 1748 6874 1782
rect 9167 -375 9201 22941
rect -17877 -435 9141 -401
<< poly >>
rect -16533 17547 -16441 17563
rect -16533 17513 -16517 17547
rect -16483 17513 -16441 17547
rect -16533 17497 -16441 17513
rect -16471 17466 -16441 17497
rect -8151 17547 -8059 17563
rect -8151 17513 -8109 17547
rect -8075 17513 -8059 17547
rect -8151 17497 -8059 17513
rect -16383 17466 -14383 17492
rect -14325 17466 -12325 17492
rect -12267 17466 -10267 17492
rect -10209 17466 -8209 17492
rect -8151 17466 -8121 17497
rect -16471 17240 -16441 17266
rect -16383 17219 -14383 17266
rect -16383 17202 -15875 17219
rect -15891 17185 -15875 17202
rect -14891 17202 -14383 17219
rect -14325 17219 -12325 17266
rect -14325 17202 -13817 17219
rect -14891 17185 -14875 17202
rect -15891 17169 -14875 17185
rect -13833 17185 -13817 17202
rect -12833 17202 -12325 17219
rect -12267 17219 -10267 17266
rect -12267 17202 -11759 17219
rect -12833 17185 -12817 17202
rect -13833 17169 -12817 17185
rect -11775 17185 -11759 17202
rect -10775 17202 -10267 17219
rect -10209 17219 -8209 17266
rect -8151 17240 -8121 17266
rect -10209 17202 -9701 17219
rect -10775 17185 -10759 17202
rect -11775 17169 -10759 17185
rect -9717 17185 -9701 17202
rect -8717 17202 -8209 17219
rect -8717 17185 -8701 17202
rect -9717 17169 -8701 17185
rect -15891 17068 -14875 17084
rect -15891 17051 -15875 17068
rect -16383 17034 -15875 17051
rect -14891 17051 -14875 17068
rect -13833 17068 -12817 17084
rect -13833 17051 -13817 17068
rect -14891 17034 -14383 17051
rect -16471 16987 -16441 17013
rect -16383 16987 -14383 17034
rect -14325 17034 -13817 17051
rect -12833 17051 -12817 17068
rect -11775 17068 -10759 17084
rect -11775 17051 -11759 17068
rect -12833 17034 -12325 17051
rect -14325 16987 -12325 17034
rect -12267 17034 -11759 17051
rect -10775 17051 -10759 17068
rect -9717 17068 -8701 17084
rect -9717 17051 -9701 17068
rect -10775 17034 -10267 17051
rect -12267 16987 -10267 17034
rect -10209 17034 -9701 17051
rect -8717 17051 -8701 17068
rect -8717 17034 -8209 17051
rect -10209 16987 -8209 17034
rect -8151 16987 -8121 17013
rect -16471 16685 -16441 16787
rect -16533 16669 -16441 16685
rect -16533 16635 -16517 16669
rect -16483 16635 -16441 16669
rect -16533 16619 -16441 16635
rect -16471 16517 -16441 16619
rect -16383 16740 -14383 16787
rect -16383 16706 -15875 16740
rect -14891 16723 -14383 16740
rect -14325 16740 -12325 16787
rect -14325 16723 -13817 16740
rect -14891 16706 -13817 16723
rect -12833 16723 -12325 16740
rect -12267 16740 -10267 16787
rect -12267 16723 -11759 16740
rect -12833 16706 -11759 16723
rect -10775 16723 -10267 16740
rect -10209 16740 -8209 16787
rect -10209 16723 -9701 16740
rect -10775 16706 -9701 16723
rect -8717 16706 -8209 16740
rect -16383 16598 -8209 16706
rect -16383 16564 -15875 16598
rect -14891 16581 -13817 16598
rect -14891 16564 -14383 16581
rect -16383 16517 -14383 16564
rect -14325 16564 -13817 16581
rect -12833 16581 -11759 16598
rect -12833 16564 -12325 16581
rect -14325 16517 -12325 16564
rect -12267 16564 -11759 16581
rect -10775 16581 -9701 16598
rect -10775 16564 -10267 16581
rect -12267 16517 -10267 16564
rect -10209 16564 -9701 16581
rect -8717 16564 -8209 16598
rect -10209 16517 -8209 16564
rect -8151 16685 -8121 16787
rect -8151 16669 -8059 16685
rect -8151 16635 -8109 16669
rect -8075 16635 -8059 16669
rect -8151 16619 -8059 16635
rect -8151 16517 -8121 16619
rect -16471 16291 -16441 16317
rect -16383 16270 -14383 16317
rect -16383 16253 -15875 16270
rect -15891 16236 -15875 16253
rect -14891 16253 -14383 16270
rect -14325 16270 -12325 16317
rect -14325 16253 -13817 16270
rect -14891 16236 -14875 16253
rect -15891 16220 -14875 16236
rect -13833 16236 -13817 16253
rect -12833 16253 -12325 16270
rect -12267 16270 -10267 16317
rect -12267 16253 -11759 16270
rect -12833 16236 -12817 16253
rect -13833 16220 -12817 16236
rect -11775 16236 -11759 16253
rect -10775 16253 -10267 16270
rect -10209 16270 -8209 16317
rect -8151 16291 -8121 16317
rect -10209 16253 -9701 16270
rect -10775 16236 -10759 16253
rect -11775 16220 -10759 16236
rect -9717 16236 -9701 16253
rect -8717 16253 -8209 16270
rect -8717 16236 -8701 16253
rect -9717 16220 -8701 16236
rect -15891 16119 -14875 16135
rect -15891 16102 -15875 16119
rect -16383 16085 -15875 16102
rect -14891 16102 -14875 16119
rect -13833 16119 -12817 16135
rect -13833 16102 -13817 16119
rect -14891 16085 -14383 16102
rect -16471 16038 -16441 16064
rect -16383 16038 -14383 16085
rect -14325 16085 -13817 16102
rect -12833 16102 -12817 16119
rect -11775 16119 -10759 16135
rect -11775 16102 -11759 16119
rect -12833 16085 -12325 16102
rect -14325 16038 -12325 16085
rect -12267 16085 -11759 16102
rect -10775 16102 -10759 16119
rect -9717 16119 -8701 16135
rect -9717 16102 -9701 16119
rect -10775 16085 -10267 16102
rect -12267 16038 -10267 16085
rect -10209 16085 -9701 16102
rect -8717 16102 -8701 16119
rect -8717 16085 -8209 16102
rect -10209 16038 -8209 16085
rect -8151 16038 -8121 16064
rect -16471 15807 -16441 15838
rect -16383 15812 -14383 15838
rect -14325 15812 -12325 15838
rect -12267 15812 -10267 15838
rect -10209 15812 -8209 15838
rect -16533 15791 -16441 15807
rect -16533 15757 -16517 15791
rect -16483 15757 -16441 15791
rect -16533 15741 -16441 15757
rect -8151 15807 -8121 15838
rect -8151 15791 -8059 15807
rect -8151 15757 -8109 15791
rect -8075 15757 -8059 15791
rect -8151 15741 -8059 15757
rect -7512 17453 -7420 17469
rect -7512 17419 -7496 17453
rect -7462 17419 -7420 17453
rect -7512 17403 -7420 17419
rect -7450 17372 -7420 17403
rect -3246 17453 -3154 17469
rect -3246 17419 -3204 17453
rect -3170 17419 -3154 17453
rect -3246 17403 -3154 17419
rect -7362 17372 -5362 17398
rect -5304 17372 -3304 17398
rect -3246 17372 -3216 17403
rect -7450 17146 -7420 17172
rect -7362 17125 -5362 17172
rect -7362 17108 -6854 17125
rect -6870 17091 -6854 17108
rect -5870 17108 -5362 17125
rect -5304 17125 -3304 17172
rect -3246 17146 -3216 17172
rect -5304 17108 -4796 17125
rect -5870 17091 -5854 17108
rect -6870 17075 -5854 17091
rect -4812 17091 -4796 17108
rect -3812 17108 -3304 17125
rect -3812 17091 -3796 17108
rect -4812 17075 -3796 17091
rect -7512 17021 -7420 17037
rect -7512 16987 -7496 17021
rect -7462 16987 -7420 17021
rect -7512 16971 -7420 16987
rect -7450 16940 -7420 16971
rect -3246 17021 -3154 17037
rect -3246 16987 -3204 17021
rect -3170 16987 -3154 17021
rect -3246 16971 -3154 16987
rect -7362 16940 -5362 16966
rect -5304 16940 -3304 16966
rect -3246 16940 -3216 16971
rect -7450 16714 -7420 16740
rect -7362 16693 -5362 16740
rect -7362 16676 -6854 16693
rect -6870 16659 -6854 16676
rect -5870 16676 -5362 16693
rect -5304 16693 -3304 16740
rect -3246 16714 -3216 16740
rect -5304 16676 -4796 16693
rect -5870 16659 -5854 16676
rect -6870 16643 -5854 16659
rect -4812 16659 -4796 16676
rect -3812 16676 -3304 16693
rect -3812 16659 -3796 16676
rect -4812 16643 -3796 16659
rect -6870 16551 -5854 16567
rect -6870 16534 -6854 16551
rect -7362 16517 -6854 16534
rect -5870 16534 -5854 16551
rect -4812 16551 -3796 16567
rect -4812 16534 -4796 16551
rect -5870 16517 -5362 16534
rect -7450 16470 -7420 16496
rect -7362 16470 -5362 16517
rect -5304 16517 -4796 16534
rect -3812 16534 -3796 16551
rect -3812 16517 -3304 16534
rect -5304 16470 -3304 16517
rect -3246 16470 -3216 16496
rect -7450 16239 -7420 16270
rect -7362 16244 -5362 16270
rect -5304 16244 -3304 16270
rect -7512 16223 -7420 16239
rect -7512 16189 -7496 16223
rect -7462 16189 -7420 16223
rect -7512 16173 -7420 16189
rect -3246 16239 -3216 16270
rect -3246 16223 -3154 16239
rect -3246 16189 -3204 16223
rect -3170 16189 -3154 16223
rect -3246 16174 -3154 16189
rect -3220 16173 -3154 16174
rect -6870 16119 -5854 16135
rect -6870 16102 -6854 16119
rect -7362 16085 -6854 16102
rect -5870 16102 -5854 16119
rect -4812 16119 -3796 16135
rect -4812 16102 -4796 16119
rect -5870 16085 -5362 16102
rect -7450 16038 -7420 16064
rect -7362 16038 -5362 16085
rect -5304 16085 -4796 16102
rect -3812 16102 -3796 16119
rect -3812 16085 -3304 16102
rect -5304 16038 -3304 16085
rect -3246 16038 -3216 16064
rect -7450 15807 -7420 15838
rect -7362 15812 -5362 15838
rect -5304 15812 -3304 15838
rect -7512 15791 -7420 15807
rect -7512 15757 -7496 15791
rect -7462 15757 -7420 15791
rect -7512 15741 -7420 15757
rect -3246 15807 -3216 15838
rect -3246 15791 -3154 15807
rect -3246 15757 -3204 15791
rect -3170 15757 -3154 15791
rect -3246 15741 -3154 15757
rect -1186 17524 -1094 17540
rect -1186 17490 -1170 17524
rect -1136 17490 -1094 17524
rect -1186 17474 -1094 17490
rect -1124 17452 -1094 17474
rect -1036 17524 -836 17540
rect -1036 17490 -1020 17524
rect -852 17490 -836 17524
rect -1036 17452 -836 17490
rect -778 17524 -578 17540
rect -778 17490 -762 17524
rect -594 17490 -578 17524
rect -778 17452 -578 17490
rect -520 17524 -428 17540
rect -520 17490 -478 17524
rect -444 17490 -428 17524
rect -520 17474 -428 17490
rect -520 17452 -490 17474
rect -1124 17226 -1094 17252
rect -1036 17237 -836 17252
rect -778 17237 -578 17252
rect -1036 17214 -578 17237
rect -520 17226 -490 17252
rect -1036 17180 -1020 17214
rect -852 17180 -762 17214
rect -594 17180 -578 17214
rect -1124 17142 -1094 17168
rect -1036 17157 -578 17180
rect -1036 17142 -836 17157
rect -778 17142 -578 17157
rect -520 17142 -490 17168
rect -1124 16920 -1094 16942
rect -1186 16904 -1094 16920
rect -1186 16870 -1170 16904
rect -1136 16870 -1094 16904
rect -1186 16854 -1094 16870
rect -1036 16904 -836 16942
rect -1036 16870 -1020 16904
rect -852 16870 -836 16904
rect -1036 16854 -836 16870
rect -778 16904 -578 16942
rect -778 16870 -762 16904
rect -594 16870 -578 16904
rect -778 16854 -578 16870
rect -520 16920 -490 16942
rect -520 16904 -428 16920
rect -520 16870 -478 16904
rect -444 16870 -428 16904
rect -520 16854 -428 16870
rect -108 17536 -16 17552
rect -108 17502 -92 17536
rect -58 17502 -16 17536
rect 5316 17536 7332 17552
rect 5316 17519 5332 17536
rect -108 17486 -16 17502
rect 4324 17502 5332 17519
rect 7316 17519 7332 17536
rect 8494 17536 8586 17552
rect 7316 17502 8324 17519
rect -46 17464 -16 17486
rect 154 17464 4154 17490
rect 4324 17464 8324 17502
rect 8494 17502 8536 17536
rect 8570 17502 8586 17536
rect 8494 17486 8586 17502
rect 8494 17464 8524 17486
rect -46 17238 -16 17264
rect 154 17239 4154 17264
rect 4324 17239 8324 17264
rect -108 17142 -16 17158
rect -108 17108 -92 17142
rect -58 17108 -16 17142
rect -108 17092 -16 17108
rect -46 17070 -16 17092
rect 154 17096 8324 17239
rect 8494 17238 8524 17264
rect 154 17070 4154 17096
rect 4324 17070 8324 17096
rect 8494 17142 8586 17158
rect 8494 17108 8536 17142
rect 8570 17108 8586 17142
rect 8494 17092 8586 17108
rect 8494 17070 8524 17092
rect -46 16844 -16 16870
rect 154 16845 4154 16870
rect 4324 16845 8324 16870
rect 154 16702 8324 16845
rect 8494 16844 8524 16870
rect -46 16676 -16 16702
rect 154 16676 4154 16702
rect 4324 16676 8324 16702
rect 8494 16676 8524 16702
rect -46 16454 -16 16476
rect -108 16438 -16 16454
rect -108 16404 -92 16438
rect -58 16404 -16 16438
rect -108 16388 -16 16404
rect 154 16451 4154 16476
rect 4324 16451 8324 16476
rect 154 16308 8324 16451
rect 8494 16454 8524 16476
rect 8494 16438 8586 16454
rect 8494 16404 8536 16438
rect 8570 16404 8586 16438
rect 8494 16388 8586 16404
rect -46 16282 -16 16308
rect 154 16282 4154 16308
rect 4324 16282 8324 16308
rect 8494 16282 8524 16308
rect -46 16060 -16 16082
rect -108 16044 -16 16060
rect -108 16010 -92 16044
rect -58 16010 -16 16044
rect 154 16044 4154 16082
rect 4324 16056 8324 16082
rect 8494 16060 8524 16082
rect 154 16027 1162 16044
rect -108 15994 -16 16010
rect 1146 16010 1162 16027
rect 3146 16027 4154 16044
rect 8494 16044 8586 16060
rect 3146 16010 3162 16027
rect 1146 15994 3162 16010
rect 8494 16010 8536 16044
rect 8570 16010 8586 16044
rect 8494 15994 8586 16010
rect -11742 15505 -10726 15521
rect -11742 15488 -11726 15505
rect -12234 15471 -11726 15488
rect -10742 15488 -10726 15505
rect -9684 15505 -8668 15521
rect -9684 15488 -9668 15505
rect -10742 15471 -10234 15488
rect -12322 15424 -12292 15450
rect -12234 15424 -10234 15471
rect -10176 15471 -9668 15488
rect -8684 15488 -8668 15505
rect -8684 15471 -8176 15488
rect -10176 15424 -8176 15471
rect -8118 15424 -8088 15450
rect -12322 15160 -12292 15224
rect -12384 15144 -12292 15160
rect -12384 15110 -12368 15144
rect -12334 15110 -12292 15144
rect -12384 15094 -12292 15110
rect -12322 15030 -12292 15094
rect -12234 15198 -10234 15224
rect -10176 15198 -8176 15224
rect -12234 15056 -8176 15198
rect -12234 15030 -10234 15056
rect -10176 15030 -8176 15056
rect -8118 15160 -8088 15224
rect -8118 15144 -8026 15160
rect -8118 15110 -8076 15144
rect -8042 15110 -8026 15144
rect -8118 15094 -8026 15110
rect -8118 15030 -8088 15094
rect -12322 14804 -12292 14830
rect -12234 14783 -10234 14830
rect -12234 14766 -11726 14783
rect -11742 14749 -11726 14766
rect -10742 14766 -10234 14783
rect -10176 14783 -8176 14830
rect -8118 14804 -8088 14830
rect -10176 14766 -9668 14783
rect -10742 14749 -10726 14766
rect -11742 14733 -10726 14749
rect -9684 14749 -9668 14766
rect -8684 14766 -8176 14783
rect -8684 14749 -8668 14766
rect -9684 14733 -8668 14749
rect -7416 15489 -7386 15515
rect -7328 15489 -5328 15515
rect -5270 15489 -3270 15515
rect -3212 15489 -3182 15515
rect -7416 15257 -7386 15289
rect -7478 15241 -7386 15257
rect -7478 15207 -7462 15241
rect -7428 15207 -7386 15241
rect -7328 15242 -5328 15289
rect -7328 15225 -6820 15242
rect -7478 15191 -7386 15207
rect -6836 15208 -6820 15225
rect -5836 15225 -5328 15242
rect -5270 15242 -3270 15289
rect -5270 15225 -4762 15242
rect -5836 15208 -5820 15225
rect -6836 15192 -5820 15208
rect -4778 15208 -4762 15225
rect -3778 15225 -3270 15242
rect -3212 15258 -3182 15289
rect -3212 15242 -3120 15258
rect -3778 15208 -3762 15225
rect -4778 15192 -3762 15208
rect -3212 15208 -3170 15242
rect -3136 15208 -3120 15242
rect -3212 15192 -3120 15208
rect -7478 15094 -7386 15110
rect -7478 15060 -7462 15094
rect -7428 15060 -7386 15094
rect -6836 15094 -5820 15110
rect -6836 15077 -6820 15094
rect -7478 15044 -7386 15060
rect -7416 15013 -7386 15044
rect -7328 15060 -6820 15077
rect -5836 15077 -5820 15094
rect -4778 15094 -3762 15110
rect -4778 15077 -4762 15094
rect -5836 15060 -5328 15077
rect -7328 15013 -5328 15060
rect -5270 15060 -4762 15077
rect -3778 15077 -3762 15094
rect -3212 15094 -3120 15110
rect -3778 15060 -3270 15077
rect -5270 15013 -3270 15060
rect -3212 15060 -3170 15094
rect -3136 15060 -3120 15094
rect -3212 15044 -3120 15060
rect -3212 15013 -3182 15044
rect -7416 14787 -7386 14813
rect -7328 14787 -5328 14813
rect -5270 14787 -3270 14813
rect -3212 14787 -3182 14813
rect 3789 15618 5105 15634
rect 3789 15601 3805 15618
rect 3147 15584 3805 15601
rect 5089 15601 5105 15618
rect 6447 15618 7763 15634
rect 6447 15601 6463 15618
rect 5089 15584 5747 15601
rect 3059 15546 3089 15572
rect 3147 15546 5747 15584
rect 5805 15584 6463 15601
rect 7747 15601 7763 15618
rect 7747 15584 8405 15601
rect 5805 15546 8405 15584
rect 8463 15546 8493 15572
rect 3059 15344 3089 15366
rect 2997 15328 3089 15344
rect 2997 15294 3013 15328
rect 3047 15294 3089 15328
rect 3147 15328 5747 15366
rect 3147 15311 3805 15328
rect 2997 15278 3089 15294
rect 3789 15294 3805 15311
rect 5089 15311 5747 15328
rect 5805 15328 8405 15366
rect 5805 15311 6463 15328
rect 5089 15294 5105 15311
rect 3789 15278 5105 15294
rect 6447 15294 6463 15311
rect 7747 15311 8405 15328
rect 8463 15344 8493 15366
rect 8463 15328 8555 15344
rect 7747 15294 7763 15311
rect 6447 15278 7763 15294
rect 8463 15294 8505 15328
rect 8539 15294 8555 15328
rect 8463 15278 8555 15294
rect 2997 15186 3089 15202
rect 2997 15152 3013 15186
rect 3047 15152 3089 15186
rect 3789 15186 5105 15202
rect 3789 15169 3805 15186
rect 2997 15136 3089 15152
rect 3059 15114 3089 15136
rect 3147 15152 3805 15169
rect 5089 15169 5105 15186
rect 6447 15186 7763 15202
rect 6447 15169 6463 15186
rect 5089 15152 5747 15169
rect 3147 15114 5747 15152
rect 5805 15152 6463 15169
rect 7747 15169 7763 15186
rect 8463 15186 8555 15202
rect 7747 15152 8405 15169
rect 5805 15114 8405 15152
rect 8463 15152 8505 15186
rect 8539 15152 8555 15186
rect 8463 15136 8555 15152
rect 8463 15114 8493 15136
rect 3059 14908 3089 14934
rect 3147 14908 5747 14934
rect 5805 14908 8405 14934
rect 8463 14908 8493 14934
rect 838 12250 1038 12266
rect 838 12216 854 12250
rect 1022 12216 1038 12250
rect 750 12178 780 12204
rect 838 12178 1038 12216
rect 1096 12250 1296 12266
rect 1096 12216 1112 12250
rect 1280 12216 1296 12250
rect 1096 12178 1296 12216
rect 1354 12178 1384 12204
rect 750 11314 780 11378
rect 688 11298 780 11314
rect 688 11264 704 11298
rect 738 11264 780 11298
rect 688 11248 780 11264
rect 750 11184 780 11248
rect 838 11352 1038 11378
rect 1096 11352 1296 11378
rect 838 11210 1296 11352
rect 838 11184 1038 11210
rect 1096 11184 1296 11210
rect 1354 11314 1384 11378
rect 1354 11298 1446 11314
rect 1354 11264 1396 11298
rect 1430 11264 1446 11298
rect 1354 11248 1446 11264
rect 1354 11184 1384 11248
rect 750 10358 780 10384
rect 838 10346 1038 10384
rect 838 10312 854 10346
rect 1022 10312 1038 10346
rect 838 10296 1038 10312
rect 1096 10346 1296 10384
rect 1354 10358 1384 10384
rect 1096 10312 1112 10346
rect 1280 10312 1296 10346
rect 1096 10296 1296 10312
rect 1730 12250 1930 12266
rect 1730 12216 1746 12250
rect 1914 12216 1930 12250
rect 1642 12178 1672 12204
rect 1730 12178 1930 12216
rect 1988 12250 2188 12266
rect 1988 12216 2004 12250
rect 2172 12216 2188 12250
rect 1988 12178 2188 12216
rect 2246 12178 2276 12204
rect 1642 11314 1672 11378
rect 1580 11298 1672 11314
rect 1580 11264 1596 11298
rect 1630 11264 1672 11298
rect 1580 11248 1672 11264
rect 1642 11184 1672 11248
rect 1730 11352 1930 11378
rect 1988 11352 2188 11378
rect 1730 11210 2188 11352
rect 1730 11184 1930 11210
rect 1988 11184 2188 11210
rect 2246 11314 2276 11378
rect 2246 11298 2338 11314
rect 2246 11264 2288 11298
rect 2322 11264 2338 11298
rect 2246 11248 2338 11264
rect 2246 11184 2276 11248
rect 1642 10358 1672 10384
rect 1730 10346 1930 10384
rect 1730 10312 1746 10346
rect 1914 10312 1930 10346
rect 1730 10296 1930 10312
rect 1988 10346 2188 10384
rect 2246 10358 2276 10384
rect 1988 10312 2004 10346
rect 2172 10312 2188 10346
rect 1988 10296 2188 10312
rect 2622 12250 2822 12266
rect 2622 12216 2638 12250
rect 2806 12216 2822 12250
rect 2534 12178 2564 12204
rect 2622 12178 2822 12216
rect 2880 12250 3080 12266
rect 2880 12216 2896 12250
rect 3064 12216 3080 12250
rect 2880 12178 3080 12216
rect 3138 12178 3168 12204
rect 2534 11314 2564 11378
rect 2472 11298 2564 11314
rect 2472 11264 2488 11298
rect 2522 11264 2564 11298
rect 2472 11248 2564 11264
rect 2534 11184 2564 11248
rect 2622 11352 2822 11378
rect 2880 11352 3080 11378
rect 2622 11210 3080 11352
rect 2622 11184 2822 11210
rect 2880 11184 3080 11210
rect 3138 11314 3168 11378
rect 3138 11298 3230 11314
rect 3138 11264 3180 11298
rect 3214 11264 3230 11298
rect 3138 11248 3230 11264
rect 3138 11184 3168 11248
rect 2534 10358 2564 10384
rect 2622 10346 2822 10384
rect 2622 10312 2638 10346
rect 2806 10312 2822 10346
rect 2622 10296 2822 10312
rect 2880 10346 3080 10384
rect 3138 10358 3168 10384
rect 2880 10312 2896 10346
rect 3064 10312 3080 10346
rect 2880 10296 3080 10312
rect 3514 12250 3714 12266
rect 3514 12216 3530 12250
rect 3698 12216 3714 12250
rect 3426 12178 3456 12204
rect 3514 12178 3714 12216
rect 3772 12250 3972 12266
rect 3772 12216 3788 12250
rect 3956 12216 3972 12250
rect 3772 12178 3972 12216
rect 4030 12178 4060 12204
rect 3426 11314 3456 11378
rect 3364 11298 3456 11314
rect 3364 11264 3380 11298
rect 3414 11264 3456 11298
rect 3364 11248 3456 11264
rect 3426 11184 3456 11248
rect 3514 11352 3714 11378
rect 3772 11352 3972 11378
rect 3514 11210 3972 11352
rect 3514 11184 3714 11210
rect 3772 11184 3972 11210
rect 4030 11314 4060 11378
rect 4030 11298 4122 11314
rect 4030 11264 4072 11298
rect 4106 11264 4122 11298
rect 4030 11248 4122 11264
rect 4030 11184 4060 11248
rect 3426 10358 3456 10384
rect 3514 10346 3714 10384
rect 3514 10312 3530 10346
rect 3698 10312 3714 10346
rect 3514 10296 3714 10312
rect 3772 10346 3972 10384
rect 4030 10358 4060 10384
rect 3772 10312 3788 10346
rect 3956 10312 3972 10346
rect 3772 10296 3972 10312
rect 4328 12201 4394 12217
rect 4328 12167 4344 12201
rect 4378 12167 4394 12201
rect 4328 12155 4394 12167
rect 4328 12125 4416 12155
rect 4616 12125 4642 12155
rect 4390 11867 4416 12067
rect 4616 12051 4704 12067
rect 4616 11883 4654 12051
rect 4688 11883 4704 12051
rect 4616 11867 4704 11883
rect 4390 11609 4416 11809
rect 4616 11793 4704 11809
rect 4616 11625 4654 11793
rect 4688 11625 4704 11793
rect 4616 11609 4704 11625
rect 4328 11521 4416 11551
rect 4616 11521 4642 11551
rect 4328 11509 4394 11521
rect 4328 11475 4344 11509
rect 4378 11475 4394 11509
rect 4328 11459 4394 11475
rect 4328 11087 4394 11103
rect 4328 11053 4344 11087
rect 4378 11053 4394 11087
rect 4328 11041 4394 11053
rect 4328 11011 4416 11041
rect 4616 11011 4642 11041
rect 4390 10753 4416 10953
rect 4616 10937 4704 10953
rect 4616 10769 4654 10937
rect 4688 10769 4704 10937
rect 4616 10753 4704 10769
rect 4390 10495 4416 10695
rect 4616 10679 4704 10695
rect 4616 10511 4654 10679
rect 4688 10511 4704 10679
rect 4616 10495 4704 10511
rect 4328 10407 4416 10437
rect 4616 10407 4642 10437
rect 4328 10395 4394 10407
rect 4328 10361 4344 10395
rect 4378 10361 4394 10395
rect 4328 10345 4394 10361
rect 5453 11812 5519 11822
rect 5453 11778 5469 11812
rect 5503 11778 5519 11812
rect 5453 11766 5519 11778
rect 4963 11736 4989 11766
rect 5389 11736 5583 11766
rect 5983 11736 6009 11766
rect 4925 11586 4989 11678
rect 4892 11570 4989 11586
rect 4892 11386 4908 11570
rect 4942 11386 4989 11570
rect 4892 11370 4989 11386
rect 4925 11278 4989 11370
rect 5389 11278 5583 11678
rect 5983 11586 6047 11678
rect 5983 11570 6080 11586
rect 5983 11386 6030 11570
rect 6064 11386 6080 11570
rect 5983 11370 6080 11386
rect 5983 11278 6047 11370
rect 5415 11220 5557 11278
rect 4925 11128 4989 11220
rect 4892 11112 4989 11128
rect 4892 10928 4908 11112
rect 4942 10928 4989 11112
rect 4892 10912 4989 10928
rect 4925 10820 4989 10912
rect 5389 10820 5583 11220
rect 5983 11128 6047 11220
rect 5983 11112 6080 11128
rect 5983 10928 6030 11112
rect 6064 10928 6080 11112
rect 5983 10912 6080 10928
rect 5983 10820 6047 10912
rect 4963 10732 4989 10762
rect 5389 10732 5583 10762
rect 5983 10732 6009 10762
rect 5453 10720 5519 10732
rect 5453 10686 5469 10720
rect 5503 10686 5519 10720
rect 5453 10676 5519 10686
<< polycont >>
rect -16517 17513 -16483 17547
rect -8109 17513 -8075 17547
rect -15875 17185 -14891 17219
rect -13817 17185 -12833 17219
rect -11759 17185 -10775 17219
rect -9701 17185 -8717 17219
rect -15875 17034 -14891 17068
rect -13817 17034 -12833 17068
rect -11759 17034 -10775 17068
rect -9701 17034 -8717 17068
rect -16517 16635 -16483 16669
rect -15875 16706 -14891 16740
rect -13817 16706 -12833 16740
rect -11759 16706 -10775 16740
rect -9701 16706 -8717 16740
rect -15875 16564 -14891 16598
rect -13817 16564 -12833 16598
rect -11759 16564 -10775 16598
rect -9701 16564 -8717 16598
rect -8109 16635 -8075 16669
rect -15875 16236 -14891 16270
rect -13817 16236 -12833 16270
rect -11759 16236 -10775 16270
rect -9701 16236 -8717 16270
rect -15875 16085 -14891 16119
rect -13817 16085 -12833 16119
rect -11759 16085 -10775 16119
rect -9701 16085 -8717 16119
rect -16517 15757 -16483 15791
rect -8109 15757 -8075 15791
rect -7496 17419 -7462 17453
rect -3204 17419 -3170 17453
rect -6854 17091 -5870 17125
rect -4796 17091 -3812 17125
rect -7496 16987 -7462 17021
rect -3204 16987 -3170 17021
rect -6854 16659 -5870 16693
rect -4796 16659 -3812 16693
rect -6854 16517 -5870 16551
rect -4796 16517 -3812 16551
rect -7496 16189 -7462 16223
rect -3204 16189 -3170 16223
rect -6854 16085 -5870 16119
rect -4796 16085 -3812 16119
rect -7496 15757 -7462 15791
rect -3204 15757 -3170 15791
rect -1170 17490 -1136 17524
rect -1020 17490 -852 17524
rect -762 17490 -594 17524
rect -478 17490 -444 17524
rect -1020 17180 -852 17214
rect -762 17180 -594 17214
rect -1170 16870 -1136 16904
rect -1020 16870 -852 16904
rect -762 16870 -594 16904
rect -478 16870 -444 16904
rect -92 17502 -58 17536
rect 5332 17502 7316 17536
rect 8536 17502 8570 17536
rect -92 17108 -58 17142
rect 8536 17108 8570 17142
rect -92 16404 -58 16438
rect 8536 16404 8570 16438
rect -92 16010 -58 16044
rect 1162 16010 3146 16044
rect 8536 16010 8570 16044
rect -11726 15471 -10742 15505
rect -9668 15471 -8684 15505
rect -12368 15110 -12334 15144
rect -8076 15110 -8042 15144
rect -11726 14749 -10742 14783
rect -9668 14749 -8684 14783
rect -7462 15207 -7428 15241
rect -6820 15208 -5836 15242
rect -4762 15208 -3778 15242
rect -3170 15208 -3136 15242
rect -7462 15060 -7428 15094
rect -6820 15060 -5836 15094
rect -4762 15060 -3778 15094
rect -3170 15060 -3136 15094
rect 3805 15584 5089 15618
rect 6463 15584 7747 15618
rect 3013 15294 3047 15328
rect 3805 15294 5089 15328
rect 6463 15294 7747 15328
rect 8505 15294 8539 15328
rect 3013 15152 3047 15186
rect 3805 15152 5089 15186
rect 6463 15152 7747 15186
rect 8505 15152 8539 15186
rect 854 12216 1022 12250
rect 1112 12216 1280 12250
rect 704 11264 738 11298
rect 1396 11264 1430 11298
rect 854 10312 1022 10346
rect 1112 10312 1280 10346
rect 1746 12216 1914 12250
rect 2004 12216 2172 12250
rect 1596 11264 1630 11298
rect 2288 11264 2322 11298
rect 1746 10312 1914 10346
rect 2004 10312 2172 10346
rect 2638 12216 2806 12250
rect 2896 12216 3064 12250
rect 2488 11264 2522 11298
rect 3180 11264 3214 11298
rect 2638 10312 2806 10346
rect 2896 10312 3064 10346
rect 3530 12216 3698 12250
rect 3788 12216 3956 12250
rect 3380 11264 3414 11298
rect 4072 11264 4106 11298
rect 3530 10312 3698 10346
rect 3788 10312 3956 10346
rect 4344 12167 4378 12201
rect 4654 11883 4688 12051
rect 4654 11625 4688 11793
rect 4344 11475 4378 11509
rect 4344 11053 4378 11087
rect 4654 10769 4688 10937
rect 4654 10511 4688 10679
rect 4344 10361 4378 10395
rect 5469 11778 5503 11812
rect 4908 11386 4942 11570
rect 6030 11386 6064 11570
rect 4908 10928 4942 11112
rect 6030 10928 6064 11112
rect 5469 10686 5503 10720
<< xpolycontact >>
rect -17355 22491 -16923 22561
rect -13555 22491 -13123 22561
rect -13019 22491 -12587 22561
rect -9219 22491 -8787 22561
rect -8683 22491 -8251 22561
rect -4883 22491 -4451 22561
rect -4347 22491 -3915 22561
rect -547 22491 -115 22561
rect -11 22491 421 22561
rect 3789 22491 4221 22561
rect 4325 22491 4757 22561
rect 8125 22491 8557 22561
rect -17355 22325 -16923 22395
rect -13555 22325 -13123 22395
rect -13019 22325 -12587 22395
rect -9219 22325 -8787 22395
rect -8683 22325 -8251 22395
rect -4883 22325 -4451 22395
rect -4347 22325 -3915 22395
rect -547 22325 -115 22395
rect -11 22325 421 22395
rect 3789 22325 4221 22395
rect 4325 22325 4757 22395
rect 8125 22325 8557 22395
rect -17355 22159 -16923 22229
rect -13555 22159 -13123 22229
rect -13019 22159 -12587 22229
rect -9219 22159 -8787 22229
rect -8683 22159 -8251 22229
rect -4883 22159 -4451 22229
rect -4347 22159 -3915 22229
rect -547 22159 -115 22229
rect -11 22159 421 22229
rect 3789 22159 4221 22229
rect 4325 22159 4757 22229
rect 8125 22159 8557 22229
rect -17355 21993 -16923 22063
rect -13555 21993 -13123 22063
rect -13019 21993 -12587 22063
rect -9219 21993 -8787 22063
rect -8683 21993 -8251 22063
rect -4883 21993 -4451 22063
rect -4347 21993 -3915 22063
rect -547 21993 -115 22063
rect -11 21993 421 22063
rect 3789 21993 4221 22063
rect 4325 21993 4757 22063
rect 8125 21993 8557 22063
rect -17355 21827 -16923 21897
rect -13555 21827 -13123 21897
rect -13019 21827 -12587 21897
rect -9219 21827 -8787 21897
rect -8683 21827 -8251 21897
rect -4883 21827 -4451 21897
rect -4347 21827 -3915 21897
rect -547 21827 -115 21897
rect -11 21827 421 21897
rect 3789 21827 4221 21897
rect 4325 21827 4757 21897
rect 8125 21827 8557 21897
rect -17355 21661 -16923 21731
rect -13555 21661 -13123 21731
rect -13019 21661 -12587 21731
rect -9219 21661 -8787 21731
rect -8683 21661 -8251 21731
rect -4883 21661 -4451 21731
rect -4347 21661 -3915 21731
rect -547 21661 -115 21731
rect -11 21661 421 21731
rect 3789 21661 4221 21731
rect 4325 21661 4757 21731
rect 8125 21661 8557 21731
rect -17355 21495 -16923 21565
rect -13555 21495 -13123 21565
rect -13019 21495 -12587 21565
rect -9219 21495 -8787 21565
rect -8683 21495 -8251 21565
rect -4883 21495 -4451 21565
rect -4347 21495 -3915 21565
rect -547 21495 -115 21565
rect -11 21495 421 21565
rect 3789 21495 4221 21565
rect 4325 21495 4757 21565
rect 8125 21495 8557 21565
rect -17355 21329 -16923 21399
rect -13555 21329 -13123 21399
rect -13019 21329 -12587 21399
rect -9219 21329 -8787 21399
rect -8683 21329 -8251 21399
rect -4883 21329 -4451 21399
rect -4347 21329 -3915 21399
rect -547 21329 -115 21399
rect -11 21329 421 21399
rect 3789 21329 4221 21399
rect 4325 21329 4757 21399
rect 8125 21329 8557 21399
rect -17355 21163 -16923 21233
rect -13555 21163 -13123 21233
rect -13019 21163 -12587 21233
rect -9219 21163 -8787 21233
rect -8683 21163 -8251 21233
rect -4883 21163 -4451 21233
rect -4347 21163 -3915 21233
rect -547 21163 -115 21233
rect -11 21163 421 21233
rect 3789 21163 4221 21233
rect 4325 21163 4757 21233
rect 8125 21163 8557 21233
rect -17355 20997 -16923 21067
rect -13555 20997 -13123 21067
rect -13019 20997 -12587 21067
rect -9219 20997 -8787 21067
rect -8683 20997 -8251 21067
rect -4883 20997 -4451 21067
rect -4347 20997 -3915 21067
rect -547 20997 -115 21067
rect -11 20997 421 21067
rect 3789 20997 4221 21067
rect 4325 20997 4757 21067
rect 8125 20997 8557 21067
rect -13019 20595 -12587 20665
rect -9219 20595 -8787 20665
rect -8683 20595 -8251 20665
rect -4883 20595 -4451 20665
rect -4347 20595 -3915 20665
rect -547 20595 -115 20665
rect -11 20595 421 20665
rect 3789 20595 4221 20665
rect 4325 20595 4757 20665
rect 8125 20595 8557 20665
rect -13019 20429 -12587 20499
rect -9219 20429 -8787 20499
rect -8683 20429 -8251 20499
rect -4883 20429 -4451 20499
rect -4347 20429 -3915 20499
rect -547 20429 -115 20499
rect -11 20429 421 20499
rect 3789 20429 4221 20499
rect 4325 20429 4757 20499
rect 8125 20429 8557 20499
rect -13019 20263 -12587 20333
rect -9219 20263 -8787 20333
rect -8683 20263 -8251 20333
rect -4883 20263 -4451 20333
rect -4347 20263 -3915 20333
rect -547 20263 -115 20333
rect -11 20263 421 20333
rect 3789 20263 4221 20333
rect 4325 20263 4757 20333
rect 8125 20263 8557 20333
rect -13019 20097 -12587 20167
rect -9219 20097 -8787 20167
rect -8683 20097 -8251 20167
rect -4883 20097 -4451 20167
rect -4347 20097 -3915 20167
rect -547 20097 -115 20167
rect -11 20097 421 20167
rect 3789 20097 4221 20167
rect 4325 20097 4757 20167
rect 8125 20097 8557 20167
rect -13019 19931 -12587 20001
rect -9219 19931 -8787 20001
rect -8683 19931 -8251 20001
rect -4883 19931 -4451 20001
rect -4347 19931 -3915 20001
rect -547 19931 -115 20001
rect -11 19931 421 20001
rect 3789 19931 4221 20001
rect 4325 19931 4757 20001
rect 8125 19931 8557 20001
rect -13019 19765 -12587 19835
rect -9219 19765 -8787 19835
rect -8683 19765 -8251 19835
rect -4883 19765 -4451 19835
rect -4347 19765 -3915 19835
rect -547 19765 -115 19835
rect -11 19765 421 19835
rect 3789 19765 4221 19835
rect 4325 19765 4757 19835
rect 8125 19765 8557 19835
rect -13019 19599 -12587 19669
rect -9219 19599 -8787 19669
rect -8683 19599 -8251 19669
rect -4883 19599 -4451 19669
rect -4347 19599 -3915 19669
rect -547 19599 -115 19669
rect -11 19599 421 19669
rect 3789 19599 4221 19669
rect 4325 19599 4757 19669
rect 8125 19599 8557 19669
rect -13019 19433 -12587 19503
rect -9219 19433 -8787 19503
rect -8683 19433 -8251 19503
rect -4883 19433 -4451 19503
rect -4347 19433 -3915 19503
rect -547 19433 -115 19503
rect -11 19433 421 19503
rect 3789 19433 4221 19503
rect 4325 19433 4757 19503
rect 8125 19433 8557 19503
rect -7035 19031 -6603 19101
rect -4955 19031 -4523 19101
rect -4419 19031 -3987 19101
rect -2339 19031 -1907 19101
rect -1803 19031 -1371 19101
rect 277 19031 709 19101
rect 813 19031 1245 19101
rect 2893 19031 3325 19101
rect 3429 19031 3861 19101
rect 5509 19031 5941 19101
rect 6045 19031 6477 19101
rect 8125 19031 8557 19101
rect -7035 18865 -6603 18935
rect -4955 18865 -4523 18935
rect -4419 18865 -3987 18935
rect -2339 18865 -1907 18935
rect -1803 18865 -1371 18935
rect 277 18865 709 18935
rect 813 18865 1245 18935
rect 2893 18865 3325 18935
rect 3429 18865 3861 18935
rect 5509 18865 5941 18935
rect 6045 18865 6477 18935
rect 8125 18865 8557 18935
rect -7035 18699 -6603 18769
rect -4955 18699 -4523 18769
rect -4419 18699 -3987 18769
rect -2339 18699 -1907 18769
rect -1803 18699 -1371 18769
rect 277 18699 709 18769
rect 813 18699 1245 18769
rect 2893 18699 3325 18769
rect 3429 18699 3861 18769
rect 5509 18699 5941 18769
rect 6045 18699 6477 18769
rect 8125 18699 8557 18769
rect -7035 18533 -6603 18603
rect -4955 18533 -4523 18603
rect -4419 18533 -3987 18603
rect -2339 18533 -1907 18603
rect -1803 18533 -1371 18603
rect 277 18533 709 18603
rect 813 18533 1245 18603
rect 2893 18533 3325 18603
rect 3429 18533 3861 18603
rect 5509 18533 5941 18603
rect 6045 18533 6477 18603
rect 8125 18533 8557 18603
rect -7035 18367 -6603 18437
rect -4955 18367 -4523 18437
rect -4419 18367 -3987 18437
rect -2339 18367 -1907 18437
rect -1803 18367 -1371 18437
rect 277 18367 709 18437
rect 813 18367 1245 18437
rect 2893 18367 3325 18437
rect 3429 18367 3861 18437
rect 5509 18367 5941 18437
rect 6045 18367 6477 18437
rect 8125 18367 8557 18437
rect -7035 18201 -6603 18271
rect -4955 18201 -4523 18271
rect -4419 18201 -3987 18271
rect -2339 18201 -1907 18271
rect -1803 18201 -1371 18271
rect 277 18201 709 18271
rect 813 18201 1245 18271
rect 2893 18201 3325 18271
rect 3429 18201 3861 18271
rect 5509 18201 5941 18271
rect 6045 18201 6477 18271
rect 8125 18201 8557 18271
rect -7035 18035 -6603 18105
rect -4955 18035 -4523 18105
rect -4419 18035 -3987 18105
rect -2339 18035 -1907 18105
rect -1803 18035 -1371 18105
rect 277 18035 709 18105
rect 813 18035 1245 18105
rect 2893 18035 3325 18105
rect 3429 18035 3861 18105
rect 5509 18035 5941 18105
rect 6045 18035 6477 18105
rect 8125 18035 8557 18105
rect -7035 17869 -6603 17939
rect -4955 17869 -4523 17939
rect -4419 17869 -3987 17939
rect -2339 17869 -1907 17939
rect -1803 17869 -1371 17939
rect 277 17869 709 17939
rect 813 17869 1245 17939
rect 2893 17869 3325 17939
rect 3429 17869 3861 17939
rect 5509 17869 5941 17939
rect 6045 17869 6477 17939
rect 8125 17869 8557 17939
rect -1080 15663 -648 15733
rect 220 15663 652 15733
rect 756 15663 1188 15733
rect 2056 15663 2488 15733
rect -1080 15497 -648 15567
rect 220 15497 652 15567
rect 756 15497 1188 15567
rect 2056 15497 2488 15567
rect -1080 15331 -648 15401
rect 220 15331 652 15401
rect 756 15331 1188 15401
rect 2056 15331 2488 15401
rect -1080 15165 -648 15235
rect 220 15165 652 15235
rect 756 15165 1188 15235
rect 2056 15165 2488 15235
rect -1080 14999 -648 15069
rect 220 14999 652 15069
rect 756 14999 1188 15069
rect 2056 14999 2488 15069
rect -1080 14833 -648 14903
rect 220 14833 652 14903
rect 756 14833 1188 14903
rect 2056 14833 2488 14903
<< ppolyres >>
rect -16923 22491 -13555 22561
rect -12587 22491 -9219 22561
rect -8251 22491 -4883 22561
rect -3915 22491 -547 22561
rect 421 22491 3789 22561
rect 4757 22491 8125 22561
rect -16923 22325 -13555 22395
rect -12587 22325 -9219 22395
rect -8251 22325 -4883 22395
rect -3915 22325 -547 22395
rect 421 22325 3789 22395
rect 4757 22325 8125 22395
rect -16923 22159 -13555 22229
rect -12587 22159 -9219 22229
rect -8251 22159 -4883 22229
rect -3915 22159 -547 22229
rect 421 22159 3789 22229
rect 4757 22159 8125 22229
rect -16923 21993 -13555 22063
rect -12587 21993 -9219 22063
rect -8251 21993 -4883 22063
rect -3915 21993 -547 22063
rect 421 21993 3789 22063
rect 4757 21993 8125 22063
rect -16923 21827 -13555 21897
rect -12587 21827 -9219 21897
rect -8251 21827 -4883 21897
rect -3915 21827 -547 21897
rect 421 21827 3789 21897
rect 4757 21827 8125 21897
rect -16923 21661 -13555 21731
rect -12587 21661 -9219 21731
rect -8251 21661 -4883 21731
rect -3915 21661 -547 21731
rect 421 21661 3789 21731
rect 4757 21661 8125 21731
rect -16923 21495 -13555 21565
rect -12587 21495 -9219 21565
rect -8251 21495 -4883 21565
rect -3915 21495 -547 21565
rect 421 21495 3789 21565
rect 4757 21495 8125 21565
rect -16923 21329 -13555 21399
rect -12587 21329 -9219 21399
rect -8251 21329 -4883 21399
rect -3915 21329 -547 21399
rect 421 21329 3789 21399
rect 4757 21329 8125 21399
rect -16923 21163 -13555 21233
rect -12587 21163 -9219 21233
rect -8251 21163 -4883 21233
rect -3915 21163 -547 21233
rect 421 21163 3789 21233
rect 4757 21163 8125 21233
rect -16923 20997 -13555 21067
rect -12587 20997 -9219 21067
rect -8251 20997 -4883 21067
rect -3915 20997 -547 21067
rect 421 20997 3789 21067
rect 4757 20997 8125 21067
rect -12587 20595 -9219 20665
rect -8251 20595 -4883 20665
rect -3915 20595 -547 20665
rect 421 20595 3789 20665
rect 4757 20595 8125 20665
rect -12587 20429 -9219 20499
rect -8251 20429 -4883 20499
rect -3915 20429 -547 20499
rect 421 20429 3789 20499
rect 4757 20429 8125 20499
rect -12587 20263 -9219 20333
rect -8251 20263 -4883 20333
rect -3915 20263 -547 20333
rect 421 20263 3789 20333
rect 4757 20263 8125 20333
rect -12587 20097 -9219 20167
rect -8251 20097 -4883 20167
rect -3915 20097 -547 20167
rect 421 20097 3789 20167
rect 4757 20097 8125 20167
rect -12587 19931 -9219 20001
rect -8251 19931 -4883 20001
rect -3915 19931 -547 20001
rect 421 19931 3789 20001
rect 4757 19931 8125 20001
rect -12587 19765 -9219 19835
rect -8251 19765 -4883 19835
rect -3915 19765 -547 19835
rect 421 19765 3789 19835
rect 4757 19765 8125 19835
rect -12587 19599 -9219 19669
rect -8251 19599 -4883 19669
rect -3915 19599 -547 19669
rect 421 19599 3789 19669
rect 4757 19599 8125 19669
rect -12587 19433 -9219 19503
rect -8251 19433 -4883 19503
rect -3915 19433 -547 19503
rect 421 19433 3789 19503
rect 4757 19433 8125 19503
rect -6603 19031 -4955 19101
rect -3987 19031 -2339 19101
rect -1371 19031 277 19101
rect 1245 19031 2893 19101
rect 3861 19031 5509 19101
rect 6477 19031 8125 19101
rect -6603 18865 -4955 18935
rect -3987 18865 -2339 18935
rect -1371 18865 277 18935
rect 1245 18865 2893 18935
rect 3861 18865 5509 18935
rect 6477 18865 8125 18935
rect -6603 18699 -4955 18769
rect -3987 18699 -2339 18769
rect -1371 18699 277 18769
rect 1245 18699 2893 18769
rect 3861 18699 5509 18769
rect 6477 18699 8125 18769
rect -6603 18533 -4955 18603
rect -3987 18533 -2339 18603
rect -1371 18533 277 18603
rect 1245 18533 2893 18603
rect 3861 18533 5509 18603
rect 6477 18533 8125 18603
rect -6603 18367 -4955 18437
rect -3987 18367 -2339 18437
rect -1371 18367 277 18437
rect 1245 18367 2893 18437
rect 3861 18367 5509 18437
rect 6477 18367 8125 18437
rect -6603 18201 -4955 18271
rect -3987 18201 -2339 18271
rect -1371 18201 277 18271
rect 1245 18201 2893 18271
rect 3861 18201 5509 18271
rect 6477 18201 8125 18271
rect -6603 18035 -4955 18105
rect -3987 18035 -2339 18105
rect -1371 18035 277 18105
rect 1245 18035 2893 18105
rect 3861 18035 5509 18105
rect 6477 18035 8125 18105
rect -6603 17869 -4955 17939
rect -3987 17869 -2339 17939
rect -1371 17869 277 17939
rect 1245 17869 2893 17939
rect 3861 17869 5509 17939
rect 6477 17869 8125 17939
rect -648 15663 220 15733
rect 1188 15663 2056 15733
rect -648 15497 220 15567
rect 1188 15497 2056 15567
rect -648 15331 220 15401
rect 1188 15331 2056 15401
rect -648 15165 220 15235
rect 1188 15165 2056 15235
rect -648 14999 220 15069
rect 1188 14999 2056 15069
rect -648 14833 220 14903
rect 1188 14833 2056 14903
<< locali >>
rect -17937 22967 -17877 23001
rect 9141 22967 9201 23001
rect -17937 22941 -17903 22967
rect 9167 22941 9201 22967
rect -7165 19197 -7069 19231
rect 8591 19197 8687 19231
rect -7165 19135 -7131 19197
rect 8653 19135 8687 19197
rect -7165 17773 -7131 17835
rect 8653 17773 8687 17835
rect -7165 17739 -7069 17773
rect 8591 17739 8687 17773
rect -16517 17547 -16483 17563
rect -16517 17454 -16483 17513
rect -8109 17547 -8075 17563
rect -16517 17262 -16483 17278
rect -16429 17454 -16395 17470
rect -16429 17262 -16395 17278
rect -14371 17454 -14337 17470
rect -14371 17262 -14337 17278
rect -12313 17454 -12279 17470
rect -12313 17262 -12279 17278
rect -10255 17454 -10221 17470
rect -10255 17262 -10221 17278
rect -8197 17454 -8163 17470
rect -8197 17262 -8163 17278
rect -8109 17454 -8075 17513
rect -8109 17262 -8075 17278
rect -15891 17185 -15875 17219
rect -14891 17185 -14875 17219
rect -13833 17185 -13817 17219
rect -12833 17185 -12817 17219
rect -11775 17185 -11759 17219
rect -10775 17185 -10759 17219
rect -9717 17185 -9701 17219
rect -8717 17185 -8701 17219
rect -15891 17034 -15875 17068
rect -14891 17034 -14875 17068
rect -13833 17034 -13817 17068
rect -12833 17034 -12817 17068
rect -11775 17034 -11759 17068
rect -10775 17034 -10759 17068
rect -9717 17034 -9701 17068
rect -8717 17034 -8701 17068
rect -16517 16975 -16483 16991
rect -16517 16783 -16483 16799
rect -16429 16975 -16395 16991
rect -16429 16783 -16395 16799
rect -14371 16975 -14337 16991
rect -14371 16783 -14337 16799
rect -12313 16975 -12279 16991
rect -12313 16783 -12279 16799
rect -10255 16975 -10221 16991
rect -10255 16783 -10221 16799
rect -8197 16975 -8163 16991
rect -8197 16783 -8163 16799
rect -8109 16975 -8075 16991
rect -8109 16783 -8075 16799
rect -15891 16706 -15875 16740
rect -14891 16706 -14875 16740
rect -13833 16706 -13817 16740
rect -12833 16706 -12817 16740
rect -11775 16706 -11759 16740
rect -10775 16706 -10759 16740
rect -9717 16706 -9701 16740
rect -8717 16706 -8701 16740
rect -16517 16669 -16483 16685
rect -16517 16619 -16483 16635
rect -8109 16669 -8075 16685
rect -8109 16619 -8075 16635
rect -15891 16564 -15875 16598
rect -14891 16564 -14875 16598
rect -13833 16564 -13817 16598
rect -12833 16564 -12817 16598
rect -11775 16564 -11759 16598
rect -10775 16564 -10759 16598
rect -9717 16564 -9701 16598
rect -8717 16564 -8701 16598
rect -16517 16505 -16483 16521
rect -16517 16313 -16483 16329
rect -16429 16505 -16395 16521
rect -16429 16313 -16395 16329
rect -14371 16505 -14337 16521
rect -14371 16313 -14337 16329
rect -12313 16505 -12279 16521
rect -12313 16313 -12279 16329
rect -10255 16505 -10221 16521
rect -10255 16313 -10221 16329
rect -8197 16505 -8163 16521
rect -8197 16313 -8163 16329
rect -8109 16505 -8075 16521
rect -8109 16313 -8075 16329
rect -15891 16236 -15875 16270
rect -14891 16236 -14875 16270
rect -13833 16236 -13817 16270
rect -12833 16236 -12817 16270
rect -11775 16236 -11759 16270
rect -10775 16236 -10759 16270
rect -9717 16236 -9701 16270
rect -8717 16236 -8701 16270
rect -15891 16085 -15875 16119
rect -14891 16085 -14875 16119
rect -13833 16085 -13817 16119
rect -12833 16085 -12817 16119
rect -11775 16085 -11759 16119
rect -10775 16085 -10759 16119
rect -9717 16085 -9701 16119
rect -8717 16085 -8701 16119
rect -16517 16026 -16483 16042
rect -16517 15791 -16483 15850
rect -16429 16026 -16395 16042
rect -16429 15834 -16395 15850
rect -14371 16026 -14337 16042
rect -14371 15834 -14337 15850
rect -12313 16026 -12279 16042
rect -12313 15834 -12279 15850
rect -10255 16026 -10221 16042
rect -10255 15834 -10221 15850
rect -8197 16026 -8163 16042
rect -8197 15834 -8163 15850
rect -8109 16026 -8075 16042
rect -16517 15741 -16483 15757
rect -8109 15791 -8075 15850
rect -8109 15741 -8075 15757
rect -7496 17453 -7462 17469
rect -7496 17360 -7462 17419
rect -3204 17453 -3170 17469
rect -7496 17168 -7462 17184
rect -7408 17360 -7374 17376
rect -7408 17168 -7374 17184
rect -5350 17360 -5316 17376
rect -5350 17168 -5316 17184
rect -3292 17360 -3258 17376
rect -3292 17168 -3258 17184
rect -3204 17360 -3170 17419
rect -3204 17168 -3170 17184
rect -6870 17091 -6854 17125
rect -5870 17091 -5854 17125
rect -4812 17091 -4796 17125
rect -3812 17091 -3796 17125
rect -7496 17021 -7462 17037
rect -7496 16928 -7462 16987
rect -3204 17021 -3170 17037
rect -7496 16736 -7462 16752
rect -7408 16928 -7374 16944
rect -7408 16736 -7374 16752
rect -5350 16928 -5316 16944
rect -5350 16736 -5316 16752
rect -3292 16928 -3258 16944
rect -3292 16736 -3258 16752
rect -3204 16928 -3170 16987
rect -3204 16736 -3170 16752
rect -6870 16659 -6854 16693
rect -5870 16659 -5854 16693
rect -4812 16659 -4796 16693
rect -3812 16659 -3796 16693
rect -6870 16517 -6854 16551
rect -5870 16517 -5854 16551
rect -4812 16517 -4796 16551
rect -3812 16517 -3796 16551
rect -7496 16458 -7462 16474
rect -7496 16223 -7462 16282
rect -7408 16458 -7374 16474
rect -7408 16266 -7374 16282
rect -5350 16458 -5316 16474
rect -5350 16266 -5316 16282
rect -3292 16458 -3258 16474
rect -3292 16266 -3258 16282
rect -3204 16458 -3170 16474
rect -7496 16173 -7462 16189
rect -3204 16223 -3170 16282
rect -3204 16173 -3170 16189
rect -6870 16085 -6854 16119
rect -5870 16085 -5854 16119
rect -4812 16085 -4796 16119
rect -3812 16085 -3796 16119
rect -7496 16026 -7462 16042
rect -7496 15791 -7462 15850
rect -7408 16026 -7374 16042
rect -7408 15834 -7374 15850
rect -5350 16026 -5316 16042
rect -5350 15834 -5316 15850
rect -3292 16026 -3258 16042
rect -3292 15834 -3258 15850
rect -3204 16026 -3170 16042
rect -7496 15741 -7462 15757
rect -3204 15791 -3170 15850
rect -3204 15741 -3170 15757
rect -1170 17524 -1136 17540
rect -478 17524 -444 17540
rect -1036 17490 -1020 17524
rect -852 17490 -836 17524
rect -778 17490 -762 17524
rect -594 17490 -578 17524
rect -1170 17440 -1136 17490
rect -1170 17248 -1136 17264
rect -1082 17440 -1048 17456
rect -1082 17248 -1048 17264
rect -824 17440 -790 17456
rect -824 17248 -790 17264
rect -566 17440 -532 17456
rect -566 17248 -532 17264
rect -478 17440 -444 17490
rect -478 17248 -444 17264
rect -1036 17180 -1020 17214
rect -852 17180 -836 17214
rect -778 17180 -762 17214
rect -594 17180 -578 17214
rect -1170 17130 -1136 17146
rect -1170 16904 -1136 16954
rect -1082 17130 -1048 17146
rect -1082 16938 -1048 16954
rect -824 17130 -790 17146
rect -824 16938 -790 16954
rect -566 17130 -532 17146
rect -566 16938 -532 16954
rect -478 17130 -444 17146
rect -478 16904 -444 16954
rect -1036 16870 -1020 16904
rect -852 16870 -836 16904
rect -778 16870 -762 16904
rect -594 16870 -578 16904
rect -1170 16854 -1136 16870
rect -478 16854 -444 16870
rect -92 17536 -58 17552
rect 8536 17536 8570 17552
rect 5316 17502 5332 17536
rect 7316 17502 7332 17536
rect -92 17452 -58 17502
rect -92 17260 -58 17276
rect -4 17452 30 17468
rect -4 17260 30 17276
rect 108 17452 142 17468
rect 108 17260 142 17276
rect 4166 17452 4200 17468
rect 4166 17260 4200 17276
rect 4278 17452 4312 17468
rect 4278 17260 4312 17276
rect 8336 17452 8370 17468
rect 8336 17260 8370 17276
rect 8448 17452 8482 17468
rect 8448 17260 8482 17276
rect 8536 17452 8570 17502
rect 8536 17260 8570 17276
rect -92 17142 -58 17158
rect -92 17058 -58 17108
rect 8536 17142 8570 17158
rect -92 16866 -58 16882
rect -4 17058 30 17074
rect -4 16866 30 16882
rect 108 17058 142 17074
rect 108 16866 142 16882
rect 4166 17058 4200 17074
rect 4166 16866 4200 16882
rect 4278 17058 4312 17074
rect 4278 16866 4312 16882
rect 8336 17058 8370 17074
rect 8336 16866 8370 16882
rect 8448 17058 8482 17074
rect 8448 16866 8482 16882
rect 8536 17058 8570 17108
rect 8536 16866 8570 16882
rect -92 16664 -58 16680
rect -92 16438 -58 16488
rect -4 16664 30 16680
rect -4 16472 30 16488
rect 108 16664 142 16680
rect 108 16472 142 16488
rect 4166 16664 4200 16680
rect 4166 16472 4200 16488
rect 4278 16664 4312 16680
rect 4278 16472 4312 16488
rect 8336 16664 8370 16680
rect 8336 16472 8370 16488
rect 8448 16664 8482 16680
rect 8448 16472 8482 16488
rect 8536 16664 8570 16680
rect -92 16388 -58 16404
rect 8536 16438 8570 16488
rect 8536 16388 8570 16404
rect -92 16270 -58 16286
rect -92 16044 -58 16094
rect -4 16270 30 16286
rect -4 16078 30 16094
rect 108 16270 142 16286
rect 108 16078 142 16094
rect 4166 16270 4200 16286
rect 4166 16078 4200 16094
rect 4278 16270 4312 16286
rect 4278 16078 4312 16094
rect 8336 16270 8370 16286
rect 8336 16078 8370 16094
rect 8448 16270 8482 16286
rect 8448 16078 8482 16094
rect 8536 16270 8570 16286
rect 8536 16044 8570 16094
rect 1146 16010 1162 16044
rect 3146 16010 3162 16044
rect -92 15994 -58 16010
rect 8536 15994 8570 16010
rect -11742 15471 -11726 15505
rect -10742 15471 -10726 15505
rect -9684 15471 -9668 15505
rect -8684 15471 -8668 15505
rect -12368 15412 -12334 15428
rect -12368 15220 -12334 15236
rect -12280 15412 -12246 15428
rect -12280 15220 -12246 15236
rect -10222 15412 -10188 15428
rect -10222 15220 -10188 15236
rect -8164 15412 -8130 15428
rect -8164 15220 -8130 15236
rect -8076 15412 -8042 15428
rect -8076 15220 -8042 15236
rect -12368 15144 -12334 15160
rect -12368 15094 -12334 15110
rect -8076 15144 -8042 15160
rect -8076 15094 -8042 15110
rect -12368 15018 -12334 15034
rect -12368 14826 -12334 14842
rect -12280 15018 -12246 15034
rect -12280 14826 -12246 14842
rect -10222 15018 -10188 15034
rect -10222 14826 -10188 14842
rect -8164 15018 -8130 15034
rect -8164 14826 -8130 14842
rect -8076 15018 -8042 15034
rect -8076 14826 -8042 14842
rect -11742 14749 -11726 14783
rect -10742 14749 -10726 14783
rect -9684 14749 -9668 14783
rect -8684 14749 -8668 14783
rect -7462 15477 -7428 15493
rect -7462 15241 -7428 15301
rect -7374 15477 -7340 15493
rect -7374 15285 -7340 15301
rect -5316 15477 -5282 15493
rect -5316 15285 -5282 15301
rect -3258 15477 -3224 15493
rect -3258 15285 -3224 15301
rect -3170 15477 -3136 15493
rect -3170 15242 -3136 15301
rect -6836 15208 -6820 15242
rect -5836 15208 -5820 15242
rect -4778 15208 -4762 15242
rect -3778 15208 -3762 15242
rect -7462 15191 -7428 15207
rect -3170 15192 -3136 15208
rect -7462 15094 -7428 15110
rect -3170 15094 -3136 15110
rect -6836 15060 -6820 15094
rect -5836 15060 -5820 15094
rect -4778 15060 -4762 15094
rect -3778 15060 -3762 15094
rect -7462 15001 -7428 15060
rect -7462 14809 -7428 14825
rect -7374 15001 -7340 15017
rect -7374 14809 -7340 14825
rect -5316 15001 -5282 15017
rect -5316 14809 -5282 14825
rect -3258 15001 -3224 15017
rect -3258 14809 -3224 14825
rect -3170 15001 -3136 15060
rect -3170 14809 -3136 14825
rect 3789 15584 3805 15618
rect 5089 15584 5105 15618
rect 6447 15584 6463 15618
rect 7747 15584 7763 15618
rect 3013 15534 3047 15550
rect 3013 15328 3047 15378
rect 3101 15534 3135 15550
rect 3101 15362 3135 15378
rect 5759 15534 5793 15550
rect 5759 15362 5793 15378
rect 8417 15534 8451 15550
rect 8417 15362 8451 15378
rect 8505 15534 8539 15550
rect 8505 15328 8539 15378
rect 3789 15294 3805 15328
rect 5089 15294 5105 15328
rect 6447 15294 6463 15328
rect 7747 15294 7763 15328
rect 3013 15278 3047 15294
rect 8505 15278 8539 15294
rect 3013 15186 3047 15202
rect 8505 15186 8539 15202
rect 3789 15152 3805 15186
rect 5089 15152 5105 15186
rect 6447 15152 6463 15186
rect 7747 15152 7763 15186
rect 3013 15102 3047 15152
rect 3013 14930 3047 14946
rect 3101 15102 3135 15118
rect 3101 14930 3135 14946
rect 5759 15102 5793 15118
rect 5759 14930 5793 14946
rect 8417 15102 8451 15118
rect 8417 14930 8451 14946
rect 8505 15102 8539 15152
rect 8505 14930 8539 14946
rect 307 12555 367 12589
rect 6341 12555 6401 12589
rect 307 12529 341 12555
rect 6367 12529 6401 12555
rect 604 12297 664 12331
rect 1470 12297 1556 12331
rect 2362 12297 2448 12331
rect 3254 12297 3340 12331
rect 4146 12297 4206 12331
rect 604 12271 638 12297
rect 1496 12271 1530 12297
rect 838 12216 854 12250
rect 1022 12216 1038 12250
rect 1096 12216 1112 12250
rect 1280 12216 1296 12250
rect 704 12166 738 12182
rect 704 11374 738 11390
rect 792 12166 826 12182
rect 792 11374 826 11390
rect 1050 12166 1084 12182
rect 1050 11374 1084 11390
rect 1308 12166 1342 12182
rect 1308 11374 1342 11390
rect 1396 12166 1430 12182
rect 1396 11374 1430 11390
rect 704 11298 738 11314
rect 704 11248 738 11264
rect 1396 11298 1430 11314
rect 1396 11248 1430 11264
rect 704 11172 738 11188
rect 704 10380 738 10396
rect 792 11172 826 11188
rect 792 10380 826 10396
rect 1050 11172 1084 11188
rect 1050 10380 1084 10396
rect 1308 11172 1342 11188
rect 1308 10380 1342 10396
rect 1396 11172 1430 11188
rect 1396 10380 1430 10396
rect 838 10312 854 10346
rect 1022 10312 1038 10346
rect 1096 10312 1112 10346
rect 1280 10312 1296 10346
rect 604 10265 638 10291
rect 2388 12271 2422 12297
rect 1730 12216 1746 12250
rect 1914 12216 1930 12250
rect 1988 12216 2004 12250
rect 2172 12216 2188 12250
rect 1596 12166 1630 12182
rect 1596 11374 1630 11390
rect 1684 12166 1718 12182
rect 1684 11374 1718 11390
rect 1942 12166 1976 12182
rect 1942 11374 1976 11390
rect 2200 12166 2234 12182
rect 2200 11374 2234 11390
rect 2288 12166 2322 12182
rect 2288 11374 2322 11390
rect 1596 11298 1630 11314
rect 1596 11248 1630 11264
rect 2288 11298 2322 11314
rect 2288 11248 2322 11264
rect 1596 11172 1630 11188
rect 1596 10380 1630 10396
rect 1684 11172 1718 11188
rect 1684 10380 1718 10396
rect 1942 11172 1976 11188
rect 1942 10380 1976 10396
rect 2200 11172 2234 11188
rect 2200 10380 2234 10396
rect 2288 11172 2322 11188
rect 2288 10380 2322 10396
rect 1730 10312 1746 10346
rect 1914 10312 1930 10346
rect 1988 10312 2004 10346
rect 2172 10312 2188 10346
rect 1496 10265 1530 10291
rect 3280 12271 3314 12297
rect 2622 12216 2638 12250
rect 2806 12216 2822 12250
rect 2880 12216 2896 12250
rect 3064 12216 3080 12250
rect 2488 12166 2522 12182
rect 2488 11374 2522 11390
rect 2576 12166 2610 12182
rect 2576 11374 2610 11390
rect 2834 12166 2868 12182
rect 2834 11374 2868 11390
rect 3092 12166 3126 12182
rect 3092 11374 3126 11390
rect 3180 12166 3214 12182
rect 3180 11374 3214 11390
rect 2488 11298 2522 11314
rect 2488 11248 2522 11264
rect 3180 11298 3214 11314
rect 3180 11248 3214 11264
rect 2488 11172 2522 11188
rect 2488 10380 2522 10396
rect 2576 11172 2610 11188
rect 2576 10380 2610 10396
rect 2834 11172 2868 11188
rect 2834 10380 2868 10396
rect 3092 11172 3126 11188
rect 3092 10380 3126 10396
rect 3180 11172 3214 11188
rect 3180 10380 3214 10396
rect 2622 10312 2638 10346
rect 2806 10312 2822 10346
rect 2880 10312 2896 10346
rect 3064 10312 3080 10346
rect 2388 10265 2422 10291
rect 4172 12271 4206 12297
rect 3514 12216 3530 12250
rect 3698 12216 3714 12250
rect 3772 12216 3788 12250
rect 3956 12216 3972 12250
rect 3380 12166 3414 12182
rect 3380 11374 3414 11390
rect 3468 12166 3502 12182
rect 3468 11374 3502 11390
rect 3726 12166 3760 12182
rect 3726 11374 3760 11390
rect 3984 12166 4018 12182
rect 3984 11374 4018 11390
rect 4072 12166 4106 12182
rect 4072 11374 4106 11390
rect 3380 11298 3414 11314
rect 3380 11248 3414 11264
rect 4072 11298 4106 11314
rect 4072 11248 4106 11264
rect 3380 11172 3414 11188
rect 3380 10380 3414 10396
rect 3468 11172 3502 11188
rect 3468 10380 3502 10396
rect 3726 11172 3760 11188
rect 3726 10380 3760 10396
rect 3984 11172 4018 11188
rect 3984 10380 4018 10396
rect 4072 11172 4106 11188
rect 4072 10380 4106 10396
rect 3514 10312 3530 10346
rect 3698 10312 3714 10346
rect 3772 10312 3788 10346
rect 3956 10312 3972 10346
rect 3280 10265 3314 10291
rect 4260 12267 4320 12301
rect 4712 12267 4772 12301
rect 4260 12241 4294 12267
rect 4738 12241 4772 12267
rect 4328 12167 4344 12201
rect 4378 12167 4428 12201
rect 4604 12167 4620 12201
rect 4412 12079 4428 12113
rect 4604 12079 4620 12113
rect 4654 12051 4688 12067
rect 4654 11867 4688 11883
rect 4412 11821 4428 11855
rect 4604 11821 4620 11855
rect 4654 11793 4688 11809
rect 4654 11609 4688 11625
rect 4412 11563 4428 11597
rect 4604 11563 4620 11597
rect 4328 11475 4344 11509
rect 4378 11475 4428 11509
rect 4604 11475 4620 11509
rect 4260 11409 4294 11435
rect 4738 11409 4772 11435
rect 4260 11375 4320 11409
rect 4712 11375 4772 11409
rect 4836 11878 4896 11912
rect 6076 11878 6136 11912
rect 4836 11852 4870 11878
rect 4172 10265 4206 10291
rect 604 10231 664 10265
rect 1470 10231 1556 10265
rect 2362 10231 2448 10265
rect 3254 10231 3340 10265
rect 4146 10231 4206 10265
rect 4260 11153 4320 11187
rect 4712 11153 4772 11187
rect 4260 11127 4294 11153
rect 4738 11127 4772 11153
rect 4328 11053 4344 11087
rect 4378 11053 4428 11087
rect 4604 11053 4620 11087
rect 4412 10965 4428 10999
rect 4604 10965 4620 10999
rect 4654 10937 4688 10953
rect 4654 10753 4688 10769
rect 4412 10707 4428 10741
rect 4604 10707 4620 10741
rect 4654 10679 4688 10695
rect 4654 10495 4688 10511
rect 4412 10449 4428 10483
rect 4604 10449 4620 10483
rect 4328 10361 4344 10395
rect 4378 10361 4428 10395
rect 4604 10361 4620 10395
rect 4260 10295 4294 10321
rect 6102 11852 6136 11878
rect 4985 11778 5001 11812
rect 5377 11778 5393 11812
rect 5453 11778 5469 11812
rect 5503 11778 5519 11812
rect 5579 11778 5595 11812
rect 5971 11778 5987 11812
rect 4985 11690 5001 11724
rect 5377 11690 5393 11724
rect 5579 11690 5595 11724
rect 5971 11690 5987 11724
rect 4908 11570 4942 11586
rect 4908 11370 4942 11386
rect 6030 11570 6064 11586
rect 6030 11370 6064 11386
rect 4985 11232 5001 11266
rect 5377 11232 5393 11266
rect 5579 11232 5595 11266
rect 5971 11232 5987 11266
rect 4908 11112 4942 11128
rect 4908 10912 4942 10928
rect 6030 11112 6064 11128
rect 6030 10912 6064 10928
rect 4985 10774 5001 10808
rect 5377 10774 5393 10808
rect 5579 10774 5595 10808
rect 5971 10774 5987 10808
rect 4985 10686 5001 10720
rect 5377 10686 5393 10720
rect 5453 10686 5469 10720
rect 5503 10686 5519 10720
rect 5579 10686 5595 10720
rect 5971 10686 5987 10720
rect 4836 10620 4870 10646
rect 6102 10620 6136 10646
rect 4836 10586 4896 10620
rect 6076 10586 6136 10620
rect 4738 10295 4772 10321
rect 4260 10261 4320 10295
rect 4712 10261 4772 10295
rect 307 10007 341 10033
rect 6367 10007 6401 10033
rect 307 9973 367 10007
rect 6341 9973 6401 10007
rect 329 8373 1617 8406
rect 329 8339 387 8373
rect 421 8339 477 8373
rect 511 8339 567 8373
rect 601 8339 657 8373
rect 691 8339 747 8373
rect 781 8339 837 8373
rect 871 8339 927 8373
rect 961 8339 1017 8373
rect 1051 8339 1107 8373
rect 1141 8339 1197 8373
rect 1231 8339 1287 8373
rect 1321 8339 1377 8373
rect 1411 8339 1467 8373
rect 1501 8339 1617 8373
rect 329 8307 1617 8339
rect 329 8272 428 8307
rect 329 8238 364 8272
rect 398 8238 428 8272
rect 1518 8272 1617 8307
rect 329 8182 428 8238
rect 329 8148 364 8182
rect 398 8148 428 8182
rect 329 8092 428 8148
rect 329 8058 364 8092
rect 398 8058 428 8092
rect 329 8002 428 8058
rect 329 7968 364 8002
rect 398 7968 428 8002
rect 329 7912 428 7968
rect 329 7878 364 7912
rect 398 7878 428 7912
rect 329 7822 428 7878
rect 329 7788 364 7822
rect 398 7788 428 7822
rect 329 7732 428 7788
rect 329 7698 364 7732
rect 398 7698 428 7732
rect 329 7642 428 7698
rect 329 7608 364 7642
rect 398 7608 428 7642
rect 329 7552 428 7608
rect 329 7518 364 7552
rect 398 7518 428 7552
rect 329 7462 428 7518
rect 329 7428 364 7462
rect 398 7428 428 7462
rect 329 7372 428 7428
rect 329 7338 364 7372
rect 398 7338 428 7372
rect 329 7282 428 7338
rect 329 7248 364 7282
rect 398 7248 428 7282
rect 492 8224 1454 8243
rect 492 8190 587 8224
rect 621 8190 677 8224
rect 711 8190 767 8224
rect 801 8190 857 8224
rect 891 8190 947 8224
rect 981 8190 1037 8224
rect 1071 8190 1127 8224
rect 1161 8190 1217 8224
rect 1251 8190 1307 8224
rect 1341 8190 1454 8224
rect 492 8171 1454 8190
rect 492 8166 564 8171
rect 492 8132 511 8166
rect 545 8132 564 8166
rect 492 8076 564 8132
rect 1382 8132 1454 8171
rect 492 8042 511 8076
rect 545 8042 564 8076
rect 492 7986 564 8042
rect 492 7952 511 7986
rect 545 7952 564 7986
rect 492 7896 564 7952
rect 492 7862 511 7896
rect 545 7862 564 7896
rect 492 7806 564 7862
rect 492 7772 511 7806
rect 545 7772 564 7806
rect 492 7716 564 7772
rect 492 7682 511 7716
rect 545 7682 564 7716
rect 492 7626 564 7682
rect 492 7592 511 7626
rect 545 7592 564 7626
rect 492 7536 564 7592
rect 492 7502 511 7536
rect 545 7502 564 7536
rect 492 7446 564 7502
rect 492 7412 511 7446
rect 545 7412 564 7446
rect 626 8050 1320 8109
rect 626 8016 685 8050
rect 719 8022 775 8050
rect 747 8016 775 8022
rect 809 8022 865 8050
rect 809 8016 813 8022
rect 626 7988 713 8016
rect 747 7988 813 8016
rect 847 8016 865 8022
rect 899 8022 955 8050
rect 899 8016 913 8022
rect 847 7988 913 8016
rect 947 8016 955 8022
rect 989 8022 1045 8050
rect 1079 8022 1135 8050
rect 1169 8022 1225 8050
rect 989 8016 1013 8022
rect 1079 8016 1113 8022
rect 1169 8016 1213 8022
rect 1259 8016 1320 8050
rect 947 7988 1013 8016
rect 1047 7988 1113 8016
rect 1147 7988 1213 8016
rect 1247 7988 1320 8016
rect 626 7960 1320 7988
rect 626 7926 685 7960
rect 719 7926 775 7960
rect 809 7926 865 7960
rect 899 7926 955 7960
rect 989 7926 1045 7960
rect 1079 7926 1135 7960
rect 1169 7926 1225 7960
rect 1259 7926 1320 7960
rect 626 7922 1320 7926
rect 626 7888 713 7922
rect 747 7888 813 7922
rect 847 7888 913 7922
rect 947 7888 1013 7922
rect 1047 7888 1113 7922
rect 1147 7888 1213 7922
rect 1247 7888 1320 7922
rect 626 7870 1320 7888
rect 626 7836 685 7870
rect 719 7836 775 7870
rect 809 7836 865 7870
rect 899 7836 955 7870
rect 989 7836 1045 7870
rect 1079 7836 1135 7870
rect 1169 7836 1225 7870
rect 1259 7836 1320 7870
rect 626 7822 1320 7836
rect 626 7788 713 7822
rect 747 7788 813 7822
rect 847 7788 913 7822
rect 947 7788 1013 7822
rect 1047 7788 1113 7822
rect 1147 7788 1213 7822
rect 1247 7788 1320 7822
rect 626 7780 1320 7788
rect 626 7746 685 7780
rect 719 7746 775 7780
rect 809 7746 865 7780
rect 899 7746 955 7780
rect 989 7746 1045 7780
rect 1079 7746 1135 7780
rect 1169 7746 1225 7780
rect 1259 7746 1320 7780
rect 626 7722 1320 7746
rect 626 7690 713 7722
rect 747 7690 813 7722
rect 626 7656 685 7690
rect 747 7688 775 7690
rect 719 7656 775 7688
rect 809 7688 813 7690
rect 847 7690 913 7722
rect 847 7688 865 7690
rect 809 7656 865 7688
rect 899 7688 913 7690
rect 947 7690 1013 7722
rect 1047 7690 1113 7722
rect 1147 7690 1213 7722
rect 1247 7690 1320 7722
rect 947 7688 955 7690
rect 899 7656 955 7688
rect 989 7688 1013 7690
rect 1079 7688 1113 7690
rect 1169 7688 1213 7690
rect 989 7656 1045 7688
rect 1079 7656 1135 7688
rect 1169 7656 1225 7688
rect 1259 7656 1320 7690
rect 626 7622 1320 7656
rect 626 7600 713 7622
rect 747 7600 813 7622
rect 626 7566 685 7600
rect 747 7588 775 7600
rect 719 7566 775 7588
rect 809 7588 813 7600
rect 847 7600 913 7622
rect 847 7588 865 7600
rect 809 7566 865 7588
rect 899 7588 913 7600
rect 947 7600 1013 7622
rect 1047 7600 1113 7622
rect 1147 7600 1213 7622
rect 1247 7600 1320 7622
rect 947 7588 955 7600
rect 899 7566 955 7588
rect 989 7588 1013 7600
rect 1079 7588 1113 7600
rect 1169 7588 1213 7600
rect 989 7566 1045 7588
rect 1079 7566 1135 7588
rect 1169 7566 1225 7588
rect 1259 7566 1320 7600
rect 626 7522 1320 7566
rect 626 7510 713 7522
rect 747 7510 813 7522
rect 626 7476 685 7510
rect 747 7488 775 7510
rect 719 7476 775 7488
rect 809 7488 813 7510
rect 847 7510 913 7522
rect 847 7488 865 7510
rect 809 7476 865 7488
rect 899 7488 913 7510
rect 947 7510 1013 7522
rect 1047 7510 1113 7522
rect 1147 7510 1213 7522
rect 1247 7510 1320 7522
rect 947 7488 955 7510
rect 899 7476 955 7488
rect 989 7488 1013 7510
rect 1079 7488 1113 7510
rect 1169 7488 1213 7510
rect 989 7476 1045 7488
rect 1079 7476 1135 7488
rect 1169 7476 1225 7488
rect 1259 7476 1320 7510
rect 626 7415 1320 7476
rect 1382 8098 1401 8132
rect 1435 8098 1454 8132
rect 1382 8042 1454 8098
rect 1382 8008 1401 8042
rect 1435 8008 1454 8042
rect 1382 7952 1454 8008
rect 1382 7918 1401 7952
rect 1435 7918 1454 7952
rect 1382 7862 1454 7918
rect 1382 7828 1401 7862
rect 1435 7828 1454 7862
rect 1382 7772 1454 7828
rect 1382 7738 1401 7772
rect 1435 7738 1454 7772
rect 1382 7682 1454 7738
rect 1382 7648 1401 7682
rect 1435 7648 1454 7682
rect 1382 7592 1454 7648
rect 1382 7558 1401 7592
rect 1435 7558 1454 7592
rect 1382 7502 1454 7558
rect 1382 7468 1401 7502
rect 1435 7468 1454 7502
rect 492 7353 564 7412
rect 1382 7412 1454 7468
rect 1382 7378 1401 7412
rect 1435 7378 1454 7412
rect 1382 7353 1454 7378
rect 492 7334 1382 7353
rect 492 7300 568 7334
rect 602 7300 658 7334
rect 692 7300 748 7334
rect 782 7300 838 7334
rect 872 7300 928 7334
rect 962 7300 1018 7334
rect 1052 7300 1108 7334
rect 1142 7300 1198 7334
rect 1232 7300 1288 7334
rect 1322 7300 1382 7334
rect 492 7281 1382 7300
rect 1518 8238 1551 8272
rect 1585 8238 1617 8272
rect 1518 8182 1617 8238
rect 1518 8148 1551 8182
rect 1585 8148 1617 8182
rect 1518 8092 1617 8148
rect 1518 8058 1551 8092
rect 1585 8058 1617 8092
rect 1518 8002 1617 8058
rect 1518 7968 1551 8002
rect 1585 7968 1617 8002
rect 1518 7912 1617 7968
rect 1518 7878 1551 7912
rect 1585 7878 1617 7912
rect 1518 7822 1617 7878
rect 1518 7788 1551 7822
rect 1585 7788 1617 7822
rect 1518 7732 1617 7788
rect 1518 7698 1551 7732
rect 1585 7698 1617 7732
rect 1518 7642 1617 7698
rect 1518 7608 1551 7642
rect 1585 7608 1617 7642
rect 1518 7552 1617 7608
rect 1518 7518 1551 7552
rect 1585 7518 1617 7552
rect 1518 7462 1617 7518
rect 1518 7428 1551 7462
rect 1585 7428 1617 7462
rect 1518 7372 1617 7428
rect 1518 7353 1551 7372
rect 1585 7353 1617 7372
rect 329 7217 428 7248
rect 1518 7248 1551 7281
rect 1585 7248 1617 7281
rect 1518 7217 1617 7248
rect 329 7186 1382 7217
rect 1454 7186 1617 7217
rect 329 7152 387 7186
rect 421 7152 477 7186
rect 511 7152 567 7186
rect 601 7152 657 7186
rect 691 7152 747 7186
rect 781 7152 837 7186
rect 871 7152 927 7186
rect 961 7152 1017 7186
rect 1051 7152 1107 7186
rect 1141 7152 1197 7186
rect 1231 7152 1287 7186
rect 1321 7152 1377 7186
rect 1454 7152 1467 7186
rect 1501 7152 1617 7186
rect 329 7118 1382 7152
rect 1454 7118 1617 7152
rect 1717 8373 3005 8406
rect 1717 8339 1775 8373
rect 1809 8339 1865 8373
rect 1899 8339 1955 8373
rect 1989 8339 2045 8373
rect 2079 8339 2135 8373
rect 2169 8339 2225 8373
rect 2259 8339 2315 8373
rect 2349 8339 2405 8373
rect 2439 8339 2495 8373
rect 2529 8339 2585 8373
rect 2619 8339 2675 8373
rect 2709 8339 2765 8373
rect 2799 8339 2855 8373
rect 2889 8339 3005 8373
rect 1717 8307 3005 8339
rect 1717 8272 1816 8307
rect 1717 8238 1752 8272
rect 1786 8238 1816 8272
rect 2906 8272 3005 8307
rect 1717 8182 1816 8238
rect 1717 8148 1752 8182
rect 1786 8148 1816 8182
rect 1717 8092 1816 8148
rect 1717 8058 1752 8092
rect 1786 8058 1816 8092
rect 1717 8002 1816 8058
rect 1717 7968 1752 8002
rect 1786 7968 1816 8002
rect 1717 7912 1816 7968
rect 1717 7878 1752 7912
rect 1786 7878 1816 7912
rect 1717 7822 1816 7878
rect 1717 7788 1752 7822
rect 1786 7788 1816 7822
rect 1717 7732 1816 7788
rect 1717 7698 1752 7732
rect 1786 7698 1816 7732
rect 1717 7642 1816 7698
rect 1717 7608 1752 7642
rect 1786 7608 1816 7642
rect 1717 7552 1816 7608
rect 1717 7518 1752 7552
rect 1786 7518 1816 7552
rect 1717 7462 1816 7518
rect 1717 7428 1752 7462
rect 1786 7428 1816 7462
rect 1717 7372 1816 7428
rect 1717 7338 1752 7372
rect 1786 7338 1816 7372
rect 1717 7282 1816 7338
rect 1717 7248 1752 7282
rect 1786 7248 1816 7282
rect 1880 8224 2842 8243
rect 1880 8190 1975 8224
rect 2009 8190 2065 8224
rect 2099 8190 2155 8224
rect 2189 8190 2245 8224
rect 2279 8190 2335 8224
rect 2369 8190 2425 8224
rect 2459 8190 2515 8224
rect 2549 8190 2605 8224
rect 2639 8190 2695 8224
rect 2729 8190 2842 8224
rect 1880 8171 2842 8190
rect 1880 8166 1952 8171
rect 1880 8132 1899 8166
rect 1933 8132 1952 8166
rect 1880 8076 1952 8132
rect 2770 8132 2842 8171
rect 1880 8042 1899 8076
rect 1933 8042 1952 8076
rect 1880 7986 1952 8042
rect 1880 7952 1899 7986
rect 1933 7952 1952 7986
rect 1880 7896 1952 7952
rect 1880 7862 1899 7896
rect 1933 7862 1952 7896
rect 1880 7806 1952 7862
rect 1880 7772 1899 7806
rect 1933 7772 1952 7806
rect 1880 7716 1952 7772
rect 1880 7682 1899 7716
rect 1933 7682 1952 7716
rect 1880 7626 1952 7682
rect 1880 7592 1899 7626
rect 1933 7592 1952 7626
rect 1880 7536 1952 7592
rect 1880 7502 1899 7536
rect 1933 7502 1952 7536
rect 1880 7446 1952 7502
rect 1880 7412 1899 7446
rect 1933 7412 1952 7446
rect 2014 8050 2708 8109
rect 2014 8016 2073 8050
rect 2107 8022 2163 8050
rect 2135 8016 2163 8022
rect 2197 8022 2253 8050
rect 2197 8016 2201 8022
rect 2014 7988 2101 8016
rect 2135 7988 2201 8016
rect 2235 8016 2253 8022
rect 2287 8022 2343 8050
rect 2287 8016 2301 8022
rect 2235 7988 2301 8016
rect 2335 8016 2343 8022
rect 2377 8022 2433 8050
rect 2467 8022 2523 8050
rect 2557 8022 2613 8050
rect 2377 8016 2401 8022
rect 2467 8016 2501 8022
rect 2557 8016 2601 8022
rect 2647 8016 2708 8050
rect 2335 7988 2401 8016
rect 2435 7988 2501 8016
rect 2535 7988 2601 8016
rect 2635 7988 2708 8016
rect 2014 7960 2708 7988
rect 2014 7926 2073 7960
rect 2107 7926 2163 7960
rect 2197 7926 2253 7960
rect 2287 7926 2343 7960
rect 2377 7926 2433 7960
rect 2467 7926 2523 7960
rect 2557 7926 2613 7960
rect 2647 7926 2708 7960
rect 2014 7922 2708 7926
rect 2014 7888 2101 7922
rect 2135 7888 2201 7922
rect 2235 7888 2301 7922
rect 2335 7888 2401 7922
rect 2435 7888 2501 7922
rect 2535 7888 2601 7922
rect 2635 7888 2708 7922
rect 2014 7870 2708 7888
rect 2014 7836 2073 7870
rect 2107 7836 2163 7870
rect 2197 7836 2253 7870
rect 2287 7836 2343 7870
rect 2377 7836 2433 7870
rect 2467 7836 2523 7870
rect 2557 7836 2613 7870
rect 2647 7836 2708 7870
rect 2014 7822 2708 7836
rect 2014 7788 2101 7822
rect 2135 7788 2201 7822
rect 2235 7788 2301 7822
rect 2335 7788 2401 7822
rect 2435 7788 2501 7822
rect 2535 7788 2601 7822
rect 2635 7788 2708 7822
rect 2014 7780 2708 7788
rect 2014 7746 2073 7780
rect 2107 7746 2163 7780
rect 2197 7746 2253 7780
rect 2287 7746 2343 7780
rect 2377 7746 2433 7780
rect 2467 7746 2523 7780
rect 2557 7746 2613 7780
rect 2647 7746 2708 7780
rect 2014 7722 2708 7746
rect 2014 7690 2101 7722
rect 2135 7690 2201 7722
rect 2014 7656 2073 7690
rect 2135 7688 2163 7690
rect 2107 7656 2163 7688
rect 2197 7688 2201 7690
rect 2235 7690 2301 7722
rect 2235 7688 2253 7690
rect 2197 7656 2253 7688
rect 2287 7688 2301 7690
rect 2335 7690 2401 7722
rect 2435 7690 2501 7722
rect 2535 7690 2601 7722
rect 2635 7690 2708 7722
rect 2335 7688 2343 7690
rect 2287 7656 2343 7688
rect 2377 7688 2401 7690
rect 2467 7688 2501 7690
rect 2557 7688 2601 7690
rect 2377 7656 2433 7688
rect 2467 7656 2523 7688
rect 2557 7656 2613 7688
rect 2647 7656 2708 7690
rect 2014 7622 2708 7656
rect 2014 7600 2101 7622
rect 2135 7600 2201 7622
rect 2014 7566 2073 7600
rect 2135 7588 2163 7600
rect 2107 7566 2163 7588
rect 2197 7588 2201 7600
rect 2235 7600 2301 7622
rect 2235 7588 2253 7600
rect 2197 7566 2253 7588
rect 2287 7588 2301 7600
rect 2335 7600 2401 7622
rect 2435 7600 2501 7622
rect 2535 7600 2601 7622
rect 2635 7600 2708 7622
rect 2335 7588 2343 7600
rect 2287 7566 2343 7588
rect 2377 7588 2401 7600
rect 2467 7588 2501 7600
rect 2557 7588 2601 7600
rect 2377 7566 2433 7588
rect 2467 7566 2523 7588
rect 2557 7566 2613 7588
rect 2647 7566 2708 7600
rect 2014 7522 2708 7566
rect 2014 7510 2101 7522
rect 2135 7510 2201 7522
rect 2014 7476 2073 7510
rect 2135 7488 2163 7510
rect 2107 7476 2163 7488
rect 2197 7488 2201 7510
rect 2235 7510 2301 7522
rect 2235 7488 2253 7510
rect 2197 7476 2253 7488
rect 2287 7488 2301 7510
rect 2335 7510 2401 7522
rect 2435 7510 2501 7522
rect 2535 7510 2601 7522
rect 2635 7510 2708 7522
rect 2335 7488 2343 7510
rect 2287 7476 2343 7488
rect 2377 7488 2401 7510
rect 2467 7488 2501 7510
rect 2557 7488 2601 7510
rect 2377 7476 2433 7488
rect 2467 7476 2523 7488
rect 2557 7476 2613 7488
rect 2647 7476 2708 7510
rect 2014 7415 2708 7476
rect 2770 8098 2789 8132
rect 2823 8098 2842 8132
rect 2770 8042 2842 8098
rect 2770 8008 2789 8042
rect 2823 8008 2842 8042
rect 2770 7952 2842 8008
rect 2770 7918 2789 7952
rect 2823 7918 2842 7952
rect 2770 7862 2842 7918
rect 2770 7828 2789 7862
rect 2823 7828 2842 7862
rect 2770 7772 2842 7828
rect 2770 7738 2789 7772
rect 2823 7738 2842 7772
rect 2770 7682 2842 7738
rect 2770 7648 2789 7682
rect 2823 7648 2842 7682
rect 2770 7592 2842 7648
rect 2770 7558 2789 7592
rect 2823 7558 2842 7592
rect 2770 7502 2842 7558
rect 2770 7468 2789 7502
rect 2823 7468 2842 7502
rect 1880 7353 1952 7412
rect 2770 7412 2842 7468
rect 2770 7378 2789 7412
rect 2823 7378 2842 7412
rect 2770 7353 2842 7378
rect 1880 7334 2770 7353
rect 1880 7300 1956 7334
rect 1990 7300 2046 7334
rect 2080 7300 2136 7334
rect 2170 7300 2226 7334
rect 2260 7300 2316 7334
rect 2350 7300 2406 7334
rect 2440 7300 2496 7334
rect 2530 7300 2586 7334
rect 2620 7300 2676 7334
rect 2710 7300 2770 7334
rect 1880 7281 2770 7300
rect 2906 8238 2939 8272
rect 2973 8238 3005 8272
rect 2906 8182 3005 8238
rect 2906 8148 2939 8182
rect 2973 8148 3005 8182
rect 2906 8092 3005 8148
rect 2906 8058 2939 8092
rect 2973 8058 3005 8092
rect 2906 8002 3005 8058
rect 2906 7968 2939 8002
rect 2973 7968 3005 8002
rect 2906 7912 3005 7968
rect 2906 7878 2939 7912
rect 2973 7878 3005 7912
rect 2906 7822 3005 7878
rect 2906 7788 2939 7822
rect 2973 7788 3005 7822
rect 2906 7732 3005 7788
rect 2906 7698 2939 7732
rect 2973 7698 3005 7732
rect 2906 7642 3005 7698
rect 2906 7608 2939 7642
rect 2973 7608 3005 7642
rect 2906 7552 3005 7608
rect 2906 7518 2939 7552
rect 2973 7518 3005 7552
rect 2906 7462 3005 7518
rect 2906 7428 2939 7462
rect 2973 7428 3005 7462
rect 2906 7372 3005 7428
rect 2906 7353 2939 7372
rect 2973 7353 3005 7372
rect 1717 7217 1816 7248
rect 2906 7248 2939 7281
rect 2973 7248 3005 7281
rect 2906 7217 3005 7248
rect 1717 7186 3005 7217
rect 1717 7152 1775 7186
rect 1809 7152 1865 7186
rect 1899 7152 1955 7186
rect 1989 7152 2045 7186
rect 2079 7152 2135 7186
rect 2169 7152 2225 7186
rect 2259 7152 2315 7186
rect 2349 7152 2405 7186
rect 2439 7152 2495 7186
rect 2529 7152 2585 7186
rect 2619 7152 2675 7186
rect 2709 7152 2765 7186
rect 2799 7152 2855 7186
rect 2889 7152 3005 7186
rect 1717 7118 3005 7152
rect 3105 8373 4393 8406
rect 3105 8339 3163 8373
rect 3197 8339 3253 8373
rect 3287 8339 3343 8373
rect 3377 8339 3433 8373
rect 3467 8339 3523 8373
rect 3557 8339 3613 8373
rect 3647 8339 3703 8373
rect 3737 8339 3793 8373
rect 3827 8339 3883 8373
rect 3917 8339 3973 8373
rect 4007 8339 4063 8373
rect 4097 8339 4153 8373
rect 4187 8339 4243 8373
rect 4277 8339 4393 8373
rect 3105 8307 4393 8339
rect 3105 8272 3204 8307
rect 3105 8238 3140 8272
rect 3174 8238 3204 8272
rect 4294 8272 4393 8307
rect 3105 8182 3204 8238
rect 3105 8148 3140 8182
rect 3174 8148 3204 8182
rect 3105 8092 3204 8148
rect 3105 8058 3140 8092
rect 3174 8058 3204 8092
rect 3105 8002 3204 8058
rect 3105 7968 3140 8002
rect 3174 7968 3204 8002
rect 3105 7912 3204 7968
rect 3105 7878 3140 7912
rect 3174 7878 3204 7912
rect 3105 7822 3204 7878
rect 3105 7788 3140 7822
rect 3174 7788 3204 7822
rect 3105 7732 3204 7788
rect 3105 7698 3140 7732
rect 3174 7698 3204 7732
rect 3105 7642 3204 7698
rect 3105 7608 3140 7642
rect 3174 7608 3204 7642
rect 3105 7552 3204 7608
rect 3105 7518 3140 7552
rect 3174 7518 3204 7552
rect 3105 7462 3204 7518
rect 3105 7428 3140 7462
rect 3174 7428 3204 7462
rect 3105 7372 3204 7428
rect 3105 7353 3140 7372
rect 3174 7353 3204 7372
rect 3268 8224 4230 8243
rect 3268 8190 3363 8224
rect 3397 8190 3453 8224
rect 3487 8190 3543 8224
rect 3577 8190 3633 8224
rect 3667 8190 3723 8224
rect 3757 8190 3813 8224
rect 3847 8190 3903 8224
rect 3937 8190 3993 8224
rect 4027 8190 4083 8224
rect 4117 8190 4230 8224
rect 3268 8171 4230 8190
rect 3268 8166 3340 8171
rect 3268 8132 3287 8166
rect 3321 8132 3340 8166
rect 3268 8076 3340 8132
rect 4158 8132 4230 8171
rect 3268 8042 3287 8076
rect 3321 8042 3340 8076
rect 3268 7986 3340 8042
rect 3268 7952 3287 7986
rect 3321 7952 3340 7986
rect 3268 7896 3340 7952
rect 3268 7862 3287 7896
rect 3321 7862 3340 7896
rect 3268 7806 3340 7862
rect 3268 7772 3287 7806
rect 3321 7772 3340 7806
rect 3268 7716 3340 7772
rect 3268 7682 3287 7716
rect 3321 7682 3340 7716
rect 3268 7626 3340 7682
rect 3268 7592 3287 7626
rect 3321 7592 3340 7626
rect 3268 7536 3340 7592
rect 3268 7502 3287 7536
rect 3321 7502 3340 7536
rect 3268 7446 3340 7502
rect 3268 7412 3287 7446
rect 3321 7412 3340 7446
rect 3402 8050 4096 8109
rect 3402 8016 3461 8050
rect 3495 8022 3551 8050
rect 3523 8016 3551 8022
rect 3585 8022 3641 8050
rect 3585 8016 3589 8022
rect 3402 7988 3489 8016
rect 3523 7988 3589 8016
rect 3623 8016 3641 8022
rect 3675 8022 3731 8050
rect 3675 8016 3689 8022
rect 3623 7988 3689 8016
rect 3723 8016 3731 8022
rect 3765 8022 3821 8050
rect 3855 8022 3911 8050
rect 3945 8022 4001 8050
rect 3765 8016 3789 8022
rect 3855 8016 3889 8022
rect 3945 8016 3989 8022
rect 4035 8016 4096 8050
rect 3723 7988 3789 8016
rect 3823 7988 3889 8016
rect 3923 7988 3989 8016
rect 4023 7988 4096 8016
rect 3402 7960 4096 7988
rect 3402 7926 3461 7960
rect 3495 7926 3551 7960
rect 3585 7926 3641 7960
rect 3675 7926 3731 7960
rect 3765 7926 3821 7960
rect 3855 7926 3911 7960
rect 3945 7926 4001 7960
rect 4035 7926 4096 7960
rect 3402 7922 4096 7926
rect 3402 7888 3489 7922
rect 3523 7888 3589 7922
rect 3623 7888 3689 7922
rect 3723 7888 3789 7922
rect 3823 7888 3889 7922
rect 3923 7888 3989 7922
rect 4023 7888 4096 7922
rect 3402 7870 4096 7888
rect 3402 7836 3461 7870
rect 3495 7836 3551 7870
rect 3585 7836 3641 7870
rect 3675 7836 3731 7870
rect 3765 7836 3821 7870
rect 3855 7836 3911 7870
rect 3945 7836 4001 7870
rect 4035 7836 4096 7870
rect 3402 7822 4096 7836
rect 3402 7788 3489 7822
rect 3523 7788 3589 7822
rect 3623 7788 3689 7822
rect 3723 7788 3789 7822
rect 3823 7788 3889 7822
rect 3923 7788 3989 7822
rect 4023 7788 4096 7822
rect 3402 7780 4096 7788
rect 3402 7746 3461 7780
rect 3495 7746 3551 7780
rect 3585 7746 3641 7780
rect 3675 7746 3731 7780
rect 3765 7746 3821 7780
rect 3855 7746 3911 7780
rect 3945 7746 4001 7780
rect 4035 7746 4096 7780
rect 3402 7722 4096 7746
rect 3402 7690 3489 7722
rect 3523 7690 3589 7722
rect 3402 7656 3461 7690
rect 3523 7688 3551 7690
rect 3495 7656 3551 7688
rect 3585 7688 3589 7690
rect 3623 7690 3689 7722
rect 3623 7688 3641 7690
rect 3585 7656 3641 7688
rect 3675 7688 3689 7690
rect 3723 7690 3789 7722
rect 3823 7690 3889 7722
rect 3923 7690 3989 7722
rect 4023 7690 4096 7722
rect 3723 7688 3731 7690
rect 3675 7656 3731 7688
rect 3765 7688 3789 7690
rect 3855 7688 3889 7690
rect 3945 7688 3989 7690
rect 3765 7656 3821 7688
rect 3855 7656 3911 7688
rect 3945 7656 4001 7688
rect 4035 7656 4096 7690
rect 3402 7622 4096 7656
rect 3402 7600 3489 7622
rect 3523 7600 3589 7622
rect 3402 7566 3461 7600
rect 3523 7588 3551 7600
rect 3495 7566 3551 7588
rect 3585 7588 3589 7600
rect 3623 7600 3689 7622
rect 3623 7588 3641 7600
rect 3585 7566 3641 7588
rect 3675 7588 3689 7600
rect 3723 7600 3789 7622
rect 3823 7600 3889 7622
rect 3923 7600 3989 7622
rect 4023 7600 4096 7622
rect 3723 7588 3731 7600
rect 3675 7566 3731 7588
rect 3765 7588 3789 7600
rect 3855 7588 3889 7600
rect 3945 7588 3989 7600
rect 3765 7566 3821 7588
rect 3855 7566 3911 7588
rect 3945 7566 4001 7588
rect 4035 7566 4096 7600
rect 3402 7522 4096 7566
rect 3402 7510 3489 7522
rect 3523 7510 3589 7522
rect 3402 7476 3461 7510
rect 3523 7488 3551 7510
rect 3495 7476 3551 7488
rect 3585 7488 3589 7510
rect 3623 7510 3689 7522
rect 3623 7488 3641 7510
rect 3585 7476 3641 7488
rect 3675 7488 3689 7510
rect 3723 7510 3789 7522
rect 3823 7510 3889 7522
rect 3923 7510 3989 7522
rect 4023 7510 4096 7522
rect 3723 7488 3731 7510
rect 3675 7476 3731 7488
rect 3765 7488 3789 7510
rect 3855 7488 3889 7510
rect 3945 7488 3989 7510
rect 3765 7476 3821 7488
rect 3855 7476 3911 7488
rect 3945 7476 4001 7488
rect 4035 7476 4096 7510
rect 3402 7415 4096 7476
rect 4158 8098 4177 8132
rect 4211 8098 4230 8132
rect 4158 8042 4230 8098
rect 4158 8008 4177 8042
rect 4211 8008 4230 8042
rect 4158 7952 4230 8008
rect 4158 7918 4177 7952
rect 4211 7918 4230 7952
rect 4158 7862 4230 7918
rect 4158 7828 4177 7862
rect 4211 7828 4230 7862
rect 4158 7772 4230 7828
rect 4158 7738 4177 7772
rect 4211 7738 4230 7772
rect 4158 7682 4230 7738
rect 4158 7648 4177 7682
rect 4211 7648 4230 7682
rect 4158 7592 4230 7648
rect 4158 7558 4177 7592
rect 4211 7558 4230 7592
rect 4158 7502 4230 7558
rect 4158 7468 4177 7502
rect 4211 7468 4230 7502
rect 3268 7353 3340 7412
rect 4158 7412 4230 7468
rect 4158 7378 4177 7412
rect 4211 7378 4230 7412
rect 4158 7353 4230 7378
rect 3340 7334 4158 7353
rect 3340 7300 3344 7334
rect 3378 7300 3434 7334
rect 3468 7300 3524 7334
rect 3558 7300 3614 7334
rect 3648 7300 3704 7334
rect 3738 7300 3794 7334
rect 3828 7300 3884 7334
rect 3918 7300 3974 7334
rect 4008 7300 4064 7334
rect 4098 7300 4158 7334
rect 3340 7281 4158 7300
rect 4294 8238 4327 8272
rect 4361 8238 4393 8272
rect 4294 8182 4393 8238
rect 4294 8148 4327 8182
rect 4361 8148 4393 8182
rect 4294 8092 4393 8148
rect 4294 8058 4327 8092
rect 4361 8058 4393 8092
rect 4294 8002 4393 8058
rect 4294 7968 4327 8002
rect 4361 7968 4393 8002
rect 4294 7912 4393 7968
rect 4294 7878 4327 7912
rect 4361 7878 4393 7912
rect 4294 7822 4393 7878
rect 4294 7788 4327 7822
rect 4361 7788 4393 7822
rect 4294 7732 4393 7788
rect 4294 7698 4327 7732
rect 4361 7698 4393 7732
rect 4294 7642 4393 7698
rect 4294 7608 4327 7642
rect 4361 7608 4393 7642
rect 4294 7552 4393 7608
rect 4294 7518 4327 7552
rect 4361 7518 4393 7552
rect 4294 7462 4393 7518
rect 4294 7428 4327 7462
rect 4361 7428 4393 7462
rect 4294 7372 4393 7428
rect 4294 7353 4327 7372
rect 4361 7353 4393 7372
rect 3105 7248 3140 7281
rect 3174 7248 3204 7281
rect 3105 7217 3204 7248
rect 4294 7248 4327 7281
rect 4361 7248 4393 7281
rect 4294 7217 4393 7248
rect 3105 7186 4393 7217
rect 3105 7152 3163 7186
rect 3197 7152 3253 7186
rect 3287 7152 3343 7186
rect 3377 7152 3433 7186
rect 3467 7152 3523 7186
rect 3557 7152 3613 7186
rect 3647 7152 3703 7186
rect 3737 7152 3793 7186
rect 3827 7152 3883 7186
rect 3917 7152 3973 7186
rect 4007 7152 4063 7186
rect 4097 7152 4153 7186
rect 4187 7152 4243 7186
rect 4277 7152 4393 7186
rect 3105 7118 4393 7152
rect 4493 8373 5781 8406
rect 4493 8339 4551 8373
rect 4585 8339 4641 8373
rect 4675 8339 4731 8373
rect 4765 8339 4821 8373
rect 4855 8339 4911 8373
rect 4945 8339 5001 8373
rect 5035 8339 5091 8373
rect 5125 8339 5181 8373
rect 5215 8339 5271 8373
rect 5305 8339 5361 8373
rect 5395 8339 5451 8373
rect 5485 8339 5541 8373
rect 5575 8339 5631 8373
rect 5665 8339 5781 8373
rect 4493 8307 5781 8339
rect 4493 8272 4592 8307
rect 4493 8238 4528 8272
rect 4562 8238 4592 8272
rect 5682 8272 5781 8307
rect 4493 8182 4592 8238
rect 4493 8148 4528 8182
rect 4562 8148 4592 8182
rect 4493 8092 4592 8148
rect 4493 8058 4528 8092
rect 4562 8058 4592 8092
rect 4493 8002 4592 8058
rect 4493 7968 4528 8002
rect 4562 7968 4592 8002
rect 4493 7912 4592 7968
rect 4493 7878 4528 7912
rect 4562 7878 4592 7912
rect 4493 7822 4592 7878
rect 4493 7788 4528 7822
rect 4562 7788 4592 7822
rect 4493 7732 4592 7788
rect 4493 7698 4528 7732
rect 4562 7698 4592 7732
rect 4493 7642 4592 7698
rect 4493 7608 4528 7642
rect 4562 7608 4592 7642
rect 4493 7552 4592 7608
rect 4493 7518 4528 7552
rect 4562 7518 4592 7552
rect 4493 7462 4592 7518
rect 4493 7428 4528 7462
rect 4562 7428 4592 7462
rect 4493 7372 4592 7428
rect 4493 7353 4528 7372
rect 4562 7353 4592 7372
rect 4656 8224 5618 8243
rect 4656 8190 4751 8224
rect 4785 8190 4841 8224
rect 4875 8190 4931 8224
rect 4965 8190 5021 8224
rect 5055 8190 5111 8224
rect 5145 8190 5201 8224
rect 5235 8190 5291 8224
rect 5325 8190 5381 8224
rect 5415 8190 5471 8224
rect 5505 8190 5618 8224
rect 4656 8171 5618 8190
rect 4656 8166 4728 8171
rect 4656 8132 4675 8166
rect 4709 8132 4728 8166
rect 4656 8076 4728 8132
rect 5546 8132 5618 8171
rect 4656 8042 4675 8076
rect 4709 8042 4728 8076
rect 4656 7986 4728 8042
rect 4656 7952 4675 7986
rect 4709 7952 4728 7986
rect 4656 7896 4728 7952
rect 4656 7862 4675 7896
rect 4709 7862 4728 7896
rect 4656 7806 4728 7862
rect 4656 7772 4675 7806
rect 4709 7772 4728 7806
rect 4656 7716 4728 7772
rect 4656 7682 4675 7716
rect 4709 7682 4728 7716
rect 4656 7626 4728 7682
rect 4656 7592 4675 7626
rect 4709 7592 4728 7626
rect 4656 7536 4728 7592
rect 4656 7502 4675 7536
rect 4709 7502 4728 7536
rect 4656 7446 4728 7502
rect 4656 7412 4675 7446
rect 4709 7412 4728 7446
rect 4790 8050 5484 8109
rect 4790 8016 4849 8050
rect 4883 8022 4939 8050
rect 4911 8016 4939 8022
rect 4973 8022 5029 8050
rect 4973 8016 4977 8022
rect 4790 7988 4877 8016
rect 4911 7988 4977 8016
rect 5011 8016 5029 8022
rect 5063 8022 5119 8050
rect 5063 8016 5077 8022
rect 5011 7988 5077 8016
rect 5111 8016 5119 8022
rect 5153 8022 5209 8050
rect 5243 8022 5299 8050
rect 5333 8022 5389 8050
rect 5153 8016 5177 8022
rect 5243 8016 5277 8022
rect 5333 8016 5377 8022
rect 5423 8016 5484 8050
rect 5111 7988 5177 8016
rect 5211 7988 5277 8016
rect 5311 7988 5377 8016
rect 5411 7988 5484 8016
rect 4790 7960 5484 7988
rect 4790 7926 4849 7960
rect 4883 7926 4939 7960
rect 4973 7926 5029 7960
rect 5063 7926 5119 7960
rect 5153 7926 5209 7960
rect 5243 7926 5299 7960
rect 5333 7926 5389 7960
rect 5423 7926 5484 7960
rect 4790 7922 5484 7926
rect 4790 7888 4877 7922
rect 4911 7888 4977 7922
rect 5011 7888 5077 7922
rect 5111 7888 5177 7922
rect 5211 7888 5277 7922
rect 5311 7888 5377 7922
rect 5411 7888 5484 7922
rect 4790 7870 5484 7888
rect 4790 7836 4849 7870
rect 4883 7836 4939 7870
rect 4973 7836 5029 7870
rect 5063 7836 5119 7870
rect 5153 7836 5209 7870
rect 5243 7836 5299 7870
rect 5333 7836 5389 7870
rect 5423 7836 5484 7870
rect 4790 7822 5484 7836
rect 4790 7788 4877 7822
rect 4911 7788 4977 7822
rect 5011 7788 5077 7822
rect 5111 7788 5177 7822
rect 5211 7788 5277 7822
rect 5311 7788 5377 7822
rect 5411 7788 5484 7822
rect 4790 7780 5484 7788
rect 4790 7746 4849 7780
rect 4883 7746 4939 7780
rect 4973 7746 5029 7780
rect 5063 7746 5119 7780
rect 5153 7746 5209 7780
rect 5243 7746 5299 7780
rect 5333 7746 5389 7780
rect 5423 7746 5484 7780
rect 4790 7722 5484 7746
rect 4790 7690 4877 7722
rect 4911 7690 4977 7722
rect 4790 7656 4849 7690
rect 4911 7688 4939 7690
rect 4883 7656 4939 7688
rect 4973 7688 4977 7690
rect 5011 7690 5077 7722
rect 5011 7688 5029 7690
rect 4973 7656 5029 7688
rect 5063 7688 5077 7690
rect 5111 7690 5177 7722
rect 5211 7690 5277 7722
rect 5311 7690 5377 7722
rect 5411 7690 5484 7722
rect 5111 7688 5119 7690
rect 5063 7656 5119 7688
rect 5153 7688 5177 7690
rect 5243 7688 5277 7690
rect 5333 7688 5377 7690
rect 5153 7656 5209 7688
rect 5243 7656 5299 7688
rect 5333 7656 5389 7688
rect 5423 7656 5484 7690
rect 4790 7622 5484 7656
rect 4790 7600 4877 7622
rect 4911 7600 4977 7622
rect 4790 7566 4849 7600
rect 4911 7588 4939 7600
rect 4883 7566 4939 7588
rect 4973 7588 4977 7600
rect 5011 7600 5077 7622
rect 5011 7588 5029 7600
rect 4973 7566 5029 7588
rect 5063 7588 5077 7600
rect 5111 7600 5177 7622
rect 5211 7600 5277 7622
rect 5311 7600 5377 7622
rect 5411 7600 5484 7622
rect 5111 7588 5119 7600
rect 5063 7566 5119 7588
rect 5153 7588 5177 7600
rect 5243 7588 5277 7600
rect 5333 7588 5377 7600
rect 5153 7566 5209 7588
rect 5243 7566 5299 7588
rect 5333 7566 5389 7588
rect 5423 7566 5484 7600
rect 4790 7522 5484 7566
rect 4790 7510 4877 7522
rect 4911 7510 4977 7522
rect 4790 7476 4849 7510
rect 4911 7488 4939 7510
rect 4883 7476 4939 7488
rect 4973 7488 4977 7510
rect 5011 7510 5077 7522
rect 5011 7488 5029 7510
rect 4973 7476 5029 7488
rect 5063 7488 5077 7510
rect 5111 7510 5177 7522
rect 5211 7510 5277 7522
rect 5311 7510 5377 7522
rect 5411 7510 5484 7522
rect 5111 7488 5119 7510
rect 5063 7476 5119 7488
rect 5153 7488 5177 7510
rect 5243 7488 5277 7510
rect 5333 7488 5377 7510
rect 5153 7476 5209 7488
rect 5243 7476 5299 7488
rect 5333 7476 5389 7488
rect 5423 7476 5484 7510
rect 4790 7415 5484 7476
rect 5546 8098 5565 8132
rect 5599 8098 5618 8132
rect 5546 8042 5618 8098
rect 5546 8008 5565 8042
rect 5599 8008 5618 8042
rect 5546 7952 5618 8008
rect 5546 7918 5565 7952
rect 5599 7918 5618 7952
rect 5546 7862 5618 7918
rect 5546 7828 5565 7862
rect 5599 7828 5618 7862
rect 5546 7772 5618 7828
rect 5546 7738 5565 7772
rect 5599 7738 5618 7772
rect 5546 7682 5618 7738
rect 5546 7648 5565 7682
rect 5599 7648 5618 7682
rect 5546 7592 5618 7648
rect 5546 7558 5565 7592
rect 5599 7558 5618 7592
rect 5546 7502 5618 7558
rect 5546 7468 5565 7502
rect 5599 7468 5618 7502
rect 4656 7353 4728 7412
rect 5546 7412 5618 7468
rect 5546 7378 5565 7412
rect 5599 7378 5618 7412
rect 5546 7353 5618 7378
rect 4728 7334 5546 7353
rect 4728 7300 4732 7334
rect 4766 7300 4822 7334
rect 4856 7300 4912 7334
rect 4946 7300 5002 7334
rect 5036 7300 5092 7334
rect 5126 7300 5182 7334
rect 5216 7300 5272 7334
rect 5306 7300 5362 7334
rect 5396 7300 5452 7334
rect 5486 7300 5546 7334
rect 4728 7281 5546 7300
rect 5682 8238 5715 8272
rect 5749 8238 5781 8272
rect 5682 8182 5781 8238
rect 5682 8148 5715 8182
rect 5749 8148 5781 8182
rect 5682 8092 5781 8148
rect 5682 8058 5715 8092
rect 5749 8058 5781 8092
rect 5682 8002 5781 8058
rect 5682 7968 5715 8002
rect 5749 7968 5781 8002
rect 5682 7912 5781 7968
rect 5682 7878 5715 7912
rect 5749 7878 5781 7912
rect 5682 7822 5781 7878
rect 5682 7788 5715 7822
rect 5749 7788 5781 7822
rect 5682 7732 5781 7788
rect 5682 7698 5715 7732
rect 5749 7698 5781 7732
rect 5682 7642 5781 7698
rect 5682 7608 5715 7642
rect 5749 7608 5781 7642
rect 5682 7552 5781 7608
rect 5682 7518 5715 7552
rect 5749 7518 5781 7552
rect 5682 7462 5781 7518
rect 5682 7428 5715 7462
rect 5749 7428 5781 7462
rect 5682 7372 5781 7428
rect 5682 7353 5715 7372
rect 5749 7353 5781 7372
rect 4493 7248 4528 7281
rect 4562 7248 4592 7281
rect 4493 7217 4592 7248
rect 5682 7248 5715 7281
rect 5749 7248 5781 7281
rect 5682 7217 5781 7248
rect 4493 7186 5781 7217
rect 4493 7152 4551 7186
rect 4585 7152 4641 7186
rect 4675 7152 4731 7186
rect 4765 7152 4821 7186
rect 4855 7152 4911 7186
rect 4945 7152 5001 7186
rect 5035 7152 5091 7186
rect 5125 7152 5181 7186
rect 5215 7152 5271 7186
rect 5305 7152 5361 7186
rect 5395 7152 5451 7186
rect 5485 7152 5541 7186
rect 5575 7152 5631 7186
rect 5665 7152 5781 7186
rect 4493 7118 5781 7152
rect 5881 8373 7169 8406
rect 5881 8339 5939 8373
rect 5973 8339 6029 8373
rect 6063 8339 6119 8373
rect 6153 8339 6209 8373
rect 6243 8339 6299 8373
rect 6333 8339 6389 8373
rect 6423 8339 6479 8373
rect 6513 8339 6569 8373
rect 6603 8339 6659 8373
rect 6693 8339 6749 8373
rect 6783 8339 6839 8373
rect 6873 8339 6929 8373
rect 6963 8339 7019 8373
rect 7053 8339 7169 8373
rect 5881 8307 7169 8339
rect 5881 8272 5980 8307
rect 5881 8238 5916 8272
rect 5950 8238 5980 8272
rect 7070 8272 7169 8307
rect 5881 8182 5980 8238
rect 5881 8148 5916 8182
rect 5950 8148 5980 8182
rect 5881 8092 5980 8148
rect 5881 8058 5916 8092
rect 5950 8058 5980 8092
rect 5881 8002 5980 8058
rect 5881 7968 5916 8002
rect 5950 7968 5980 8002
rect 5881 7912 5980 7968
rect 5881 7878 5916 7912
rect 5950 7878 5980 7912
rect 5881 7822 5980 7878
rect 5881 7788 5916 7822
rect 5950 7788 5980 7822
rect 5881 7732 5980 7788
rect 5881 7698 5916 7732
rect 5950 7698 5980 7732
rect 5881 7642 5980 7698
rect 5881 7608 5916 7642
rect 5950 7608 5980 7642
rect 5881 7552 5980 7608
rect 5881 7518 5916 7552
rect 5950 7518 5980 7552
rect 5881 7462 5980 7518
rect 5881 7428 5916 7462
rect 5950 7428 5980 7462
rect 5881 7372 5980 7428
rect 5881 7353 5916 7372
rect 5950 7353 5980 7372
rect 6044 8224 7006 8243
rect 6044 8190 6139 8224
rect 6173 8190 6229 8224
rect 6263 8190 6319 8224
rect 6353 8190 6409 8224
rect 6443 8190 6499 8224
rect 6533 8190 6589 8224
rect 6623 8190 6679 8224
rect 6713 8190 6769 8224
rect 6803 8190 6859 8224
rect 6893 8190 7006 8224
rect 6044 8171 7006 8190
rect 6044 8166 6116 8171
rect 6044 8132 6063 8166
rect 6097 8132 6116 8166
rect 6044 8076 6116 8132
rect 6934 8132 7006 8171
rect 6044 8042 6063 8076
rect 6097 8042 6116 8076
rect 6044 7986 6116 8042
rect 6044 7952 6063 7986
rect 6097 7952 6116 7986
rect 6044 7896 6116 7952
rect 6044 7862 6063 7896
rect 6097 7862 6116 7896
rect 6044 7806 6116 7862
rect 6044 7772 6063 7806
rect 6097 7772 6116 7806
rect 6044 7716 6116 7772
rect 6044 7682 6063 7716
rect 6097 7682 6116 7716
rect 6044 7626 6116 7682
rect 6044 7592 6063 7626
rect 6097 7592 6116 7626
rect 6044 7536 6116 7592
rect 6044 7502 6063 7536
rect 6097 7502 6116 7536
rect 6044 7446 6116 7502
rect 6044 7412 6063 7446
rect 6097 7412 6116 7446
rect 6178 8050 6872 8109
rect 6178 8016 6237 8050
rect 6271 8022 6327 8050
rect 6299 8016 6327 8022
rect 6361 8022 6417 8050
rect 6361 8016 6365 8022
rect 6178 7988 6265 8016
rect 6299 7988 6365 8016
rect 6399 8016 6417 8022
rect 6451 8022 6507 8050
rect 6451 8016 6465 8022
rect 6399 7988 6465 8016
rect 6499 8016 6507 8022
rect 6541 8022 6597 8050
rect 6631 8022 6687 8050
rect 6721 8022 6777 8050
rect 6541 8016 6565 8022
rect 6631 8016 6665 8022
rect 6721 8016 6765 8022
rect 6811 8016 6872 8050
rect 6499 7988 6565 8016
rect 6599 7988 6665 8016
rect 6699 7988 6765 8016
rect 6799 7988 6872 8016
rect 6178 7960 6872 7988
rect 6178 7926 6237 7960
rect 6271 7926 6327 7960
rect 6361 7926 6417 7960
rect 6451 7926 6507 7960
rect 6541 7926 6597 7960
rect 6631 7926 6687 7960
rect 6721 7926 6777 7960
rect 6811 7926 6872 7960
rect 6178 7922 6872 7926
rect 6178 7888 6265 7922
rect 6299 7888 6365 7922
rect 6399 7888 6465 7922
rect 6499 7888 6565 7922
rect 6599 7888 6665 7922
rect 6699 7888 6765 7922
rect 6799 7888 6872 7922
rect 6178 7870 6872 7888
rect 6178 7836 6237 7870
rect 6271 7836 6327 7870
rect 6361 7836 6417 7870
rect 6451 7836 6507 7870
rect 6541 7836 6597 7870
rect 6631 7836 6687 7870
rect 6721 7836 6777 7870
rect 6811 7836 6872 7870
rect 6178 7822 6872 7836
rect 6178 7788 6265 7822
rect 6299 7788 6365 7822
rect 6399 7788 6465 7822
rect 6499 7788 6565 7822
rect 6599 7788 6665 7822
rect 6699 7788 6765 7822
rect 6799 7788 6872 7822
rect 6178 7780 6872 7788
rect 6178 7746 6237 7780
rect 6271 7746 6327 7780
rect 6361 7746 6417 7780
rect 6451 7746 6507 7780
rect 6541 7746 6597 7780
rect 6631 7746 6687 7780
rect 6721 7746 6777 7780
rect 6811 7746 6872 7780
rect 6178 7722 6872 7746
rect 6178 7690 6265 7722
rect 6299 7690 6365 7722
rect 6178 7656 6237 7690
rect 6299 7688 6327 7690
rect 6271 7656 6327 7688
rect 6361 7688 6365 7690
rect 6399 7690 6465 7722
rect 6399 7688 6417 7690
rect 6361 7656 6417 7688
rect 6451 7688 6465 7690
rect 6499 7690 6565 7722
rect 6599 7690 6665 7722
rect 6699 7690 6765 7722
rect 6799 7690 6872 7722
rect 6499 7688 6507 7690
rect 6451 7656 6507 7688
rect 6541 7688 6565 7690
rect 6631 7688 6665 7690
rect 6721 7688 6765 7690
rect 6541 7656 6597 7688
rect 6631 7656 6687 7688
rect 6721 7656 6777 7688
rect 6811 7656 6872 7690
rect 6178 7622 6872 7656
rect 6178 7600 6265 7622
rect 6299 7600 6365 7622
rect 6178 7566 6237 7600
rect 6299 7588 6327 7600
rect 6271 7566 6327 7588
rect 6361 7588 6365 7600
rect 6399 7600 6465 7622
rect 6399 7588 6417 7600
rect 6361 7566 6417 7588
rect 6451 7588 6465 7600
rect 6499 7600 6565 7622
rect 6599 7600 6665 7622
rect 6699 7600 6765 7622
rect 6799 7600 6872 7622
rect 6499 7588 6507 7600
rect 6451 7566 6507 7588
rect 6541 7588 6565 7600
rect 6631 7588 6665 7600
rect 6721 7588 6765 7600
rect 6541 7566 6597 7588
rect 6631 7566 6687 7588
rect 6721 7566 6777 7588
rect 6811 7566 6872 7600
rect 6178 7522 6872 7566
rect 6178 7510 6265 7522
rect 6299 7510 6365 7522
rect 6178 7476 6237 7510
rect 6299 7488 6327 7510
rect 6271 7476 6327 7488
rect 6361 7488 6365 7510
rect 6399 7510 6465 7522
rect 6399 7488 6417 7510
rect 6361 7476 6417 7488
rect 6451 7488 6465 7510
rect 6499 7510 6565 7522
rect 6599 7510 6665 7522
rect 6699 7510 6765 7522
rect 6799 7510 6872 7522
rect 6499 7488 6507 7510
rect 6451 7476 6507 7488
rect 6541 7488 6565 7510
rect 6631 7488 6665 7510
rect 6721 7488 6765 7510
rect 6541 7476 6597 7488
rect 6631 7476 6687 7488
rect 6721 7476 6777 7488
rect 6811 7476 6872 7510
rect 6178 7415 6872 7476
rect 6934 8098 6953 8132
rect 6987 8098 7006 8132
rect 6934 8042 7006 8098
rect 6934 8008 6953 8042
rect 6987 8008 7006 8042
rect 6934 7952 7006 8008
rect 6934 7918 6953 7952
rect 6987 7918 7006 7952
rect 6934 7862 7006 7918
rect 6934 7828 6953 7862
rect 6987 7828 7006 7862
rect 6934 7772 7006 7828
rect 6934 7738 6953 7772
rect 6987 7738 7006 7772
rect 6934 7682 7006 7738
rect 6934 7648 6953 7682
rect 6987 7648 7006 7682
rect 6934 7592 7006 7648
rect 6934 7558 6953 7592
rect 6987 7558 7006 7592
rect 6934 7502 7006 7558
rect 6934 7468 6953 7502
rect 6987 7468 7006 7502
rect 6044 7353 6116 7412
rect 6934 7412 7006 7468
rect 6934 7378 6953 7412
rect 6987 7378 7006 7412
rect 6934 7353 7006 7378
rect 6116 7334 7006 7353
rect 6116 7300 6120 7334
rect 6154 7300 6210 7334
rect 6244 7300 6300 7334
rect 6334 7300 6390 7334
rect 6424 7300 6480 7334
rect 6514 7300 6570 7334
rect 6604 7300 6660 7334
rect 6694 7300 6750 7334
rect 6784 7300 6840 7334
rect 6874 7300 7006 7334
rect 6116 7281 7006 7300
rect 7070 8238 7103 8272
rect 7137 8238 7169 8272
rect 7070 8182 7169 8238
rect 7070 8148 7103 8182
rect 7137 8148 7169 8182
rect 7070 8092 7169 8148
rect 7070 8058 7103 8092
rect 7137 8058 7169 8092
rect 7070 8002 7169 8058
rect 7070 7968 7103 8002
rect 7137 7968 7169 8002
rect 7070 7912 7169 7968
rect 7070 7878 7103 7912
rect 7137 7878 7169 7912
rect 7070 7822 7169 7878
rect 7070 7788 7103 7822
rect 7137 7788 7169 7822
rect 7070 7732 7169 7788
rect 7070 7698 7103 7732
rect 7137 7698 7169 7732
rect 7070 7642 7169 7698
rect 7070 7608 7103 7642
rect 7137 7608 7169 7642
rect 7070 7552 7169 7608
rect 7070 7518 7103 7552
rect 7137 7518 7169 7552
rect 7070 7462 7169 7518
rect 7070 7428 7103 7462
rect 7137 7428 7169 7462
rect 7070 7372 7169 7428
rect 7070 7338 7103 7372
rect 7137 7338 7169 7372
rect 7070 7282 7169 7338
rect 5881 7248 5916 7281
rect 5950 7248 5980 7281
rect 5881 7217 5980 7248
rect 7070 7248 7103 7282
rect 7137 7248 7169 7282
rect 7070 7217 7169 7248
rect 5881 7186 6044 7217
rect 6116 7186 7169 7217
rect 5881 7152 5939 7186
rect 5973 7152 6029 7186
rect 6116 7152 6119 7186
rect 6153 7152 6209 7186
rect 6243 7152 6299 7186
rect 6333 7152 6389 7186
rect 6423 7152 6479 7186
rect 6513 7152 6569 7186
rect 6603 7152 6659 7186
rect 6693 7152 6749 7186
rect 6783 7152 6839 7186
rect 6873 7152 6929 7186
rect 6963 7152 7019 7186
rect 7053 7152 7169 7186
rect 5881 7118 6044 7152
rect 6116 7118 7169 7152
rect 329 6985 1382 7018
rect 1454 6985 1617 7018
rect 329 6951 387 6985
rect 421 6951 477 6985
rect 511 6951 567 6985
rect 601 6951 657 6985
rect 691 6951 747 6985
rect 781 6951 837 6985
rect 871 6951 927 6985
rect 961 6951 1017 6985
rect 1051 6951 1107 6985
rect 1141 6951 1197 6985
rect 1231 6951 1287 6985
rect 1321 6951 1377 6985
rect 1454 6951 1467 6985
rect 1501 6951 1617 6985
rect 329 6919 1382 6951
rect 1454 6919 1617 6951
rect 329 6884 428 6919
rect 329 6850 364 6884
rect 398 6850 428 6884
rect 1518 6884 1617 6919
rect 329 6794 428 6850
rect 329 6760 364 6794
rect 398 6760 428 6794
rect 329 6704 428 6760
rect 329 6670 364 6704
rect 398 6670 428 6704
rect 329 6614 428 6670
rect 329 6580 364 6614
rect 398 6580 428 6614
rect 329 6524 428 6580
rect 329 6490 364 6524
rect 398 6490 428 6524
rect 329 6434 428 6490
rect 329 6400 364 6434
rect 398 6400 428 6434
rect 329 6344 428 6400
rect 329 6310 364 6344
rect 398 6310 428 6344
rect 329 6254 428 6310
rect 329 6220 364 6254
rect 398 6220 428 6254
rect 329 6164 428 6220
rect 329 6130 364 6164
rect 398 6130 428 6164
rect 329 6074 428 6130
rect 329 6040 364 6074
rect 398 6040 428 6074
rect 329 5984 428 6040
rect 329 5950 364 5984
rect 398 5950 428 5984
rect 329 5894 428 5950
rect 329 5860 364 5894
rect 398 5860 428 5894
rect 492 6836 1382 6855
rect 492 6802 587 6836
rect 621 6802 677 6836
rect 711 6802 767 6836
rect 801 6802 857 6836
rect 891 6802 947 6836
rect 981 6802 1037 6836
rect 1071 6802 1127 6836
rect 1161 6802 1217 6836
rect 1251 6802 1307 6836
rect 1341 6802 1382 6836
rect 492 6783 1382 6802
rect 492 6778 564 6783
rect 492 6744 511 6778
rect 545 6744 564 6778
rect 492 6688 564 6744
rect 1382 6744 1454 6783
rect 492 6654 511 6688
rect 545 6654 564 6688
rect 492 6598 564 6654
rect 492 6564 511 6598
rect 545 6564 564 6598
rect 492 6508 564 6564
rect 492 6474 511 6508
rect 545 6474 564 6508
rect 492 6418 564 6474
rect 492 6384 511 6418
rect 545 6384 564 6418
rect 492 6328 564 6384
rect 492 6294 511 6328
rect 545 6294 564 6328
rect 492 6238 564 6294
rect 492 6204 511 6238
rect 545 6204 564 6238
rect 492 6148 564 6204
rect 492 6114 511 6148
rect 545 6114 564 6148
rect 492 6058 564 6114
rect 492 6024 511 6058
rect 545 6024 564 6058
rect 626 6662 1320 6721
rect 626 6628 685 6662
rect 719 6634 775 6662
rect 747 6628 775 6634
rect 809 6634 865 6662
rect 809 6628 813 6634
rect 626 6600 713 6628
rect 747 6600 813 6628
rect 847 6628 865 6634
rect 899 6634 955 6662
rect 899 6628 913 6634
rect 847 6600 913 6628
rect 947 6628 955 6634
rect 989 6634 1045 6662
rect 1079 6634 1135 6662
rect 1169 6634 1225 6662
rect 989 6628 1013 6634
rect 1079 6628 1113 6634
rect 1169 6628 1213 6634
rect 1259 6628 1320 6662
rect 947 6600 1013 6628
rect 1047 6600 1113 6628
rect 1147 6600 1213 6628
rect 1247 6600 1320 6628
rect 626 6572 1320 6600
rect 626 6538 685 6572
rect 719 6538 775 6572
rect 809 6538 865 6572
rect 899 6538 955 6572
rect 989 6538 1045 6572
rect 1079 6538 1135 6572
rect 1169 6538 1225 6572
rect 1259 6538 1320 6572
rect 626 6534 1320 6538
rect 626 6500 713 6534
rect 747 6500 813 6534
rect 847 6500 913 6534
rect 947 6500 1013 6534
rect 1047 6500 1113 6534
rect 1147 6500 1213 6534
rect 1247 6500 1320 6534
rect 626 6482 1320 6500
rect 626 6448 685 6482
rect 719 6448 775 6482
rect 809 6448 865 6482
rect 899 6448 955 6482
rect 989 6448 1045 6482
rect 1079 6448 1135 6482
rect 1169 6448 1225 6482
rect 1259 6448 1320 6482
rect 626 6434 1320 6448
rect 626 6400 713 6434
rect 747 6400 813 6434
rect 847 6400 913 6434
rect 947 6400 1013 6434
rect 1047 6400 1113 6434
rect 1147 6400 1213 6434
rect 1247 6400 1320 6434
rect 626 6392 1320 6400
rect 626 6358 685 6392
rect 719 6358 775 6392
rect 809 6358 865 6392
rect 899 6358 955 6392
rect 989 6358 1045 6392
rect 1079 6358 1135 6392
rect 1169 6358 1225 6392
rect 1259 6358 1320 6392
rect 626 6334 1320 6358
rect 626 6302 713 6334
rect 747 6302 813 6334
rect 626 6268 685 6302
rect 747 6300 775 6302
rect 719 6268 775 6300
rect 809 6300 813 6302
rect 847 6302 913 6334
rect 847 6300 865 6302
rect 809 6268 865 6300
rect 899 6300 913 6302
rect 947 6302 1013 6334
rect 1047 6302 1113 6334
rect 1147 6302 1213 6334
rect 1247 6302 1320 6334
rect 947 6300 955 6302
rect 899 6268 955 6300
rect 989 6300 1013 6302
rect 1079 6300 1113 6302
rect 1169 6300 1213 6302
rect 989 6268 1045 6300
rect 1079 6268 1135 6300
rect 1169 6268 1225 6300
rect 1259 6268 1320 6302
rect 626 6234 1320 6268
rect 626 6212 713 6234
rect 747 6212 813 6234
rect 626 6178 685 6212
rect 747 6200 775 6212
rect 719 6178 775 6200
rect 809 6200 813 6212
rect 847 6212 913 6234
rect 847 6200 865 6212
rect 809 6178 865 6200
rect 899 6200 913 6212
rect 947 6212 1013 6234
rect 1047 6212 1113 6234
rect 1147 6212 1213 6234
rect 1247 6212 1320 6234
rect 947 6200 955 6212
rect 899 6178 955 6200
rect 989 6200 1013 6212
rect 1079 6200 1113 6212
rect 1169 6200 1213 6212
rect 989 6178 1045 6200
rect 1079 6178 1135 6200
rect 1169 6178 1225 6200
rect 1259 6178 1320 6212
rect 626 6134 1320 6178
rect 626 6122 713 6134
rect 747 6122 813 6134
rect 626 6088 685 6122
rect 747 6100 775 6122
rect 719 6088 775 6100
rect 809 6100 813 6122
rect 847 6122 913 6134
rect 847 6100 865 6122
rect 809 6088 865 6100
rect 899 6100 913 6122
rect 947 6122 1013 6134
rect 1047 6122 1113 6134
rect 1147 6122 1213 6134
rect 1247 6122 1320 6134
rect 947 6100 955 6122
rect 899 6088 955 6100
rect 989 6100 1013 6122
rect 1079 6100 1113 6122
rect 1169 6100 1213 6122
rect 989 6088 1045 6100
rect 1079 6088 1135 6100
rect 1169 6088 1225 6100
rect 1259 6088 1320 6122
rect 626 6027 1320 6088
rect 1382 6710 1401 6744
rect 1435 6710 1454 6744
rect 1382 6654 1454 6710
rect 1382 6620 1401 6654
rect 1435 6620 1454 6654
rect 1382 6564 1454 6620
rect 1382 6530 1401 6564
rect 1435 6530 1454 6564
rect 1382 6474 1454 6530
rect 1382 6440 1401 6474
rect 1435 6440 1454 6474
rect 1382 6384 1454 6440
rect 1382 6350 1401 6384
rect 1435 6350 1454 6384
rect 1382 6294 1454 6350
rect 1382 6260 1401 6294
rect 1435 6260 1454 6294
rect 1382 6204 1454 6260
rect 1382 6170 1401 6204
rect 1435 6170 1454 6204
rect 1382 6114 1454 6170
rect 1382 6080 1401 6114
rect 1435 6080 1454 6114
rect 492 5965 564 6024
rect 1382 6024 1454 6080
rect 1382 5990 1401 6024
rect 1435 5990 1454 6024
rect 1382 5965 1454 5990
rect 492 5946 1382 5965
rect 492 5912 568 5946
rect 602 5912 658 5946
rect 692 5912 748 5946
rect 782 5912 838 5946
rect 872 5912 928 5946
rect 962 5912 1018 5946
rect 1052 5912 1108 5946
rect 1142 5912 1198 5946
rect 1232 5912 1288 5946
rect 1322 5912 1382 5946
rect 492 5893 1382 5912
rect 1518 6850 1551 6884
rect 1585 6850 1617 6884
rect 1518 6794 1617 6850
rect 1518 6760 1551 6794
rect 1585 6760 1617 6794
rect 1518 6704 1617 6760
rect 1518 6670 1551 6704
rect 1585 6670 1617 6704
rect 1518 6614 1617 6670
rect 1518 6580 1551 6614
rect 1585 6580 1617 6614
rect 1518 6524 1617 6580
rect 1518 6490 1551 6524
rect 1585 6490 1617 6524
rect 1518 6434 1617 6490
rect 1518 6400 1551 6434
rect 1585 6400 1617 6434
rect 1518 6344 1617 6400
rect 1518 6310 1551 6344
rect 1585 6310 1617 6344
rect 1518 6254 1617 6310
rect 1518 6220 1551 6254
rect 1585 6220 1617 6254
rect 1518 6164 1617 6220
rect 1518 6130 1551 6164
rect 1585 6130 1617 6164
rect 1518 6074 1617 6130
rect 1518 6040 1551 6074
rect 1585 6040 1617 6074
rect 1518 5984 1617 6040
rect 1518 5950 1551 5984
rect 1585 5950 1617 5984
rect 1518 5894 1617 5950
rect 329 5829 428 5860
rect 1518 5860 1551 5894
rect 1585 5860 1617 5894
rect 1518 5829 1617 5860
rect 329 5798 1382 5829
rect 1454 5798 1617 5829
rect 329 5764 387 5798
rect 421 5764 477 5798
rect 511 5764 567 5798
rect 601 5764 657 5798
rect 691 5764 747 5798
rect 781 5764 837 5798
rect 871 5764 927 5798
rect 961 5764 1017 5798
rect 1051 5764 1107 5798
rect 1141 5764 1197 5798
rect 1231 5764 1287 5798
rect 1321 5764 1377 5798
rect 1454 5764 1467 5798
rect 1501 5764 1617 5798
rect 329 5730 1382 5764
rect 1454 5730 1617 5764
rect 1717 6985 3005 7018
rect 1717 6951 1775 6985
rect 1809 6951 1865 6985
rect 1899 6951 1955 6985
rect 1989 6951 2045 6985
rect 2079 6951 2135 6985
rect 2169 6951 2225 6985
rect 2259 6951 2315 6985
rect 2349 6951 2405 6985
rect 2439 6951 2495 6985
rect 2529 6951 2585 6985
rect 2619 6951 2675 6985
rect 2709 6951 2765 6985
rect 2799 6951 2855 6985
rect 2889 6951 3005 6985
rect 1717 6919 3005 6951
rect 1717 6884 1816 6919
rect 1717 6850 1752 6884
rect 1786 6850 1816 6884
rect 2906 6884 3005 6919
rect 1717 6794 1816 6850
rect 1717 6760 1752 6794
rect 1786 6760 1816 6794
rect 1717 6704 1816 6760
rect 1717 6670 1752 6704
rect 1786 6670 1816 6704
rect 1717 6614 1816 6670
rect 1717 6580 1752 6614
rect 1786 6580 1816 6614
rect 1717 6524 1816 6580
rect 1717 6490 1752 6524
rect 1786 6490 1816 6524
rect 1717 6434 1816 6490
rect 1717 6400 1752 6434
rect 1786 6400 1816 6434
rect 1717 6344 1816 6400
rect 1717 6310 1752 6344
rect 1786 6310 1816 6344
rect 1717 6254 1816 6310
rect 1717 6220 1752 6254
rect 1786 6220 1816 6254
rect 1717 6164 1816 6220
rect 1717 6130 1752 6164
rect 1786 6130 1816 6164
rect 1717 6074 1816 6130
rect 1717 6040 1752 6074
rect 1786 6040 1816 6074
rect 1717 5984 1816 6040
rect 1717 5950 1752 5984
rect 1786 5950 1816 5984
rect 1717 5894 1816 5950
rect 1717 5860 1752 5894
rect 1786 5860 1816 5894
rect 1880 6836 2842 6855
rect 1880 6802 1975 6836
rect 2009 6802 2065 6836
rect 2099 6802 2155 6836
rect 2189 6802 2245 6836
rect 2279 6802 2335 6836
rect 2369 6802 2425 6836
rect 2459 6802 2515 6836
rect 2549 6802 2605 6836
rect 2639 6802 2695 6836
rect 2729 6802 2842 6836
rect 1880 6783 2842 6802
rect 1880 6778 1952 6783
rect 1880 6744 1899 6778
rect 1933 6744 1952 6778
rect 1880 6688 1952 6744
rect 2770 6744 2842 6783
rect 1880 6654 1899 6688
rect 1933 6654 1952 6688
rect 1880 6598 1952 6654
rect 1880 6564 1899 6598
rect 1933 6564 1952 6598
rect 1880 6508 1952 6564
rect 1880 6474 1899 6508
rect 1933 6474 1952 6508
rect 1880 6418 1952 6474
rect 1880 6384 1899 6418
rect 1933 6384 1952 6418
rect 1880 6328 1952 6384
rect 1880 6294 1899 6328
rect 1933 6294 1952 6328
rect 1880 6238 1952 6294
rect 1880 6204 1899 6238
rect 1933 6204 1952 6238
rect 1880 6148 1952 6204
rect 1880 6114 1899 6148
rect 1933 6114 1952 6148
rect 1880 6058 1952 6114
rect 1880 6024 1899 6058
rect 1933 6024 1952 6058
rect 2014 6662 2708 6721
rect 2014 6628 2073 6662
rect 2107 6634 2163 6662
rect 2135 6628 2163 6634
rect 2197 6634 2253 6662
rect 2197 6628 2201 6634
rect 2014 6600 2101 6628
rect 2135 6600 2201 6628
rect 2235 6628 2253 6634
rect 2287 6634 2343 6662
rect 2287 6628 2301 6634
rect 2235 6600 2301 6628
rect 2335 6628 2343 6634
rect 2377 6634 2433 6662
rect 2467 6634 2523 6662
rect 2557 6634 2613 6662
rect 2377 6628 2401 6634
rect 2467 6628 2501 6634
rect 2557 6628 2601 6634
rect 2647 6628 2708 6662
rect 2335 6600 2401 6628
rect 2435 6600 2501 6628
rect 2535 6600 2601 6628
rect 2635 6600 2708 6628
rect 2014 6572 2708 6600
rect 2014 6538 2073 6572
rect 2107 6538 2163 6572
rect 2197 6538 2253 6572
rect 2287 6538 2343 6572
rect 2377 6538 2433 6572
rect 2467 6538 2523 6572
rect 2557 6538 2613 6572
rect 2647 6538 2708 6572
rect 2014 6534 2708 6538
rect 2014 6500 2101 6534
rect 2135 6500 2201 6534
rect 2235 6500 2301 6534
rect 2335 6500 2401 6534
rect 2435 6500 2501 6534
rect 2535 6500 2601 6534
rect 2635 6500 2708 6534
rect 2014 6482 2708 6500
rect 2014 6448 2073 6482
rect 2107 6448 2163 6482
rect 2197 6448 2253 6482
rect 2287 6448 2343 6482
rect 2377 6448 2433 6482
rect 2467 6448 2523 6482
rect 2557 6448 2613 6482
rect 2647 6448 2708 6482
rect 2014 6434 2708 6448
rect 2014 6400 2101 6434
rect 2135 6400 2201 6434
rect 2235 6400 2301 6434
rect 2335 6400 2401 6434
rect 2435 6400 2501 6434
rect 2535 6400 2601 6434
rect 2635 6400 2708 6434
rect 2014 6392 2708 6400
rect 2014 6358 2073 6392
rect 2107 6358 2163 6392
rect 2197 6358 2253 6392
rect 2287 6358 2343 6392
rect 2377 6358 2433 6392
rect 2467 6358 2523 6392
rect 2557 6358 2613 6392
rect 2647 6358 2708 6392
rect 2014 6334 2708 6358
rect 2014 6302 2101 6334
rect 2135 6302 2201 6334
rect 2014 6268 2073 6302
rect 2135 6300 2163 6302
rect 2107 6268 2163 6300
rect 2197 6300 2201 6302
rect 2235 6302 2301 6334
rect 2235 6300 2253 6302
rect 2197 6268 2253 6300
rect 2287 6300 2301 6302
rect 2335 6302 2401 6334
rect 2435 6302 2501 6334
rect 2535 6302 2601 6334
rect 2635 6302 2708 6334
rect 2335 6300 2343 6302
rect 2287 6268 2343 6300
rect 2377 6300 2401 6302
rect 2467 6300 2501 6302
rect 2557 6300 2601 6302
rect 2377 6268 2433 6300
rect 2467 6268 2523 6300
rect 2557 6268 2613 6300
rect 2647 6268 2708 6302
rect 2014 6234 2708 6268
rect 2014 6212 2101 6234
rect 2135 6212 2201 6234
rect 2014 6178 2073 6212
rect 2135 6200 2163 6212
rect 2107 6178 2163 6200
rect 2197 6200 2201 6212
rect 2235 6212 2301 6234
rect 2235 6200 2253 6212
rect 2197 6178 2253 6200
rect 2287 6200 2301 6212
rect 2335 6212 2401 6234
rect 2435 6212 2501 6234
rect 2535 6212 2601 6234
rect 2635 6212 2708 6234
rect 2335 6200 2343 6212
rect 2287 6178 2343 6200
rect 2377 6200 2401 6212
rect 2467 6200 2501 6212
rect 2557 6200 2601 6212
rect 2377 6178 2433 6200
rect 2467 6178 2523 6200
rect 2557 6178 2613 6200
rect 2647 6178 2708 6212
rect 2014 6134 2708 6178
rect 2014 6122 2101 6134
rect 2135 6122 2201 6134
rect 2014 6088 2073 6122
rect 2135 6100 2163 6122
rect 2107 6088 2163 6100
rect 2197 6100 2201 6122
rect 2235 6122 2301 6134
rect 2235 6100 2253 6122
rect 2197 6088 2253 6100
rect 2287 6100 2301 6122
rect 2335 6122 2401 6134
rect 2435 6122 2501 6134
rect 2535 6122 2601 6134
rect 2635 6122 2708 6134
rect 2335 6100 2343 6122
rect 2287 6088 2343 6100
rect 2377 6100 2401 6122
rect 2467 6100 2501 6122
rect 2557 6100 2601 6122
rect 2377 6088 2433 6100
rect 2467 6088 2523 6100
rect 2557 6088 2613 6100
rect 2647 6088 2708 6122
rect 2014 6027 2708 6088
rect 2770 6710 2789 6744
rect 2823 6710 2842 6744
rect 2770 6654 2842 6710
rect 2770 6620 2789 6654
rect 2823 6620 2842 6654
rect 2770 6564 2842 6620
rect 2770 6530 2789 6564
rect 2823 6530 2842 6564
rect 2770 6474 2842 6530
rect 2770 6440 2789 6474
rect 2823 6440 2842 6474
rect 2770 6384 2842 6440
rect 2770 6350 2789 6384
rect 2823 6350 2842 6384
rect 2770 6294 2842 6350
rect 2770 6260 2789 6294
rect 2823 6260 2842 6294
rect 2770 6204 2842 6260
rect 2770 6170 2789 6204
rect 2823 6170 2842 6204
rect 2770 6114 2842 6170
rect 2770 6080 2789 6114
rect 2823 6080 2842 6114
rect 1880 5965 1952 6024
rect 2770 6024 2842 6080
rect 2770 5990 2789 6024
rect 2823 5990 2842 6024
rect 2770 5965 2842 5990
rect 1880 5946 2770 5965
rect 1880 5912 1956 5946
rect 1990 5912 2046 5946
rect 2080 5912 2136 5946
rect 2170 5912 2226 5946
rect 2260 5912 2316 5946
rect 2350 5912 2406 5946
rect 2440 5912 2496 5946
rect 2530 5912 2586 5946
rect 2620 5912 2676 5946
rect 2710 5912 2770 5946
rect 1880 5893 2770 5912
rect 2906 6850 2939 6884
rect 2973 6850 3005 6884
rect 2906 6794 3005 6850
rect 2906 6760 2939 6794
rect 2973 6760 3005 6794
rect 2906 6704 3005 6760
rect 2906 6670 2939 6704
rect 2973 6670 3005 6704
rect 2906 6614 3005 6670
rect 2906 6580 2939 6614
rect 2973 6580 3005 6614
rect 2906 6524 3005 6580
rect 2906 6490 2939 6524
rect 2973 6490 3005 6524
rect 2906 6434 3005 6490
rect 2906 6400 2939 6434
rect 2973 6400 3005 6434
rect 2906 6344 3005 6400
rect 2906 6310 2939 6344
rect 2973 6310 3005 6344
rect 2906 6254 3005 6310
rect 2906 6220 2939 6254
rect 2973 6220 3005 6254
rect 2906 6164 3005 6220
rect 2906 6130 2939 6164
rect 2973 6130 3005 6164
rect 2906 6074 3005 6130
rect 2906 6040 2939 6074
rect 2973 6040 3005 6074
rect 2906 5984 3005 6040
rect 2906 5965 2939 5984
rect 2973 5965 3005 5984
rect 1717 5829 1816 5860
rect 2906 5860 2939 5893
rect 2973 5860 3005 5893
rect 2906 5829 3005 5860
rect 1717 5798 2770 5829
rect 2842 5798 3005 5829
rect 1717 5764 1775 5798
rect 1809 5764 1865 5798
rect 1899 5764 1955 5798
rect 1989 5764 2045 5798
rect 2079 5764 2135 5798
rect 2169 5764 2225 5798
rect 2259 5764 2315 5798
rect 2349 5764 2405 5798
rect 2439 5764 2495 5798
rect 2529 5764 2585 5798
rect 2619 5764 2675 5798
rect 2709 5764 2765 5798
rect 2842 5764 2855 5798
rect 2889 5764 3005 5798
rect 1717 5730 2770 5764
rect 2842 5730 3005 5764
rect 3105 6985 4393 7018
rect 3105 6951 3163 6985
rect 3197 6951 3253 6985
rect 3287 6951 3343 6985
rect 3377 6951 3433 6985
rect 3467 6951 3523 6985
rect 3557 6951 3613 6985
rect 3647 6951 3703 6985
rect 3737 6951 3793 6985
rect 3827 6951 3883 6985
rect 3917 6951 3973 6985
rect 4007 6951 4063 6985
rect 4097 6951 4153 6985
rect 4187 6951 4243 6985
rect 4277 6951 4393 6985
rect 3105 6919 4393 6951
rect 3105 6884 3204 6919
rect 3105 6850 3140 6884
rect 3174 6850 3204 6884
rect 4294 6884 4393 6919
rect 3105 6794 3204 6850
rect 3105 6760 3140 6794
rect 3174 6760 3204 6794
rect 3105 6704 3204 6760
rect 3105 6670 3140 6704
rect 3174 6670 3204 6704
rect 3105 6614 3204 6670
rect 3105 6580 3140 6614
rect 3174 6580 3204 6614
rect 3105 6524 3204 6580
rect 3105 6490 3140 6524
rect 3174 6490 3204 6524
rect 3105 6434 3204 6490
rect 3105 6400 3140 6434
rect 3174 6400 3204 6434
rect 3105 6344 3204 6400
rect 3105 6310 3140 6344
rect 3174 6310 3204 6344
rect 3105 6254 3204 6310
rect 3105 6220 3140 6254
rect 3174 6220 3204 6254
rect 3105 6164 3204 6220
rect 3105 6130 3140 6164
rect 3174 6130 3204 6164
rect 3105 6074 3204 6130
rect 3105 6040 3140 6074
rect 3174 6040 3204 6074
rect 3105 5984 3204 6040
rect 3105 5965 3140 5984
rect 3174 5965 3204 5984
rect 3268 6836 4230 6855
rect 3268 6802 3363 6836
rect 3397 6802 3453 6836
rect 3487 6802 3543 6836
rect 3577 6802 3633 6836
rect 3667 6802 3723 6836
rect 3757 6802 3813 6836
rect 3847 6802 3903 6836
rect 3937 6802 3993 6836
rect 4027 6802 4083 6836
rect 4117 6802 4230 6836
rect 3268 6783 4230 6802
rect 3268 6778 3340 6783
rect 3268 6744 3287 6778
rect 3321 6744 3340 6778
rect 3268 6688 3340 6744
rect 4158 6744 4230 6783
rect 3268 6654 3287 6688
rect 3321 6654 3340 6688
rect 3268 6598 3340 6654
rect 3268 6564 3287 6598
rect 3321 6564 3340 6598
rect 3268 6508 3340 6564
rect 3268 6474 3287 6508
rect 3321 6474 3340 6508
rect 3268 6418 3340 6474
rect 3268 6384 3287 6418
rect 3321 6384 3340 6418
rect 3268 6328 3340 6384
rect 3268 6294 3287 6328
rect 3321 6294 3340 6328
rect 3268 6238 3340 6294
rect 3268 6204 3287 6238
rect 3321 6204 3340 6238
rect 3268 6148 3340 6204
rect 3268 6114 3287 6148
rect 3321 6114 3340 6148
rect 3268 6058 3340 6114
rect 3268 6024 3287 6058
rect 3321 6024 3340 6058
rect 3402 6662 4096 6721
rect 3402 6628 3461 6662
rect 3495 6634 3551 6662
rect 3523 6628 3551 6634
rect 3585 6634 3641 6662
rect 3585 6628 3589 6634
rect 3402 6600 3489 6628
rect 3523 6600 3589 6628
rect 3623 6628 3641 6634
rect 3675 6634 3731 6662
rect 3675 6628 3689 6634
rect 3623 6600 3689 6628
rect 3723 6628 3731 6634
rect 3765 6634 3821 6662
rect 3855 6634 3911 6662
rect 3945 6634 4001 6662
rect 3765 6628 3789 6634
rect 3855 6628 3889 6634
rect 3945 6628 3989 6634
rect 4035 6628 4096 6662
rect 3723 6600 3789 6628
rect 3823 6600 3889 6628
rect 3923 6600 3989 6628
rect 4023 6600 4096 6628
rect 3402 6572 4096 6600
rect 3402 6538 3461 6572
rect 3495 6538 3551 6572
rect 3585 6538 3641 6572
rect 3675 6538 3731 6572
rect 3765 6538 3821 6572
rect 3855 6538 3911 6572
rect 3945 6538 4001 6572
rect 4035 6538 4096 6572
rect 3402 6534 4096 6538
rect 3402 6500 3489 6534
rect 3523 6500 3589 6534
rect 3623 6500 3689 6534
rect 3723 6500 3789 6534
rect 3823 6500 3889 6534
rect 3923 6500 3989 6534
rect 4023 6500 4096 6534
rect 3402 6482 4096 6500
rect 3402 6448 3461 6482
rect 3495 6448 3551 6482
rect 3585 6448 3641 6482
rect 3675 6448 3731 6482
rect 3765 6448 3821 6482
rect 3855 6448 3911 6482
rect 3945 6448 4001 6482
rect 4035 6448 4096 6482
rect 3402 6434 4096 6448
rect 3402 6400 3489 6434
rect 3523 6400 3589 6434
rect 3623 6400 3689 6434
rect 3723 6400 3789 6434
rect 3823 6400 3889 6434
rect 3923 6400 3989 6434
rect 4023 6400 4096 6434
rect 3402 6392 4096 6400
rect 3402 6358 3461 6392
rect 3495 6358 3551 6392
rect 3585 6358 3641 6392
rect 3675 6358 3731 6392
rect 3765 6358 3821 6392
rect 3855 6358 3911 6392
rect 3945 6358 4001 6392
rect 4035 6358 4096 6392
rect 3402 6334 4096 6358
rect 3402 6302 3489 6334
rect 3523 6302 3589 6334
rect 3402 6268 3461 6302
rect 3523 6300 3551 6302
rect 3495 6268 3551 6300
rect 3585 6300 3589 6302
rect 3623 6302 3689 6334
rect 3623 6300 3641 6302
rect 3585 6268 3641 6300
rect 3675 6300 3689 6302
rect 3723 6302 3789 6334
rect 3823 6302 3889 6334
rect 3923 6302 3989 6334
rect 4023 6302 4096 6334
rect 3723 6300 3731 6302
rect 3675 6268 3731 6300
rect 3765 6300 3789 6302
rect 3855 6300 3889 6302
rect 3945 6300 3989 6302
rect 3765 6268 3821 6300
rect 3855 6268 3911 6300
rect 3945 6268 4001 6300
rect 4035 6268 4096 6302
rect 3402 6234 4096 6268
rect 3402 6212 3489 6234
rect 3523 6212 3589 6234
rect 3402 6178 3461 6212
rect 3523 6200 3551 6212
rect 3495 6178 3551 6200
rect 3585 6200 3589 6212
rect 3623 6212 3689 6234
rect 3623 6200 3641 6212
rect 3585 6178 3641 6200
rect 3675 6200 3689 6212
rect 3723 6212 3789 6234
rect 3823 6212 3889 6234
rect 3923 6212 3989 6234
rect 4023 6212 4096 6234
rect 3723 6200 3731 6212
rect 3675 6178 3731 6200
rect 3765 6200 3789 6212
rect 3855 6200 3889 6212
rect 3945 6200 3989 6212
rect 3765 6178 3821 6200
rect 3855 6178 3911 6200
rect 3945 6178 4001 6200
rect 4035 6178 4096 6212
rect 3402 6134 4096 6178
rect 3402 6122 3489 6134
rect 3523 6122 3589 6134
rect 3402 6088 3461 6122
rect 3523 6100 3551 6122
rect 3495 6088 3551 6100
rect 3585 6100 3589 6122
rect 3623 6122 3689 6134
rect 3623 6100 3641 6122
rect 3585 6088 3641 6100
rect 3675 6100 3689 6122
rect 3723 6122 3789 6134
rect 3823 6122 3889 6134
rect 3923 6122 3989 6134
rect 4023 6122 4096 6134
rect 3723 6100 3731 6122
rect 3675 6088 3731 6100
rect 3765 6100 3789 6122
rect 3855 6100 3889 6122
rect 3945 6100 3989 6122
rect 3765 6088 3821 6100
rect 3855 6088 3911 6100
rect 3945 6088 4001 6100
rect 4035 6088 4096 6122
rect 3402 6027 4096 6088
rect 4158 6710 4177 6744
rect 4211 6710 4230 6744
rect 4158 6654 4230 6710
rect 4158 6620 4177 6654
rect 4211 6620 4230 6654
rect 4158 6564 4230 6620
rect 4158 6530 4177 6564
rect 4211 6530 4230 6564
rect 4158 6474 4230 6530
rect 4158 6440 4177 6474
rect 4211 6440 4230 6474
rect 4158 6384 4230 6440
rect 4158 6350 4177 6384
rect 4211 6350 4230 6384
rect 4158 6294 4230 6350
rect 4158 6260 4177 6294
rect 4211 6260 4230 6294
rect 4158 6204 4230 6260
rect 4158 6170 4177 6204
rect 4211 6170 4230 6204
rect 4158 6114 4230 6170
rect 4158 6080 4177 6114
rect 4211 6080 4230 6114
rect 3268 5965 3340 6024
rect 4158 6024 4230 6080
rect 4158 5990 4177 6024
rect 4211 5990 4230 6024
rect 4158 5965 4230 5990
rect 3340 5946 4158 5965
rect 3340 5912 3344 5946
rect 3378 5912 3434 5946
rect 3468 5912 3524 5946
rect 3558 5912 3614 5946
rect 3648 5912 3704 5946
rect 3738 5912 3794 5946
rect 3828 5912 3884 5946
rect 3918 5912 3974 5946
rect 4008 5912 4064 5946
rect 4098 5912 4158 5946
rect 3340 5893 4158 5912
rect 4294 6850 4327 6884
rect 4361 6850 4393 6884
rect 4294 6794 4393 6850
rect 4294 6760 4327 6794
rect 4361 6760 4393 6794
rect 4294 6704 4393 6760
rect 4294 6670 4327 6704
rect 4361 6670 4393 6704
rect 4294 6614 4393 6670
rect 4294 6580 4327 6614
rect 4361 6580 4393 6614
rect 4294 6524 4393 6580
rect 4294 6490 4327 6524
rect 4361 6490 4393 6524
rect 4294 6434 4393 6490
rect 4294 6400 4327 6434
rect 4361 6400 4393 6434
rect 4294 6344 4393 6400
rect 4294 6310 4327 6344
rect 4361 6310 4393 6344
rect 4294 6254 4393 6310
rect 4294 6220 4327 6254
rect 4361 6220 4393 6254
rect 4294 6164 4393 6220
rect 4294 6130 4327 6164
rect 4361 6130 4393 6164
rect 4294 6074 4393 6130
rect 4294 6040 4327 6074
rect 4361 6040 4393 6074
rect 4294 5984 4393 6040
rect 4294 5965 4327 5984
rect 4361 5965 4393 5984
rect 3105 5860 3140 5893
rect 3174 5860 3204 5893
rect 3105 5829 3204 5860
rect 4294 5860 4327 5893
rect 4361 5860 4393 5893
rect 4294 5829 4393 5860
rect 3105 5798 4393 5829
rect 3105 5764 3163 5798
rect 3197 5764 3253 5798
rect 3287 5764 3343 5798
rect 3377 5764 3433 5798
rect 3467 5764 3523 5798
rect 3557 5764 3613 5798
rect 3647 5764 3703 5798
rect 3737 5764 3793 5798
rect 3827 5764 3883 5798
rect 3917 5764 3973 5798
rect 4007 5764 4063 5798
rect 4097 5764 4153 5798
rect 4187 5764 4243 5798
rect 4277 5764 4393 5798
rect 3105 5730 4393 5764
rect 4493 6985 5781 7018
rect 4493 6951 4551 6985
rect 4585 6951 4641 6985
rect 4675 6951 4731 6985
rect 4765 6951 4821 6985
rect 4855 6951 4911 6985
rect 4945 6951 5001 6985
rect 5035 6951 5091 6985
rect 5125 6951 5181 6985
rect 5215 6951 5271 6985
rect 5305 6951 5361 6985
rect 5395 6951 5451 6985
rect 5485 6951 5541 6985
rect 5575 6951 5631 6985
rect 5665 6951 5781 6985
rect 4493 6919 5781 6951
rect 4493 6884 4592 6919
rect 4493 6850 4528 6884
rect 4562 6850 4592 6884
rect 5682 6884 5781 6919
rect 4493 6794 4592 6850
rect 4493 6760 4528 6794
rect 4562 6760 4592 6794
rect 4493 6704 4592 6760
rect 4493 6670 4528 6704
rect 4562 6670 4592 6704
rect 4493 6614 4592 6670
rect 4493 6580 4528 6614
rect 4562 6580 4592 6614
rect 4493 6524 4592 6580
rect 4493 6490 4528 6524
rect 4562 6490 4592 6524
rect 4493 6434 4592 6490
rect 4493 6400 4528 6434
rect 4562 6400 4592 6434
rect 4493 6344 4592 6400
rect 4493 6310 4528 6344
rect 4562 6310 4592 6344
rect 4493 6254 4592 6310
rect 4493 6220 4528 6254
rect 4562 6220 4592 6254
rect 4493 6164 4592 6220
rect 4493 6130 4528 6164
rect 4562 6130 4592 6164
rect 4493 6074 4592 6130
rect 4493 6040 4528 6074
rect 4562 6040 4592 6074
rect 4493 5984 4592 6040
rect 4493 5965 4528 5984
rect 4562 5965 4592 5984
rect 4656 6836 5618 6855
rect 4656 6802 4751 6836
rect 4785 6802 4841 6836
rect 4875 6802 4931 6836
rect 4965 6802 5021 6836
rect 5055 6802 5111 6836
rect 5145 6802 5201 6836
rect 5235 6802 5291 6836
rect 5325 6802 5381 6836
rect 5415 6802 5471 6836
rect 5505 6802 5618 6836
rect 4656 6783 5618 6802
rect 4656 6778 4728 6783
rect 4656 6744 4675 6778
rect 4709 6744 4728 6778
rect 4656 6688 4728 6744
rect 5546 6744 5618 6783
rect 4656 6654 4675 6688
rect 4709 6654 4728 6688
rect 4656 6598 4728 6654
rect 4656 6564 4675 6598
rect 4709 6564 4728 6598
rect 4656 6508 4728 6564
rect 4656 6474 4675 6508
rect 4709 6474 4728 6508
rect 4656 6418 4728 6474
rect 4656 6384 4675 6418
rect 4709 6384 4728 6418
rect 4656 6328 4728 6384
rect 4656 6294 4675 6328
rect 4709 6294 4728 6328
rect 4656 6238 4728 6294
rect 4656 6204 4675 6238
rect 4709 6204 4728 6238
rect 4656 6148 4728 6204
rect 4656 6114 4675 6148
rect 4709 6114 4728 6148
rect 4656 6058 4728 6114
rect 4656 6024 4675 6058
rect 4709 6024 4728 6058
rect 4790 6662 5484 6721
rect 4790 6628 4849 6662
rect 4883 6634 4939 6662
rect 4911 6628 4939 6634
rect 4973 6634 5029 6662
rect 4973 6628 4977 6634
rect 4790 6600 4877 6628
rect 4911 6600 4977 6628
rect 5011 6628 5029 6634
rect 5063 6634 5119 6662
rect 5063 6628 5077 6634
rect 5011 6600 5077 6628
rect 5111 6628 5119 6634
rect 5153 6634 5209 6662
rect 5243 6634 5299 6662
rect 5333 6634 5389 6662
rect 5153 6628 5177 6634
rect 5243 6628 5277 6634
rect 5333 6628 5377 6634
rect 5423 6628 5484 6662
rect 5111 6600 5177 6628
rect 5211 6600 5277 6628
rect 5311 6600 5377 6628
rect 5411 6600 5484 6628
rect 4790 6572 5484 6600
rect 4790 6538 4849 6572
rect 4883 6538 4939 6572
rect 4973 6538 5029 6572
rect 5063 6538 5119 6572
rect 5153 6538 5209 6572
rect 5243 6538 5299 6572
rect 5333 6538 5389 6572
rect 5423 6538 5484 6572
rect 4790 6534 5484 6538
rect 4790 6500 4877 6534
rect 4911 6500 4977 6534
rect 5011 6500 5077 6534
rect 5111 6500 5177 6534
rect 5211 6500 5277 6534
rect 5311 6500 5377 6534
rect 5411 6500 5484 6534
rect 4790 6482 5484 6500
rect 4790 6448 4849 6482
rect 4883 6448 4939 6482
rect 4973 6448 5029 6482
rect 5063 6448 5119 6482
rect 5153 6448 5209 6482
rect 5243 6448 5299 6482
rect 5333 6448 5389 6482
rect 5423 6448 5484 6482
rect 4790 6434 5484 6448
rect 4790 6400 4877 6434
rect 4911 6400 4977 6434
rect 5011 6400 5077 6434
rect 5111 6400 5177 6434
rect 5211 6400 5277 6434
rect 5311 6400 5377 6434
rect 5411 6400 5484 6434
rect 4790 6392 5484 6400
rect 4790 6358 4849 6392
rect 4883 6358 4939 6392
rect 4973 6358 5029 6392
rect 5063 6358 5119 6392
rect 5153 6358 5209 6392
rect 5243 6358 5299 6392
rect 5333 6358 5389 6392
rect 5423 6358 5484 6392
rect 4790 6334 5484 6358
rect 4790 6302 4877 6334
rect 4911 6302 4977 6334
rect 4790 6268 4849 6302
rect 4911 6300 4939 6302
rect 4883 6268 4939 6300
rect 4973 6300 4977 6302
rect 5011 6302 5077 6334
rect 5011 6300 5029 6302
rect 4973 6268 5029 6300
rect 5063 6300 5077 6302
rect 5111 6302 5177 6334
rect 5211 6302 5277 6334
rect 5311 6302 5377 6334
rect 5411 6302 5484 6334
rect 5111 6300 5119 6302
rect 5063 6268 5119 6300
rect 5153 6300 5177 6302
rect 5243 6300 5277 6302
rect 5333 6300 5377 6302
rect 5153 6268 5209 6300
rect 5243 6268 5299 6300
rect 5333 6268 5389 6300
rect 5423 6268 5484 6302
rect 4790 6234 5484 6268
rect 4790 6212 4877 6234
rect 4911 6212 4977 6234
rect 4790 6178 4849 6212
rect 4911 6200 4939 6212
rect 4883 6178 4939 6200
rect 4973 6200 4977 6212
rect 5011 6212 5077 6234
rect 5011 6200 5029 6212
rect 4973 6178 5029 6200
rect 5063 6200 5077 6212
rect 5111 6212 5177 6234
rect 5211 6212 5277 6234
rect 5311 6212 5377 6234
rect 5411 6212 5484 6234
rect 5111 6200 5119 6212
rect 5063 6178 5119 6200
rect 5153 6200 5177 6212
rect 5243 6200 5277 6212
rect 5333 6200 5377 6212
rect 5153 6178 5209 6200
rect 5243 6178 5299 6200
rect 5333 6178 5389 6200
rect 5423 6178 5484 6212
rect 4790 6134 5484 6178
rect 4790 6122 4877 6134
rect 4911 6122 4977 6134
rect 4790 6088 4849 6122
rect 4911 6100 4939 6122
rect 4883 6088 4939 6100
rect 4973 6100 4977 6122
rect 5011 6122 5077 6134
rect 5011 6100 5029 6122
rect 4973 6088 5029 6100
rect 5063 6100 5077 6122
rect 5111 6122 5177 6134
rect 5211 6122 5277 6134
rect 5311 6122 5377 6134
rect 5411 6122 5484 6134
rect 5111 6100 5119 6122
rect 5063 6088 5119 6100
rect 5153 6100 5177 6122
rect 5243 6100 5277 6122
rect 5333 6100 5377 6122
rect 5153 6088 5209 6100
rect 5243 6088 5299 6100
rect 5333 6088 5389 6100
rect 5423 6088 5484 6122
rect 4790 6027 5484 6088
rect 5546 6710 5565 6744
rect 5599 6710 5618 6744
rect 5546 6654 5618 6710
rect 5546 6620 5565 6654
rect 5599 6620 5618 6654
rect 5546 6564 5618 6620
rect 5546 6530 5565 6564
rect 5599 6530 5618 6564
rect 5546 6474 5618 6530
rect 5546 6440 5565 6474
rect 5599 6440 5618 6474
rect 5546 6384 5618 6440
rect 5546 6350 5565 6384
rect 5599 6350 5618 6384
rect 5546 6294 5618 6350
rect 5546 6260 5565 6294
rect 5599 6260 5618 6294
rect 5546 6204 5618 6260
rect 5546 6170 5565 6204
rect 5599 6170 5618 6204
rect 5546 6114 5618 6170
rect 5546 6080 5565 6114
rect 5599 6080 5618 6114
rect 4656 5965 4728 6024
rect 5546 6024 5618 6080
rect 5546 5990 5565 6024
rect 5599 5990 5618 6024
rect 5546 5965 5618 5990
rect 4728 5946 5618 5965
rect 4728 5912 4732 5946
rect 4766 5912 4822 5946
rect 4856 5912 4912 5946
rect 4946 5912 5002 5946
rect 5036 5912 5092 5946
rect 5126 5912 5182 5946
rect 5216 5912 5272 5946
rect 5306 5912 5362 5946
rect 5396 5912 5452 5946
rect 5486 5912 5618 5946
rect 4728 5893 5618 5912
rect 5682 6850 5715 6884
rect 5749 6850 5781 6884
rect 5682 6794 5781 6850
rect 5682 6760 5715 6794
rect 5749 6760 5781 6794
rect 5682 6704 5781 6760
rect 5682 6670 5715 6704
rect 5749 6670 5781 6704
rect 5682 6614 5781 6670
rect 5682 6580 5715 6614
rect 5749 6580 5781 6614
rect 5682 6524 5781 6580
rect 5682 6490 5715 6524
rect 5749 6490 5781 6524
rect 5682 6434 5781 6490
rect 5682 6400 5715 6434
rect 5749 6400 5781 6434
rect 5682 6344 5781 6400
rect 5682 6310 5715 6344
rect 5749 6310 5781 6344
rect 5682 6254 5781 6310
rect 5682 6220 5715 6254
rect 5749 6220 5781 6254
rect 5682 6164 5781 6220
rect 5682 6130 5715 6164
rect 5749 6130 5781 6164
rect 5682 6074 5781 6130
rect 5682 6040 5715 6074
rect 5749 6040 5781 6074
rect 5682 5984 5781 6040
rect 5682 5950 5715 5984
rect 5749 5950 5781 5984
rect 5682 5894 5781 5950
rect 4493 5860 4528 5893
rect 4562 5860 4592 5893
rect 4493 5829 4592 5860
rect 5682 5860 5715 5894
rect 5749 5860 5781 5894
rect 5682 5829 5781 5860
rect 4493 5798 4656 5829
rect 4728 5798 5781 5829
rect 4493 5764 4551 5798
rect 4585 5764 4641 5798
rect 4728 5764 4731 5798
rect 4765 5764 4821 5798
rect 4855 5764 4911 5798
rect 4945 5764 5001 5798
rect 5035 5764 5091 5798
rect 5125 5764 5181 5798
rect 5215 5764 5271 5798
rect 5305 5764 5361 5798
rect 5395 5764 5451 5798
rect 5485 5764 5541 5798
rect 5575 5764 5631 5798
rect 5665 5764 5781 5798
rect 4493 5730 4656 5764
rect 4728 5730 5781 5764
rect 5881 6985 6044 7018
rect 6116 6985 7169 7018
rect 5881 6951 5939 6985
rect 5973 6951 6029 6985
rect 6116 6951 6119 6985
rect 6153 6951 6209 6985
rect 6243 6951 6299 6985
rect 6333 6951 6389 6985
rect 6423 6951 6479 6985
rect 6513 6951 6569 6985
rect 6603 6951 6659 6985
rect 6693 6951 6749 6985
rect 6783 6951 6839 6985
rect 6873 6951 6929 6985
rect 6963 6951 7019 6985
rect 7053 6951 7169 6985
rect 5881 6919 6044 6951
rect 6116 6919 7169 6951
rect 5881 6884 5980 6919
rect 5881 6850 5916 6884
rect 5950 6850 5980 6884
rect 7070 6884 7169 6919
rect 5881 6794 5980 6850
rect 5881 6760 5916 6794
rect 5950 6760 5980 6794
rect 5881 6704 5980 6760
rect 5881 6670 5916 6704
rect 5950 6670 5980 6704
rect 5881 6614 5980 6670
rect 5881 6580 5916 6614
rect 5950 6580 5980 6614
rect 5881 6524 5980 6580
rect 5881 6490 5916 6524
rect 5950 6490 5980 6524
rect 5881 6434 5980 6490
rect 5881 6400 5916 6434
rect 5950 6400 5980 6434
rect 5881 6344 5980 6400
rect 5881 6310 5916 6344
rect 5950 6310 5980 6344
rect 5881 6254 5980 6310
rect 5881 6220 5916 6254
rect 5950 6220 5980 6254
rect 5881 6164 5980 6220
rect 5881 6130 5916 6164
rect 5950 6130 5980 6164
rect 5881 6074 5980 6130
rect 5881 6040 5916 6074
rect 5950 6040 5980 6074
rect 5881 5984 5980 6040
rect 5881 5950 5916 5984
rect 5950 5950 5980 5984
rect 5881 5894 5980 5950
rect 5881 5860 5916 5894
rect 5950 5860 5980 5894
rect 6116 6836 7006 6855
rect 6116 6802 6139 6836
rect 6173 6802 6229 6836
rect 6263 6802 6319 6836
rect 6353 6802 6409 6836
rect 6443 6802 6499 6836
rect 6533 6802 6589 6836
rect 6623 6802 6679 6836
rect 6713 6802 6769 6836
rect 6803 6802 6859 6836
rect 6893 6802 7006 6836
rect 6116 6783 7006 6802
rect 6044 6778 6116 6783
rect 6044 6744 6063 6778
rect 6097 6744 6116 6778
rect 6044 6688 6116 6744
rect 6934 6744 7006 6783
rect 6044 6654 6063 6688
rect 6097 6654 6116 6688
rect 6044 6598 6116 6654
rect 6044 6564 6063 6598
rect 6097 6564 6116 6598
rect 6044 6508 6116 6564
rect 6044 6474 6063 6508
rect 6097 6474 6116 6508
rect 6044 6418 6116 6474
rect 6044 6384 6063 6418
rect 6097 6384 6116 6418
rect 6044 6328 6116 6384
rect 6044 6294 6063 6328
rect 6097 6294 6116 6328
rect 6044 6238 6116 6294
rect 6044 6204 6063 6238
rect 6097 6204 6116 6238
rect 6044 6148 6116 6204
rect 6044 6114 6063 6148
rect 6097 6114 6116 6148
rect 6044 6058 6116 6114
rect 6044 6024 6063 6058
rect 6097 6024 6116 6058
rect 6178 6662 6872 6721
rect 6178 6628 6237 6662
rect 6271 6634 6327 6662
rect 6299 6628 6327 6634
rect 6361 6634 6417 6662
rect 6361 6628 6365 6634
rect 6178 6600 6265 6628
rect 6299 6600 6365 6628
rect 6399 6628 6417 6634
rect 6451 6634 6507 6662
rect 6451 6628 6465 6634
rect 6399 6600 6465 6628
rect 6499 6628 6507 6634
rect 6541 6634 6597 6662
rect 6631 6634 6687 6662
rect 6721 6634 6777 6662
rect 6541 6628 6565 6634
rect 6631 6628 6665 6634
rect 6721 6628 6765 6634
rect 6811 6628 6872 6662
rect 6499 6600 6565 6628
rect 6599 6600 6665 6628
rect 6699 6600 6765 6628
rect 6799 6600 6872 6628
rect 6178 6572 6872 6600
rect 6178 6538 6237 6572
rect 6271 6538 6327 6572
rect 6361 6538 6417 6572
rect 6451 6538 6507 6572
rect 6541 6538 6597 6572
rect 6631 6538 6687 6572
rect 6721 6538 6777 6572
rect 6811 6538 6872 6572
rect 6178 6534 6872 6538
rect 6178 6500 6265 6534
rect 6299 6500 6365 6534
rect 6399 6500 6465 6534
rect 6499 6500 6565 6534
rect 6599 6500 6665 6534
rect 6699 6500 6765 6534
rect 6799 6500 6872 6534
rect 6178 6482 6872 6500
rect 6178 6448 6237 6482
rect 6271 6448 6327 6482
rect 6361 6448 6417 6482
rect 6451 6448 6507 6482
rect 6541 6448 6597 6482
rect 6631 6448 6687 6482
rect 6721 6448 6777 6482
rect 6811 6448 6872 6482
rect 6178 6434 6872 6448
rect 6178 6400 6265 6434
rect 6299 6400 6365 6434
rect 6399 6400 6465 6434
rect 6499 6400 6565 6434
rect 6599 6400 6665 6434
rect 6699 6400 6765 6434
rect 6799 6400 6872 6434
rect 6178 6392 6872 6400
rect 6178 6358 6237 6392
rect 6271 6358 6327 6392
rect 6361 6358 6417 6392
rect 6451 6358 6507 6392
rect 6541 6358 6597 6392
rect 6631 6358 6687 6392
rect 6721 6358 6777 6392
rect 6811 6358 6872 6392
rect 6178 6334 6872 6358
rect 6178 6302 6265 6334
rect 6299 6302 6365 6334
rect 6178 6268 6237 6302
rect 6299 6300 6327 6302
rect 6271 6268 6327 6300
rect 6361 6300 6365 6302
rect 6399 6302 6465 6334
rect 6399 6300 6417 6302
rect 6361 6268 6417 6300
rect 6451 6300 6465 6302
rect 6499 6302 6565 6334
rect 6599 6302 6665 6334
rect 6699 6302 6765 6334
rect 6799 6302 6872 6334
rect 6499 6300 6507 6302
rect 6451 6268 6507 6300
rect 6541 6300 6565 6302
rect 6631 6300 6665 6302
rect 6721 6300 6765 6302
rect 6541 6268 6597 6300
rect 6631 6268 6687 6300
rect 6721 6268 6777 6300
rect 6811 6268 6872 6302
rect 6178 6234 6872 6268
rect 6178 6212 6265 6234
rect 6299 6212 6365 6234
rect 6178 6178 6237 6212
rect 6299 6200 6327 6212
rect 6271 6178 6327 6200
rect 6361 6200 6365 6212
rect 6399 6212 6465 6234
rect 6399 6200 6417 6212
rect 6361 6178 6417 6200
rect 6451 6200 6465 6212
rect 6499 6212 6565 6234
rect 6599 6212 6665 6234
rect 6699 6212 6765 6234
rect 6799 6212 6872 6234
rect 6499 6200 6507 6212
rect 6451 6178 6507 6200
rect 6541 6200 6565 6212
rect 6631 6200 6665 6212
rect 6721 6200 6765 6212
rect 6541 6178 6597 6200
rect 6631 6178 6687 6200
rect 6721 6178 6777 6200
rect 6811 6178 6872 6212
rect 6178 6134 6872 6178
rect 6178 6122 6265 6134
rect 6299 6122 6365 6134
rect 6178 6088 6237 6122
rect 6299 6100 6327 6122
rect 6271 6088 6327 6100
rect 6361 6100 6365 6122
rect 6399 6122 6465 6134
rect 6399 6100 6417 6122
rect 6361 6088 6417 6100
rect 6451 6100 6465 6122
rect 6499 6122 6565 6134
rect 6599 6122 6665 6134
rect 6699 6122 6765 6134
rect 6799 6122 6872 6134
rect 6499 6100 6507 6122
rect 6451 6088 6507 6100
rect 6541 6100 6565 6122
rect 6631 6100 6665 6122
rect 6721 6100 6765 6122
rect 6541 6088 6597 6100
rect 6631 6088 6687 6100
rect 6721 6088 6777 6100
rect 6811 6088 6872 6122
rect 6178 6027 6872 6088
rect 6934 6710 6953 6744
rect 6987 6710 7006 6744
rect 6934 6654 7006 6710
rect 6934 6620 6953 6654
rect 6987 6620 7006 6654
rect 6934 6564 7006 6620
rect 6934 6530 6953 6564
rect 6987 6530 7006 6564
rect 6934 6474 7006 6530
rect 6934 6440 6953 6474
rect 6987 6440 7006 6474
rect 6934 6384 7006 6440
rect 6934 6350 6953 6384
rect 6987 6350 7006 6384
rect 6934 6294 7006 6350
rect 6934 6260 6953 6294
rect 6987 6260 7006 6294
rect 6934 6204 7006 6260
rect 6934 6170 6953 6204
rect 6987 6170 7006 6204
rect 6934 6114 7006 6170
rect 6934 6080 6953 6114
rect 6987 6080 7006 6114
rect 6044 5965 6116 6024
rect 6934 6024 7006 6080
rect 6934 5990 6953 6024
rect 6987 5990 7006 6024
rect 6934 5965 7006 5990
rect 6116 5946 7006 5965
rect 6116 5912 6120 5946
rect 6154 5912 6210 5946
rect 6244 5912 6300 5946
rect 6334 5912 6390 5946
rect 6424 5912 6480 5946
rect 6514 5912 6570 5946
rect 6604 5912 6660 5946
rect 6694 5912 6750 5946
rect 6784 5912 6840 5946
rect 6874 5912 7006 5946
rect 6116 5893 7006 5912
rect 7070 6850 7103 6884
rect 7137 6850 7169 6884
rect 7070 6794 7169 6850
rect 7070 6760 7103 6794
rect 7137 6760 7169 6794
rect 7070 6704 7169 6760
rect 7070 6670 7103 6704
rect 7137 6670 7169 6704
rect 7070 6614 7169 6670
rect 7070 6580 7103 6614
rect 7137 6580 7169 6614
rect 7070 6524 7169 6580
rect 7070 6490 7103 6524
rect 7137 6490 7169 6524
rect 7070 6434 7169 6490
rect 7070 6400 7103 6434
rect 7137 6400 7169 6434
rect 7070 6344 7169 6400
rect 7070 6310 7103 6344
rect 7137 6310 7169 6344
rect 7070 6254 7169 6310
rect 7070 6220 7103 6254
rect 7137 6220 7169 6254
rect 7070 6164 7169 6220
rect 7070 6130 7103 6164
rect 7137 6130 7169 6164
rect 7070 6074 7169 6130
rect 7070 6040 7103 6074
rect 7137 6040 7169 6074
rect 7070 5984 7169 6040
rect 7070 5950 7103 5984
rect 7137 5950 7169 5984
rect 7070 5894 7169 5950
rect 5881 5829 5980 5860
rect 7070 5860 7103 5894
rect 7137 5860 7169 5894
rect 7070 5829 7169 5860
rect 5881 5798 6044 5829
rect 6116 5798 7169 5829
rect 5881 5764 5939 5798
rect 5973 5764 6029 5798
rect 6116 5764 6119 5798
rect 6153 5764 6209 5798
rect 6243 5764 6299 5798
rect 6333 5764 6389 5798
rect 6423 5764 6479 5798
rect 6513 5764 6569 5798
rect 6603 5764 6659 5798
rect 6693 5764 6749 5798
rect 6783 5764 6839 5798
rect 6873 5764 6929 5798
rect 6963 5764 7019 5798
rect 7053 5764 7169 5798
rect 5881 5730 6044 5764
rect 6116 5730 7169 5764
rect 329 5597 1382 5630
rect 1454 5597 1617 5630
rect 329 5563 387 5597
rect 421 5563 477 5597
rect 511 5563 567 5597
rect 601 5563 657 5597
rect 691 5563 747 5597
rect 781 5563 837 5597
rect 871 5563 927 5597
rect 961 5563 1017 5597
rect 1051 5563 1107 5597
rect 1141 5563 1197 5597
rect 1231 5563 1287 5597
rect 1321 5563 1377 5597
rect 1454 5563 1467 5597
rect 1501 5563 1617 5597
rect 329 5531 1382 5563
rect 1454 5531 1617 5563
rect 329 5496 428 5531
rect 329 5462 364 5496
rect 398 5462 428 5496
rect 1518 5496 1617 5531
rect 329 5406 428 5462
rect 329 5372 364 5406
rect 398 5372 428 5406
rect 329 5316 428 5372
rect 329 5282 364 5316
rect 398 5282 428 5316
rect 329 5226 428 5282
rect 329 5192 364 5226
rect 398 5192 428 5226
rect 329 5136 428 5192
rect 329 5102 364 5136
rect 398 5102 428 5136
rect 329 5046 428 5102
rect 329 5012 364 5046
rect 398 5012 428 5046
rect 329 4956 428 5012
rect 329 4922 364 4956
rect 398 4922 428 4956
rect 329 4866 428 4922
rect 329 4832 364 4866
rect 398 4832 428 4866
rect 329 4776 428 4832
rect 329 4742 364 4776
rect 398 4742 428 4776
rect 329 4686 428 4742
rect 329 4652 364 4686
rect 398 4652 428 4686
rect 329 4596 428 4652
rect 329 4562 364 4596
rect 398 4562 428 4596
rect 329 4506 428 4562
rect 329 4472 364 4506
rect 398 4472 428 4506
rect 492 5448 1382 5467
rect 492 5414 587 5448
rect 621 5414 677 5448
rect 711 5414 767 5448
rect 801 5414 857 5448
rect 891 5414 947 5448
rect 981 5414 1037 5448
rect 1071 5414 1127 5448
rect 1161 5414 1217 5448
rect 1251 5414 1307 5448
rect 1341 5414 1382 5448
rect 492 5395 1382 5414
rect 492 5390 564 5395
rect 492 5356 511 5390
rect 545 5356 564 5390
rect 492 5300 564 5356
rect 1382 5356 1454 5395
rect 492 5266 511 5300
rect 545 5266 564 5300
rect 492 5210 564 5266
rect 492 5176 511 5210
rect 545 5176 564 5210
rect 492 5120 564 5176
rect 492 5086 511 5120
rect 545 5086 564 5120
rect 492 5030 564 5086
rect 492 4996 511 5030
rect 545 4996 564 5030
rect 492 4940 564 4996
rect 492 4906 511 4940
rect 545 4906 564 4940
rect 492 4850 564 4906
rect 492 4816 511 4850
rect 545 4816 564 4850
rect 492 4760 564 4816
rect 492 4726 511 4760
rect 545 4726 564 4760
rect 492 4670 564 4726
rect 492 4636 511 4670
rect 545 4636 564 4670
rect 626 5274 1320 5333
rect 626 5240 685 5274
rect 719 5246 775 5274
rect 747 5240 775 5246
rect 809 5246 865 5274
rect 809 5240 813 5246
rect 626 5212 713 5240
rect 747 5212 813 5240
rect 847 5240 865 5246
rect 899 5246 955 5274
rect 899 5240 913 5246
rect 847 5212 913 5240
rect 947 5240 955 5246
rect 989 5246 1045 5274
rect 1079 5246 1135 5274
rect 1169 5246 1225 5274
rect 989 5240 1013 5246
rect 1079 5240 1113 5246
rect 1169 5240 1213 5246
rect 1259 5240 1320 5274
rect 947 5212 1013 5240
rect 1047 5212 1113 5240
rect 1147 5212 1213 5240
rect 1247 5212 1320 5240
rect 626 5184 1320 5212
rect 626 5150 685 5184
rect 719 5150 775 5184
rect 809 5150 865 5184
rect 899 5150 955 5184
rect 989 5150 1045 5184
rect 1079 5150 1135 5184
rect 1169 5150 1225 5184
rect 1259 5150 1320 5184
rect 626 5146 1320 5150
rect 626 5112 713 5146
rect 747 5112 813 5146
rect 847 5112 913 5146
rect 947 5112 1013 5146
rect 1047 5112 1113 5146
rect 1147 5112 1213 5146
rect 1247 5112 1320 5146
rect 626 5094 1320 5112
rect 626 5060 685 5094
rect 719 5060 775 5094
rect 809 5060 865 5094
rect 899 5060 955 5094
rect 989 5060 1045 5094
rect 1079 5060 1135 5094
rect 1169 5060 1225 5094
rect 1259 5060 1320 5094
rect 626 5046 1320 5060
rect 626 5012 713 5046
rect 747 5012 813 5046
rect 847 5012 913 5046
rect 947 5012 1013 5046
rect 1047 5012 1113 5046
rect 1147 5012 1213 5046
rect 1247 5012 1320 5046
rect 626 5004 1320 5012
rect 626 4970 685 5004
rect 719 4970 775 5004
rect 809 4970 865 5004
rect 899 4970 955 5004
rect 989 4970 1045 5004
rect 1079 4970 1135 5004
rect 1169 4970 1225 5004
rect 1259 4970 1320 5004
rect 626 4946 1320 4970
rect 626 4914 713 4946
rect 747 4914 813 4946
rect 626 4880 685 4914
rect 747 4912 775 4914
rect 719 4880 775 4912
rect 809 4912 813 4914
rect 847 4914 913 4946
rect 847 4912 865 4914
rect 809 4880 865 4912
rect 899 4912 913 4914
rect 947 4914 1013 4946
rect 1047 4914 1113 4946
rect 1147 4914 1213 4946
rect 1247 4914 1320 4946
rect 947 4912 955 4914
rect 899 4880 955 4912
rect 989 4912 1013 4914
rect 1079 4912 1113 4914
rect 1169 4912 1213 4914
rect 989 4880 1045 4912
rect 1079 4880 1135 4912
rect 1169 4880 1225 4912
rect 1259 4880 1320 4914
rect 626 4846 1320 4880
rect 626 4824 713 4846
rect 747 4824 813 4846
rect 626 4790 685 4824
rect 747 4812 775 4824
rect 719 4790 775 4812
rect 809 4812 813 4824
rect 847 4824 913 4846
rect 847 4812 865 4824
rect 809 4790 865 4812
rect 899 4812 913 4824
rect 947 4824 1013 4846
rect 1047 4824 1113 4846
rect 1147 4824 1213 4846
rect 1247 4824 1320 4846
rect 947 4812 955 4824
rect 899 4790 955 4812
rect 989 4812 1013 4824
rect 1079 4812 1113 4824
rect 1169 4812 1213 4824
rect 989 4790 1045 4812
rect 1079 4790 1135 4812
rect 1169 4790 1225 4812
rect 1259 4790 1320 4824
rect 626 4746 1320 4790
rect 626 4734 713 4746
rect 747 4734 813 4746
rect 626 4700 685 4734
rect 747 4712 775 4734
rect 719 4700 775 4712
rect 809 4712 813 4734
rect 847 4734 913 4746
rect 847 4712 865 4734
rect 809 4700 865 4712
rect 899 4712 913 4734
rect 947 4734 1013 4746
rect 1047 4734 1113 4746
rect 1147 4734 1213 4746
rect 1247 4734 1320 4746
rect 947 4712 955 4734
rect 899 4700 955 4712
rect 989 4712 1013 4734
rect 1079 4712 1113 4734
rect 1169 4712 1213 4734
rect 989 4700 1045 4712
rect 1079 4700 1135 4712
rect 1169 4700 1225 4712
rect 1259 4700 1320 4734
rect 626 4639 1320 4700
rect 1382 5322 1401 5356
rect 1435 5322 1454 5356
rect 1382 5266 1454 5322
rect 1382 5232 1401 5266
rect 1435 5232 1454 5266
rect 1382 5176 1454 5232
rect 1382 5142 1401 5176
rect 1435 5142 1454 5176
rect 1382 5086 1454 5142
rect 1382 5052 1401 5086
rect 1435 5052 1454 5086
rect 1382 4996 1454 5052
rect 1382 4962 1401 4996
rect 1435 4962 1454 4996
rect 1382 4906 1454 4962
rect 1382 4872 1401 4906
rect 1435 4872 1454 4906
rect 1382 4816 1454 4872
rect 1382 4782 1401 4816
rect 1435 4782 1454 4816
rect 1382 4726 1454 4782
rect 1382 4692 1401 4726
rect 1435 4692 1454 4726
rect 492 4577 564 4636
rect 1382 4636 1454 4692
rect 1382 4602 1401 4636
rect 1435 4602 1454 4636
rect 1382 4577 1454 4602
rect 492 4558 1382 4577
rect 492 4524 568 4558
rect 602 4524 658 4558
rect 692 4524 748 4558
rect 782 4524 838 4558
rect 872 4524 928 4558
rect 962 4524 1018 4558
rect 1052 4524 1108 4558
rect 1142 4524 1198 4558
rect 1232 4524 1288 4558
rect 1322 4524 1382 4558
rect 492 4505 1382 4524
rect 1518 5462 1551 5496
rect 1585 5462 1617 5496
rect 1518 5406 1617 5462
rect 1518 5372 1551 5406
rect 1585 5372 1617 5406
rect 1518 5316 1617 5372
rect 1518 5282 1551 5316
rect 1585 5282 1617 5316
rect 1518 5226 1617 5282
rect 1518 5192 1551 5226
rect 1585 5192 1617 5226
rect 1518 5136 1617 5192
rect 1518 5102 1551 5136
rect 1585 5102 1617 5136
rect 1518 5046 1617 5102
rect 1518 5012 1551 5046
rect 1585 5012 1617 5046
rect 1518 4956 1617 5012
rect 1518 4922 1551 4956
rect 1585 4922 1617 4956
rect 1518 4866 1617 4922
rect 1518 4832 1551 4866
rect 1585 4832 1617 4866
rect 1518 4776 1617 4832
rect 1518 4742 1551 4776
rect 1585 4742 1617 4776
rect 1518 4686 1617 4742
rect 1518 4652 1551 4686
rect 1585 4652 1617 4686
rect 1518 4596 1617 4652
rect 1518 4562 1551 4596
rect 1585 4562 1617 4596
rect 1518 4506 1617 4562
rect 329 4441 428 4472
rect 1518 4472 1551 4506
rect 1585 4472 1617 4506
rect 1518 4441 1617 4472
rect 329 4410 1382 4441
rect 1454 4410 1617 4441
rect 329 4376 387 4410
rect 421 4376 477 4410
rect 511 4376 567 4410
rect 601 4376 657 4410
rect 691 4376 747 4410
rect 781 4376 837 4410
rect 871 4376 927 4410
rect 961 4376 1017 4410
rect 1051 4376 1107 4410
rect 1141 4376 1197 4410
rect 1231 4376 1287 4410
rect 1321 4376 1377 4410
rect 1454 4376 1467 4410
rect 1501 4376 1617 4410
rect 329 4342 1382 4376
rect 1454 4342 1617 4376
rect 1717 5597 2770 5630
rect 2842 5597 3005 5630
rect 1717 5563 1775 5597
rect 1809 5563 1865 5597
rect 1899 5563 1955 5597
rect 1989 5563 2045 5597
rect 2079 5563 2135 5597
rect 2169 5563 2225 5597
rect 2259 5563 2315 5597
rect 2349 5563 2405 5597
rect 2439 5563 2495 5597
rect 2529 5563 2585 5597
rect 2619 5563 2675 5597
rect 2709 5563 2765 5597
rect 2842 5563 2855 5597
rect 2889 5563 3005 5597
rect 1717 5531 2770 5563
rect 2842 5531 3005 5563
rect 1717 5496 1816 5531
rect 1717 5462 1752 5496
rect 1786 5462 1816 5496
rect 2906 5496 3005 5531
rect 1717 5406 1816 5462
rect 1717 5372 1752 5406
rect 1786 5372 1816 5406
rect 1717 5316 1816 5372
rect 1717 5282 1752 5316
rect 1786 5282 1816 5316
rect 1717 5226 1816 5282
rect 1717 5192 1752 5226
rect 1786 5192 1816 5226
rect 1717 5136 1816 5192
rect 1717 5102 1752 5136
rect 1786 5102 1816 5136
rect 1717 5046 1816 5102
rect 1717 5012 1752 5046
rect 1786 5012 1816 5046
rect 1717 4956 1816 5012
rect 1717 4922 1752 4956
rect 1786 4922 1816 4956
rect 1717 4866 1816 4922
rect 1717 4832 1752 4866
rect 1786 4832 1816 4866
rect 1717 4776 1816 4832
rect 1717 4742 1752 4776
rect 1786 4742 1816 4776
rect 1717 4686 1816 4742
rect 1717 4652 1752 4686
rect 1786 4652 1816 4686
rect 1717 4596 1816 4652
rect 1717 4562 1752 4596
rect 1786 4562 1816 4596
rect 1717 4506 1816 4562
rect 1717 4472 1752 4506
rect 1786 4472 1816 4506
rect 1880 5448 2770 5467
rect 1880 5414 1975 5448
rect 2009 5414 2065 5448
rect 2099 5414 2155 5448
rect 2189 5414 2245 5448
rect 2279 5414 2335 5448
rect 2369 5414 2425 5448
rect 2459 5414 2515 5448
rect 2549 5414 2605 5448
rect 2639 5414 2695 5448
rect 2729 5414 2770 5448
rect 1880 5395 2770 5414
rect 1880 5390 1952 5395
rect 1880 5356 1899 5390
rect 1933 5356 1952 5390
rect 1880 5300 1952 5356
rect 2770 5356 2842 5395
rect 1880 5266 1899 5300
rect 1933 5266 1952 5300
rect 1880 5210 1952 5266
rect 1880 5176 1899 5210
rect 1933 5176 1952 5210
rect 1880 5120 1952 5176
rect 1880 5086 1899 5120
rect 1933 5086 1952 5120
rect 1880 5030 1952 5086
rect 1880 4996 1899 5030
rect 1933 4996 1952 5030
rect 1880 4940 1952 4996
rect 1880 4906 1899 4940
rect 1933 4906 1952 4940
rect 1880 4850 1952 4906
rect 1880 4816 1899 4850
rect 1933 4816 1952 4850
rect 1880 4760 1952 4816
rect 1880 4726 1899 4760
rect 1933 4726 1952 4760
rect 1880 4670 1952 4726
rect 1880 4636 1899 4670
rect 1933 4636 1952 4670
rect 2014 5274 2708 5333
rect 2014 5240 2073 5274
rect 2107 5246 2163 5274
rect 2135 5240 2163 5246
rect 2197 5246 2253 5274
rect 2197 5240 2201 5246
rect 2014 5212 2101 5240
rect 2135 5212 2201 5240
rect 2235 5240 2253 5246
rect 2287 5246 2343 5274
rect 2287 5240 2301 5246
rect 2235 5212 2301 5240
rect 2335 5240 2343 5246
rect 2377 5246 2433 5274
rect 2467 5246 2523 5274
rect 2557 5246 2613 5274
rect 2377 5240 2401 5246
rect 2467 5240 2501 5246
rect 2557 5240 2601 5246
rect 2647 5240 2708 5274
rect 2335 5212 2401 5240
rect 2435 5212 2501 5240
rect 2535 5212 2601 5240
rect 2635 5212 2708 5240
rect 2014 5184 2708 5212
rect 2014 5150 2073 5184
rect 2107 5150 2163 5184
rect 2197 5150 2253 5184
rect 2287 5150 2343 5184
rect 2377 5150 2433 5184
rect 2467 5150 2523 5184
rect 2557 5150 2613 5184
rect 2647 5150 2708 5184
rect 2014 5146 2708 5150
rect 2014 5112 2101 5146
rect 2135 5112 2201 5146
rect 2235 5112 2301 5146
rect 2335 5112 2401 5146
rect 2435 5112 2501 5146
rect 2535 5112 2601 5146
rect 2635 5112 2708 5146
rect 2014 5094 2708 5112
rect 2014 5060 2073 5094
rect 2107 5060 2163 5094
rect 2197 5060 2253 5094
rect 2287 5060 2343 5094
rect 2377 5060 2433 5094
rect 2467 5060 2523 5094
rect 2557 5060 2613 5094
rect 2647 5060 2708 5094
rect 2014 5046 2708 5060
rect 2014 5012 2101 5046
rect 2135 5012 2201 5046
rect 2235 5012 2301 5046
rect 2335 5012 2401 5046
rect 2435 5012 2501 5046
rect 2535 5012 2601 5046
rect 2635 5012 2708 5046
rect 2014 5004 2708 5012
rect 2014 4970 2073 5004
rect 2107 4970 2163 5004
rect 2197 4970 2253 5004
rect 2287 4970 2343 5004
rect 2377 4970 2433 5004
rect 2467 4970 2523 5004
rect 2557 4970 2613 5004
rect 2647 4970 2708 5004
rect 2014 4946 2708 4970
rect 2014 4914 2101 4946
rect 2135 4914 2201 4946
rect 2014 4880 2073 4914
rect 2135 4912 2163 4914
rect 2107 4880 2163 4912
rect 2197 4912 2201 4914
rect 2235 4914 2301 4946
rect 2235 4912 2253 4914
rect 2197 4880 2253 4912
rect 2287 4912 2301 4914
rect 2335 4914 2401 4946
rect 2435 4914 2501 4946
rect 2535 4914 2601 4946
rect 2635 4914 2708 4946
rect 2335 4912 2343 4914
rect 2287 4880 2343 4912
rect 2377 4912 2401 4914
rect 2467 4912 2501 4914
rect 2557 4912 2601 4914
rect 2377 4880 2433 4912
rect 2467 4880 2523 4912
rect 2557 4880 2613 4912
rect 2647 4880 2708 4914
rect 2014 4846 2708 4880
rect 2014 4824 2101 4846
rect 2135 4824 2201 4846
rect 2014 4790 2073 4824
rect 2135 4812 2163 4824
rect 2107 4790 2163 4812
rect 2197 4812 2201 4824
rect 2235 4824 2301 4846
rect 2235 4812 2253 4824
rect 2197 4790 2253 4812
rect 2287 4812 2301 4824
rect 2335 4824 2401 4846
rect 2435 4824 2501 4846
rect 2535 4824 2601 4846
rect 2635 4824 2708 4846
rect 2335 4812 2343 4824
rect 2287 4790 2343 4812
rect 2377 4812 2401 4824
rect 2467 4812 2501 4824
rect 2557 4812 2601 4824
rect 2377 4790 2433 4812
rect 2467 4790 2523 4812
rect 2557 4790 2613 4812
rect 2647 4790 2708 4824
rect 2014 4746 2708 4790
rect 2014 4734 2101 4746
rect 2135 4734 2201 4746
rect 2014 4700 2073 4734
rect 2135 4712 2163 4734
rect 2107 4700 2163 4712
rect 2197 4712 2201 4734
rect 2235 4734 2301 4746
rect 2235 4712 2253 4734
rect 2197 4700 2253 4712
rect 2287 4712 2301 4734
rect 2335 4734 2401 4746
rect 2435 4734 2501 4746
rect 2535 4734 2601 4746
rect 2635 4734 2708 4746
rect 2335 4712 2343 4734
rect 2287 4700 2343 4712
rect 2377 4712 2401 4734
rect 2467 4712 2501 4734
rect 2557 4712 2601 4734
rect 2377 4700 2433 4712
rect 2467 4700 2523 4712
rect 2557 4700 2613 4712
rect 2647 4700 2708 4734
rect 2014 4639 2708 4700
rect 2770 5322 2789 5356
rect 2823 5322 2842 5356
rect 2770 5266 2842 5322
rect 2770 5232 2789 5266
rect 2823 5232 2842 5266
rect 2770 5176 2842 5232
rect 2770 5142 2789 5176
rect 2823 5142 2842 5176
rect 2770 5086 2842 5142
rect 2770 5052 2789 5086
rect 2823 5052 2842 5086
rect 2770 4996 2842 5052
rect 2770 4962 2789 4996
rect 2823 4962 2842 4996
rect 2770 4906 2842 4962
rect 2770 4872 2789 4906
rect 2823 4872 2842 4906
rect 2770 4816 2842 4872
rect 2770 4782 2789 4816
rect 2823 4782 2842 4816
rect 2770 4726 2842 4782
rect 2770 4692 2789 4726
rect 2823 4692 2842 4726
rect 1880 4577 1952 4636
rect 2770 4636 2842 4692
rect 2770 4602 2789 4636
rect 2823 4602 2842 4636
rect 2770 4577 2842 4602
rect 1880 4558 2770 4577
rect 1880 4524 1956 4558
rect 1990 4524 2046 4558
rect 2080 4524 2136 4558
rect 2170 4524 2226 4558
rect 2260 4524 2316 4558
rect 2350 4524 2406 4558
rect 2440 4524 2496 4558
rect 2530 4524 2586 4558
rect 2620 4524 2676 4558
rect 2710 4524 2770 4558
rect 1880 4505 2770 4524
rect 2906 5462 2939 5496
rect 2973 5462 3005 5496
rect 2906 5406 3005 5462
rect 2906 5372 2939 5406
rect 2973 5372 3005 5406
rect 2906 5316 3005 5372
rect 2906 5282 2939 5316
rect 2973 5282 3005 5316
rect 2906 5226 3005 5282
rect 2906 5192 2939 5226
rect 2973 5192 3005 5226
rect 2906 5136 3005 5192
rect 2906 5102 2939 5136
rect 2973 5102 3005 5136
rect 2906 5046 3005 5102
rect 2906 5012 2939 5046
rect 2973 5012 3005 5046
rect 2906 4956 3005 5012
rect 2906 4922 2939 4956
rect 2973 4922 3005 4956
rect 2906 4866 3005 4922
rect 2906 4832 2939 4866
rect 2973 4832 3005 4866
rect 2906 4776 3005 4832
rect 2906 4742 2939 4776
rect 2973 4742 3005 4776
rect 2906 4686 3005 4742
rect 2906 4652 2939 4686
rect 2973 4652 3005 4686
rect 2906 4596 3005 4652
rect 2906 4562 2939 4596
rect 2973 4562 3005 4596
rect 2906 4506 3005 4562
rect 1717 4441 1816 4472
rect 2906 4472 2939 4506
rect 2973 4472 3005 4506
rect 2906 4441 3005 4472
rect 1717 4410 2770 4441
rect 2842 4410 3005 4441
rect 1717 4376 1775 4410
rect 1809 4376 1865 4410
rect 1899 4376 1955 4410
rect 1989 4376 2045 4410
rect 2079 4376 2135 4410
rect 2169 4376 2225 4410
rect 2259 4376 2315 4410
rect 2349 4376 2405 4410
rect 2439 4376 2495 4410
rect 2529 4376 2585 4410
rect 2619 4376 2675 4410
rect 2709 4376 2765 4410
rect 2842 4376 2855 4410
rect 2889 4376 3005 4410
rect 1717 4342 2770 4376
rect 2842 4342 3005 4376
rect 3105 5597 3268 5630
rect 3340 5597 4158 5630
rect 4230 5597 4393 5630
rect 3105 5563 3163 5597
rect 3197 5563 3253 5597
rect 3340 5563 3343 5597
rect 3377 5563 3433 5597
rect 3467 5563 3523 5597
rect 3557 5563 3613 5597
rect 3647 5563 3703 5597
rect 3737 5563 3793 5597
rect 3827 5563 3883 5597
rect 3917 5563 3973 5597
rect 4007 5563 4063 5597
rect 4097 5563 4153 5597
rect 4230 5563 4243 5597
rect 4277 5563 4393 5597
rect 3105 5531 3268 5563
rect 3340 5531 4158 5563
rect 4230 5531 4393 5563
rect 3105 5496 3204 5531
rect 3105 5467 3140 5496
rect 3174 5467 3204 5496
rect 4294 5496 4393 5531
rect 4294 5467 4327 5496
rect 4361 5467 4393 5496
rect 3105 5372 3140 5395
rect 3174 5372 3204 5395
rect 3105 5316 3204 5372
rect 3105 5282 3140 5316
rect 3174 5282 3204 5316
rect 3105 5226 3204 5282
rect 3105 5192 3140 5226
rect 3174 5192 3204 5226
rect 3105 5136 3204 5192
rect 3105 5102 3140 5136
rect 3174 5102 3204 5136
rect 3105 5046 3204 5102
rect 3105 5012 3140 5046
rect 3174 5012 3204 5046
rect 3105 4956 3204 5012
rect 3105 4922 3140 4956
rect 3174 4922 3204 4956
rect 3105 4866 3204 4922
rect 3105 4832 3140 4866
rect 3174 4832 3204 4866
rect 3105 4776 3204 4832
rect 3105 4742 3140 4776
rect 3174 4742 3204 4776
rect 3105 4686 3204 4742
rect 3105 4652 3140 4686
rect 3174 4652 3204 4686
rect 3105 4596 3204 4652
rect 3105 4577 3140 4596
rect 3174 4577 3204 4596
rect 3340 5448 4158 5467
rect 3340 5414 3363 5448
rect 3397 5414 3453 5448
rect 3487 5414 3543 5448
rect 3577 5414 3633 5448
rect 3667 5414 3723 5448
rect 3757 5414 3813 5448
rect 3847 5414 3903 5448
rect 3937 5414 3993 5448
rect 4027 5414 4083 5448
rect 4117 5414 4158 5448
rect 3340 5395 4158 5414
rect 3268 5390 3340 5395
rect 3268 5356 3287 5390
rect 3321 5356 3340 5390
rect 3268 5300 3340 5356
rect 4158 5356 4230 5395
rect 3268 5266 3287 5300
rect 3321 5266 3340 5300
rect 3268 5210 3340 5266
rect 3268 5176 3287 5210
rect 3321 5176 3340 5210
rect 3268 5120 3340 5176
rect 3268 5086 3287 5120
rect 3321 5086 3340 5120
rect 3268 5030 3340 5086
rect 3268 4996 3287 5030
rect 3321 4996 3340 5030
rect 3268 4940 3340 4996
rect 3268 4906 3287 4940
rect 3321 4906 3340 4940
rect 3268 4850 3340 4906
rect 3268 4816 3287 4850
rect 3321 4816 3340 4850
rect 3268 4760 3340 4816
rect 3268 4726 3287 4760
rect 3321 4726 3340 4760
rect 3268 4670 3340 4726
rect 3268 4636 3287 4670
rect 3321 4636 3340 4670
rect 3402 5274 4096 5333
rect 3402 5240 3461 5274
rect 3495 5246 3551 5274
rect 3523 5240 3551 5246
rect 3585 5246 3641 5274
rect 3585 5240 3589 5246
rect 3402 5212 3489 5240
rect 3523 5212 3589 5240
rect 3623 5240 3641 5246
rect 3675 5246 3731 5274
rect 3675 5240 3689 5246
rect 3623 5212 3689 5240
rect 3723 5240 3731 5246
rect 3765 5246 3821 5274
rect 3855 5246 3911 5274
rect 3945 5246 4001 5274
rect 3765 5240 3789 5246
rect 3855 5240 3889 5246
rect 3945 5240 3989 5246
rect 4035 5240 4096 5274
rect 3723 5212 3789 5240
rect 3823 5212 3889 5240
rect 3923 5212 3989 5240
rect 4023 5212 4096 5240
rect 3402 5184 4096 5212
rect 3402 5150 3461 5184
rect 3495 5150 3551 5184
rect 3585 5150 3641 5184
rect 3675 5150 3731 5184
rect 3765 5150 3821 5184
rect 3855 5150 3911 5184
rect 3945 5150 4001 5184
rect 4035 5150 4096 5184
rect 3402 5146 4096 5150
rect 3402 5112 3489 5146
rect 3523 5112 3589 5146
rect 3623 5112 3689 5146
rect 3723 5112 3789 5146
rect 3823 5112 3889 5146
rect 3923 5112 3989 5146
rect 4023 5112 4096 5146
rect 3402 5094 4096 5112
rect 3402 5060 3461 5094
rect 3495 5060 3551 5094
rect 3585 5060 3641 5094
rect 3675 5060 3731 5094
rect 3765 5060 3821 5094
rect 3855 5060 3911 5094
rect 3945 5060 4001 5094
rect 4035 5060 4096 5094
rect 3402 5046 4096 5060
rect 3402 5012 3489 5046
rect 3523 5012 3589 5046
rect 3623 5012 3689 5046
rect 3723 5012 3789 5046
rect 3823 5012 3889 5046
rect 3923 5012 3989 5046
rect 4023 5012 4096 5046
rect 3402 5004 4096 5012
rect 3402 4970 3461 5004
rect 3495 4970 3551 5004
rect 3585 4970 3641 5004
rect 3675 4970 3731 5004
rect 3765 4970 3821 5004
rect 3855 4970 3911 5004
rect 3945 4970 4001 5004
rect 4035 4970 4096 5004
rect 3402 4946 4096 4970
rect 3402 4914 3489 4946
rect 3523 4914 3589 4946
rect 3402 4880 3461 4914
rect 3523 4912 3551 4914
rect 3495 4880 3551 4912
rect 3585 4912 3589 4914
rect 3623 4914 3689 4946
rect 3623 4912 3641 4914
rect 3585 4880 3641 4912
rect 3675 4912 3689 4914
rect 3723 4914 3789 4946
rect 3823 4914 3889 4946
rect 3923 4914 3989 4946
rect 4023 4914 4096 4946
rect 3723 4912 3731 4914
rect 3675 4880 3731 4912
rect 3765 4912 3789 4914
rect 3855 4912 3889 4914
rect 3945 4912 3989 4914
rect 3765 4880 3821 4912
rect 3855 4880 3911 4912
rect 3945 4880 4001 4912
rect 4035 4880 4096 4914
rect 3402 4846 4096 4880
rect 3402 4824 3489 4846
rect 3523 4824 3589 4846
rect 3402 4790 3461 4824
rect 3523 4812 3551 4824
rect 3495 4790 3551 4812
rect 3585 4812 3589 4824
rect 3623 4824 3689 4846
rect 3623 4812 3641 4824
rect 3585 4790 3641 4812
rect 3675 4812 3689 4824
rect 3723 4824 3789 4846
rect 3823 4824 3889 4846
rect 3923 4824 3989 4846
rect 4023 4824 4096 4846
rect 3723 4812 3731 4824
rect 3675 4790 3731 4812
rect 3765 4812 3789 4824
rect 3855 4812 3889 4824
rect 3945 4812 3989 4824
rect 3765 4790 3821 4812
rect 3855 4790 3911 4812
rect 3945 4790 4001 4812
rect 4035 4790 4096 4824
rect 3402 4746 4096 4790
rect 3402 4734 3489 4746
rect 3523 4734 3589 4746
rect 3402 4700 3461 4734
rect 3523 4712 3551 4734
rect 3495 4700 3551 4712
rect 3585 4712 3589 4734
rect 3623 4734 3689 4746
rect 3623 4712 3641 4734
rect 3585 4700 3641 4712
rect 3675 4712 3689 4734
rect 3723 4734 3789 4746
rect 3823 4734 3889 4746
rect 3923 4734 3989 4746
rect 4023 4734 4096 4746
rect 3723 4712 3731 4734
rect 3675 4700 3731 4712
rect 3765 4712 3789 4734
rect 3855 4712 3889 4734
rect 3945 4712 3989 4734
rect 3765 4700 3821 4712
rect 3855 4700 3911 4712
rect 3945 4700 4001 4712
rect 4035 4700 4096 4734
rect 3402 4639 4096 4700
rect 4158 5322 4177 5356
rect 4211 5322 4230 5356
rect 4158 5266 4230 5322
rect 4158 5232 4177 5266
rect 4211 5232 4230 5266
rect 4158 5176 4230 5232
rect 4158 5142 4177 5176
rect 4211 5142 4230 5176
rect 4158 5086 4230 5142
rect 4158 5052 4177 5086
rect 4211 5052 4230 5086
rect 4158 4996 4230 5052
rect 4158 4962 4177 4996
rect 4211 4962 4230 4996
rect 4158 4906 4230 4962
rect 4158 4872 4177 4906
rect 4211 4872 4230 4906
rect 4158 4816 4230 4872
rect 4158 4782 4177 4816
rect 4211 4782 4230 4816
rect 4158 4726 4230 4782
rect 4158 4692 4177 4726
rect 4211 4692 4230 4726
rect 3268 4577 3340 4636
rect 4158 4636 4230 4692
rect 4158 4602 4177 4636
rect 4211 4602 4230 4636
rect 4158 4577 4230 4602
rect 3340 4558 4158 4577
rect 3340 4524 3344 4558
rect 3378 4524 3434 4558
rect 3468 4524 3524 4558
rect 3558 4524 3614 4558
rect 3648 4524 3704 4558
rect 3738 4524 3794 4558
rect 3828 4524 3884 4558
rect 3918 4524 3974 4558
rect 4008 4524 4064 4558
rect 4098 4524 4158 4558
rect 3340 4505 4158 4524
rect 4294 5372 4327 5395
rect 4361 5372 4393 5395
rect 4294 5316 4393 5372
rect 4294 5282 4327 5316
rect 4361 5282 4393 5316
rect 4294 5226 4393 5282
rect 4294 5192 4327 5226
rect 4361 5192 4393 5226
rect 4294 5136 4393 5192
rect 4294 5102 4327 5136
rect 4361 5102 4393 5136
rect 4294 5046 4393 5102
rect 4294 5012 4327 5046
rect 4361 5012 4393 5046
rect 4294 4956 4393 5012
rect 4294 4922 4327 4956
rect 4361 4922 4393 4956
rect 4294 4866 4393 4922
rect 4294 4832 4327 4866
rect 4361 4832 4393 4866
rect 4294 4776 4393 4832
rect 4294 4742 4327 4776
rect 4361 4742 4393 4776
rect 4294 4686 4393 4742
rect 4294 4652 4327 4686
rect 4361 4652 4393 4686
rect 4294 4596 4393 4652
rect 4294 4577 4327 4596
rect 4361 4577 4393 4596
rect 3105 4472 3140 4505
rect 3174 4472 3204 4505
rect 3105 4441 3204 4472
rect 4294 4472 4327 4505
rect 4361 4472 4393 4505
rect 4294 4441 4393 4472
rect 3105 4410 3268 4441
rect 3340 4410 4158 4441
rect 4230 4410 4393 4441
rect 3105 4376 3163 4410
rect 3197 4376 3253 4410
rect 3340 4376 3343 4410
rect 3377 4376 3433 4410
rect 3467 4376 3523 4410
rect 3557 4376 3613 4410
rect 3647 4376 3703 4410
rect 3737 4376 3793 4410
rect 3827 4376 3883 4410
rect 3917 4376 3973 4410
rect 4007 4376 4063 4410
rect 4097 4376 4153 4410
rect 4230 4376 4243 4410
rect 4277 4376 4393 4410
rect 3105 4342 3268 4376
rect 3340 4342 4158 4376
rect 4230 4342 4393 4376
rect 4493 5597 4656 5630
rect 4728 5597 5781 5630
rect 4493 5563 4551 5597
rect 4585 5563 4641 5597
rect 4728 5563 4731 5597
rect 4765 5563 4821 5597
rect 4855 5563 4911 5597
rect 4945 5563 5001 5597
rect 5035 5563 5091 5597
rect 5125 5563 5181 5597
rect 5215 5563 5271 5597
rect 5305 5563 5361 5597
rect 5395 5563 5451 5597
rect 5485 5563 5541 5597
rect 5575 5563 5631 5597
rect 5665 5563 5781 5597
rect 4493 5531 4656 5563
rect 4728 5531 5781 5563
rect 4493 5496 4592 5531
rect 4493 5462 4528 5496
rect 4562 5462 4592 5496
rect 5682 5496 5781 5531
rect 4493 5406 4592 5462
rect 4493 5372 4528 5406
rect 4562 5372 4592 5406
rect 4493 5316 4592 5372
rect 4493 5282 4528 5316
rect 4562 5282 4592 5316
rect 4493 5226 4592 5282
rect 4493 5192 4528 5226
rect 4562 5192 4592 5226
rect 4493 5136 4592 5192
rect 4493 5102 4528 5136
rect 4562 5102 4592 5136
rect 4493 5046 4592 5102
rect 4493 5012 4528 5046
rect 4562 5012 4592 5046
rect 4493 4956 4592 5012
rect 4493 4922 4528 4956
rect 4562 4922 4592 4956
rect 4493 4866 4592 4922
rect 4493 4832 4528 4866
rect 4562 4832 4592 4866
rect 4493 4776 4592 4832
rect 4493 4742 4528 4776
rect 4562 4742 4592 4776
rect 4493 4686 4592 4742
rect 4493 4652 4528 4686
rect 4562 4652 4592 4686
rect 4493 4596 4592 4652
rect 4493 4562 4528 4596
rect 4562 4562 4592 4596
rect 4493 4506 4592 4562
rect 4493 4472 4528 4506
rect 4562 4472 4592 4506
rect 4728 5448 5618 5467
rect 4728 5414 4751 5448
rect 4785 5414 4841 5448
rect 4875 5414 4931 5448
rect 4965 5414 5021 5448
rect 5055 5414 5111 5448
rect 5145 5414 5201 5448
rect 5235 5414 5291 5448
rect 5325 5414 5381 5448
rect 5415 5414 5471 5448
rect 5505 5414 5618 5448
rect 4728 5395 5618 5414
rect 4656 5390 4728 5395
rect 4656 5356 4675 5390
rect 4709 5356 4728 5390
rect 4656 5300 4728 5356
rect 5546 5356 5618 5395
rect 4656 5266 4675 5300
rect 4709 5266 4728 5300
rect 4656 5210 4728 5266
rect 4656 5176 4675 5210
rect 4709 5176 4728 5210
rect 4656 5120 4728 5176
rect 4656 5086 4675 5120
rect 4709 5086 4728 5120
rect 4656 5030 4728 5086
rect 4656 4996 4675 5030
rect 4709 4996 4728 5030
rect 4656 4940 4728 4996
rect 4656 4906 4675 4940
rect 4709 4906 4728 4940
rect 4656 4850 4728 4906
rect 4656 4816 4675 4850
rect 4709 4816 4728 4850
rect 4656 4760 4728 4816
rect 4656 4726 4675 4760
rect 4709 4726 4728 4760
rect 4656 4670 4728 4726
rect 4656 4636 4675 4670
rect 4709 4636 4728 4670
rect 4790 5274 5484 5333
rect 4790 5240 4849 5274
rect 4883 5246 4939 5274
rect 4911 5240 4939 5246
rect 4973 5246 5029 5274
rect 4973 5240 4977 5246
rect 4790 5212 4877 5240
rect 4911 5212 4977 5240
rect 5011 5240 5029 5246
rect 5063 5246 5119 5274
rect 5063 5240 5077 5246
rect 5011 5212 5077 5240
rect 5111 5240 5119 5246
rect 5153 5246 5209 5274
rect 5243 5246 5299 5274
rect 5333 5246 5389 5274
rect 5153 5240 5177 5246
rect 5243 5240 5277 5246
rect 5333 5240 5377 5246
rect 5423 5240 5484 5274
rect 5111 5212 5177 5240
rect 5211 5212 5277 5240
rect 5311 5212 5377 5240
rect 5411 5212 5484 5240
rect 4790 5184 5484 5212
rect 4790 5150 4849 5184
rect 4883 5150 4939 5184
rect 4973 5150 5029 5184
rect 5063 5150 5119 5184
rect 5153 5150 5209 5184
rect 5243 5150 5299 5184
rect 5333 5150 5389 5184
rect 5423 5150 5484 5184
rect 4790 5146 5484 5150
rect 4790 5112 4877 5146
rect 4911 5112 4977 5146
rect 5011 5112 5077 5146
rect 5111 5112 5177 5146
rect 5211 5112 5277 5146
rect 5311 5112 5377 5146
rect 5411 5112 5484 5146
rect 4790 5094 5484 5112
rect 4790 5060 4849 5094
rect 4883 5060 4939 5094
rect 4973 5060 5029 5094
rect 5063 5060 5119 5094
rect 5153 5060 5209 5094
rect 5243 5060 5299 5094
rect 5333 5060 5389 5094
rect 5423 5060 5484 5094
rect 4790 5046 5484 5060
rect 4790 5012 4877 5046
rect 4911 5012 4977 5046
rect 5011 5012 5077 5046
rect 5111 5012 5177 5046
rect 5211 5012 5277 5046
rect 5311 5012 5377 5046
rect 5411 5012 5484 5046
rect 4790 5004 5484 5012
rect 4790 4970 4849 5004
rect 4883 4970 4939 5004
rect 4973 4970 5029 5004
rect 5063 4970 5119 5004
rect 5153 4970 5209 5004
rect 5243 4970 5299 5004
rect 5333 4970 5389 5004
rect 5423 4970 5484 5004
rect 4790 4946 5484 4970
rect 4790 4914 4877 4946
rect 4911 4914 4977 4946
rect 4790 4880 4849 4914
rect 4911 4912 4939 4914
rect 4883 4880 4939 4912
rect 4973 4912 4977 4914
rect 5011 4914 5077 4946
rect 5011 4912 5029 4914
rect 4973 4880 5029 4912
rect 5063 4912 5077 4914
rect 5111 4914 5177 4946
rect 5211 4914 5277 4946
rect 5311 4914 5377 4946
rect 5411 4914 5484 4946
rect 5111 4912 5119 4914
rect 5063 4880 5119 4912
rect 5153 4912 5177 4914
rect 5243 4912 5277 4914
rect 5333 4912 5377 4914
rect 5153 4880 5209 4912
rect 5243 4880 5299 4912
rect 5333 4880 5389 4912
rect 5423 4880 5484 4914
rect 4790 4846 5484 4880
rect 4790 4824 4877 4846
rect 4911 4824 4977 4846
rect 4790 4790 4849 4824
rect 4911 4812 4939 4824
rect 4883 4790 4939 4812
rect 4973 4812 4977 4824
rect 5011 4824 5077 4846
rect 5011 4812 5029 4824
rect 4973 4790 5029 4812
rect 5063 4812 5077 4824
rect 5111 4824 5177 4846
rect 5211 4824 5277 4846
rect 5311 4824 5377 4846
rect 5411 4824 5484 4846
rect 5111 4812 5119 4824
rect 5063 4790 5119 4812
rect 5153 4812 5177 4824
rect 5243 4812 5277 4824
rect 5333 4812 5377 4824
rect 5153 4790 5209 4812
rect 5243 4790 5299 4812
rect 5333 4790 5389 4812
rect 5423 4790 5484 4824
rect 4790 4746 5484 4790
rect 4790 4734 4877 4746
rect 4911 4734 4977 4746
rect 4790 4700 4849 4734
rect 4911 4712 4939 4734
rect 4883 4700 4939 4712
rect 4973 4712 4977 4734
rect 5011 4734 5077 4746
rect 5011 4712 5029 4734
rect 4973 4700 5029 4712
rect 5063 4712 5077 4734
rect 5111 4734 5177 4746
rect 5211 4734 5277 4746
rect 5311 4734 5377 4746
rect 5411 4734 5484 4746
rect 5111 4712 5119 4734
rect 5063 4700 5119 4712
rect 5153 4712 5177 4734
rect 5243 4712 5277 4734
rect 5333 4712 5377 4734
rect 5153 4700 5209 4712
rect 5243 4700 5299 4712
rect 5333 4700 5389 4712
rect 5423 4700 5484 4734
rect 4790 4639 5484 4700
rect 5546 5322 5565 5356
rect 5599 5322 5618 5356
rect 5546 5266 5618 5322
rect 5546 5232 5565 5266
rect 5599 5232 5618 5266
rect 5546 5176 5618 5232
rect 5546 5142 5565 5176
rect 5599 5142 5618 5176
rect 5546 5086 5618 5142
rect 5546 5052 5565 5086
rect 5599 5052 5618 5086
rect 5546 4996 5618 5052
rect 5546 4962 5565 4996
rect 5599 4962 5618 4996
rect 5546 4906 5618 4962
rect 5546 4872 5565 4906
rect 5599 4872 5618 4906
rect 5546 4816 5618 4872
rect 5546 4782 5565 4816
rect 5599 4782 5618 4816
rect 5546 4726 5618 4782
rect 5546 4692 5565 4726
rect 5599 4692 5618 4726
rect 4656 4577 4728 4636
rect 5546 4636 5618 4692
rect 5546 4602 5565 4636
rect 5599 4602 5618 4636
rect 5546 4577 5618 4602
rect 4728 4558 5618 4577
rect 4728 4524 4732 4558
rect 4766 4524 4822 4558
rect 4856 4524 4912 4558
rect 4946 4524 5002 4558
rect 5036 4524 5092 4558
rect 5126 4524 5182 4558
rect 5216 4524 5272 4558
rect 5306 4524 5362 4558
rect 5396 4524 5452 4558
rect 5486 4524 5618 4558
rect 4728 4505 5618 4524
rect 5682 5462 5715 5496
rect 5749 5462 5781 5496
rect 5682 5406 5781 5462
rect 5682 5372 5715 5406
rect 5749 5372 5781 5406
rect 5682 5316 5781 5372
rect 5682 5282 5715 5316
rect 5749 5282 5781 5316
rect 5682 5226 5781 5282
rect 5682 5192 5715 5226
rect 5749 5192 5781 5226
rect 5682 5136 5781 5192
rect 5682 5102 5715 5136
rect 5749 5102 5781 5136
rect 5682 5046 5781 5102
rect 5682 5012 5715 5046
rect 5749 5012 5781 5046
rect 5682 4956 5781 5012
rect 5682 4922 5715 4956
rect 5749 4922 5781 4956
rect 5682 4866 5781 4922
rect 5682 4832 5715 4866
rect 5749 4832 5781 4866
rect 5682 4776 5781 4832
rect 5682 4742 5715 4776
rect 5749 4742 5781 4776
rect 5682 4686 5781 4742
rect 5682 4652 5715 4686
rect 5749 4652 5781 4686
rect 5682 4596 5781 4652
rect 5682 4562 5715 4596
rect 5749 4562 5781 4596
rect 5682 4506 5781 4562
rect 4493 4441 4592 4472
rect 5682 4472 5715 4506
rect 5749 4472 5781 4506
rect 5682 4441 5781 4472
rect 4493 4410 4656 4441
rect 4728 4410 5781 4441
rect 4493 4376 4551 4410
rect 4585 4376 4641 4410
rect 4728 4376 4731 4410
rect 4765 4376 4821 4410
rect 4855 4376 4911 4410
rect 4945 4376 5001 4410
rect 5035 4376 5091 4410
rect 5125 4376 5181 4410
rect 5215 4376 5271 4410
rect 5305 4376 5361 4410
rect 5395 4376 5451 4410
rect 5485 4376 5541 4410
rect 5575 4376 5631 4410
rect 5665 4376 5781 4410
rect 4493 4342 4656 4376
rect 4728 4342 5781 4376
rect 5881 5597 6044 5630
rect 6116 5597 7169 5630
rect 5881 5563 5939 5597
rect 5973 5563 6029 5597
rect 6116 5563 6119 5597
rect 6153 5563 6209 5597
rect 6243 5563 6299 5597
rect 6333 5563 6389 5597
rect 6423 5563 6479 5597
rect 6513 5563 6569 5597
rect 6603 5563 6659 5597
rect 6693 5563 6749 5597
rect 6783 5563 6839 5597
rect 6873 5563 6929 5597
rect 6963 5563 7019 5597
rect 7053 5563 7169 5597
rect 5881 5531 6044 5563
rect 6116 5531 7169 5563
rect 5881 5496 5980 5531
rect 5881 5462 5916 5496
rect 5950 5462 5980 5496
rect 7070 5496 7169 5531
rect 5881 5406 5980 5462
rect 5881 5372 5916 5406
rect 5950 5372 5980 5406
rect 5881 5316 5980 5372
rect 5881 5282 5916 5316
rect 5950 5282 5980 5316
rect 5881 5226 5980 5282
rect 5881 5192 5916 5226
rect 5950 5192 5980 5226
rect 5881 5136 5980 5192
rect 5881 5102 5916 5136
rect 5950 5102 5980 5136
rect 5881 5046 5980 5102
rect 5881 5012 5916 5046
rect 5950 5012 5980 5046
rect 5881 4956 5980 5012
rect 5881 4922 5916 4956
rect 5950 4922 5980 4956
rect 5881 4866 5980 4922
rect 5881 4832 5916 4866
rect 5950 4832 5980 4866
rect 5881 4776 5980 4832
rect 5881 4742 5916 4776
rect 5950 4742 5980 4776
rect 5881 4686 5980 4742
rect 5881 4652 5916 4686
rect 5950 4652 5980 4686
rect 5881 4596 5980 4652
rect 5881 4562 5916 4596
rect 5950 4562 5980 4596
rect 5881 4506 5980 4562
rect 5881 4472 5916 4506
rect 5950 4472 5980 4506
rect 6116 5448 7006 5467
rect 6116 5414 6139 5448
rect 6173 5414 6229 5448
rect 6263 5414 6319 5448
rect 6353 5414 6409 5448
rect 6443 5414 6499 5448
rect 6533 5414 6589 5448
rect 6623 5414 6679 5448
rect 6713 5414 6769 5448
rect 6803 5414 6859 5448
rect 6893 5414 7006 5448
rect 6116 5395 7006 5414
rect 6044 5390 6116 5395
rect 6044 5356 6063 5390
rect 6097 5356 6116 5390
rect 6044 5300 6116 5356
rect 6934 5356 7006 5395
rect 6044 5266 6063 5300
rect 6097 5266 6116 5300
rect 6044 5210 6116 5266
rect 6044 5176 6063 5210
rect 6097 5176 6116 5210
rect 6044 5120 6116 5176
rect 6044 5086 6063 5120
rect 6097 5086 6116 5120
rect 6044 5030 6116 5086
rect 6044 4996 6063 5030
rect 6097 4996 6116 5030
rect 6044 4940 6116 4996
rect 6044 4906 6063 4940
rect 6097 4906 6116 4940
rect 6044 4850 6116 4906
rect 6044 4816 6063 4850
rect 6097 4816 6116 4850
rect 6044 4760 6116 4816
rect 6044 4726 6063 4760
rect 6097 4726 6116 4760
rect 6044 4670 6116 4726
rect 6044 4636 6063 4670
rect 6097 4636 6116 4670
rect 6178 5274 6872 5333
rect 6178 5240 6237 5274
rect 6271 5246 6327 5274
rect 6299 5240 6327 5246
rect 6361 5246 6417 5274
rect 6361 5240 6365 5246
rect 6178 5212 6265 5240
rect 6299 5212 6365 5240
rect 6399 5240 6417 5246
rect 6451 5246 6507 5274
rect 6451 5240 6465 5246
rect 6399 5212 6465 5240
rect 6499 5240 6507 5246
rect 6541 5246 6597 5274
rect 6631 5246 6687 5274
rect 6721 5246 6777 5274
rect 6541 5240 6565 5246
rect 6631 5240 6665 5246
rect 6721 5240 6765 5246
rect 6811 5240 6872 5274
rect 6499 5212 6565 5240
rect 6599 5212 6665 5240
rect 6699 5212 6765 5240
rect 6799 5212 6872 5240
rect 6178 5184 6872 5212
rect 6178 5150 6237 5184
rect 6271 5150 6327 5184
rect 6361 5150 6417 5184
rect 6451 5150 6507 5184
rect 6541 5150 6597 5184
rect 6631 5150 6687 5184
rect 6721 5150 6777 5184
rect 6811 5150 6872 5184
rect 6178 5146 6872 5150
rect 6178 5112 6265 5146
rect 6299 5112 6365 5146
rect 6399 5112 6465 5146
rect 6499 5112 6565 5146
rect 6599 5112 6665 5146
rect 6699 5112 6765 5146
rect 6799 5112 6872 5146
rect 6178 5094 6872 5112
rect 6178 5060 6237 5094
rect 6271 5060 6327 5094
rect 6361 5060 6417 5094
rect 6451 5060 6507 5094
rect 6541 5060 6597 5094
rect 6631 5060 6687 5094
rect 6721 5060 6777 5094
rect 6811 5060 6872 5094
rect 6178 5046 6872 5060
rect 6178 5012 6265 5046
rect 6299 5012 6365 5046
rect 6399 5012 6465 5046
rect 6499 5012 6565 5046
rect 6599 5012 6665 5046
rect 6699 5012 6765 5046
rect 6799 5012 6872 5046
rect 6178 5004 6872 5012
rect 6178 4970 6237 5004
rect 6271 4970 6327 5004
rect 6361 4970 6417 5004
rect 6451 4970 6507 5004
rect 6541 4970 6597 5004
rect 6631 4970 6687 5004
rect 6721 4970 6777 5004
rect 6811 4970 6872 5004
rect 6178 4946 6872 4970
rect 6178 4914 6265 4946
rect 6299 4914 6365 4946
rect 6178 4880 6237 4914
rect 6299 4912 6327 4914
rect 6271 4880 6327 4912
rect 6361 4912 6365 4914
rect 6399 4914 6465 4946
rect 6399 4912 6417 4914
rect 6361 4880 6417 4912
rect 6451 4912 6465 4914
rect 6499 4914 6565 4946
rect 6599 4914 6665 4946
rect 6699 4914 6765 4946
rect 6799 4914 6872 4946
rect 6499 4912 6507 4914
rect 6451 4880 6507 4912
rect 6541 4912 6565 4914
rect 6631 4912 6665 4914
rect 6721 4912 6765 4914
rect 6541 4880 6597 4912
rect 6631 4880 6687 4912
rect 6721 4880 6777 4912
rect 6811 4880 6872 4914
rect 6178 4846 6872 4880
rect 6178 4824 6265 4846
rect 6299 4824 6365 4846
rect 6178 4790 6237 4824
rect 6299 4812 6327 4824
rect 6271 4790 6327 4812
rect 6361 4812 6365 4824
rect 6399 4824 6465 4846
rect 6399 4812 6417 4824
rect 6361 4790 6417 4812
rect 6451 4812 6465 4824
rect 6499 4824 6565 4846
rect 6599 4824 6665 4846
rect 6699 4824 6765 4846
rect 6799 4824 6872 4846
rect 6499 4812 6507 4824
rect 6451 4790 6507 4812
rect 6541 4812 6565 4824
rect 6631 4812 6665 4824
rect 6721 4812 6765 4824
rect 6541 4790 6597 4812
rect 6631 4790 6687 4812
rect 6721 4790 6777 4812
rect 6811 4790 6872 4824
rect 6178 4746 6872 4790
rect 6178 4734 6265 4746
rect 6299 4734 6365 4746
rect 6178 4700 6237 4734
rect 6299 4712 6327 4734
rect 6271 4700 6327 4712
rect 6361 4712 6365 4734
rect 6399 4734 6465 4746
rect 6399 4712 6417 4734
rect 6361 4700 6417 4712
rect 6451 4712 6465 4734
rect 6499 4734 6565 4746
rect 6599 4734 6665 4746
rect 6699 4734 6765 4746
rect 6799 4734 6872 4746
rect 6499 4712 6507 4734
rect 6451 4700 6507 4712
rect 6541 4712 6565 4734
rect 6631 4712 6665 4734
rect 6721 4712 6765 4734
rect 6541 4700 6597 4712
rect 6631 4700 6687 4712
rect 6721 4700 6777 4712
rect 6811 4700 6872 4734
rect 6178 4639 6872 4700
rect 6934 5322 6953 5356
rect 6987 5322 7006 5356
rect 6934 5266 7006 5322
rect 6934 5232 6953 5266
rect 6987 5232 7006 5266
rect 6934 5176 7006 5232
rect 6934 5142 6953 5176
rect 6987 5142 7006 5176
rect 6934 5086 7006 5142
rect 6934 5052 6953 5086
rect 6987 5052 7006 5086
rect 6934 4996 7006 5052
rect 6934 4962 6953 4996
rect 6987 4962 7006 4996
rect 6934 4906 7006 4962
rect 6934 4872 6953 4906
rect 6987 4872 7006 4906
rect 6934 4816 7006 4872
rect 6934 4782 6953 4816
rect 6987 4782 7006 4816
rect 6934 4726 7006 4782
rect 6934 4692 6953 4726
rect 6987 4692 7006 4726
rect 6044 4577 6116 4636
rect 6934 4636 7006 4692
rect 6934 4602 6953 4636
rect 6987 4602 7006 4636
rect 6934 4577 7006 4602
rect 6116 4558 7006 4577
rect 6116 4524 6120 4558
rect 6154 4524 6210 4558
rect 6244 4524 6300 4558
rect 6334 4524 6390 4558
rect 6424 4524 6480 4558
rect 6514 4524 6570 4558
rect 6604 4524 6660 4558
rect 6694 4524 6750 4558
rect 6784 4524 6840 4558
rect 6874 4524 7006 4558
rect 6116 4505 7006 4524
rect 7070 5462 7103 5496
rect 7137 5462 7169 5496
rect 7070 5406 7169 5462
rect 7070 5372 7103 5406
rect 7137 5372 7169 5406
rect 7070 5316 7169 5372
rect 7070 5282 7103 5316
rect 7137 5282 7169 5316
rect 7070 5226 7169 5282
rect 7070 5192 7103 5226
rect 7137 5192 7169 5226
rect 7070 5136 7169 5192
rect 7070 5102 7103 5136
rect 7137 5102 7169 5136
rect 7070 5046 7169 5102
rect 7070 5012 7103 5046
rect 7137 5012 7169 5046
rect 7070 4956 7169 5012
rect 7070 4922 7103 4956
rect 7137 4922 7169 4956
rect 7070 4866 7169 4922
rect 7070 4832 7103 4866
rect 7137 4832 7169 4866
rect 7070 4776 7169 4832
rect 7070 4742 7103 4776
rect 7137 4742 7169 4776
rect 7070 4686 7169 4742
rect 7070 4652 7103 4686
rect 7137 4652 7169 4686
rect 7070 4596 7169 4652
rect 7070 4562 7103 4596
rect 7137 4562 7169 4596
rect 7070 4506 7169 4562
rect 5881 4441 5980 4472
rect 7070 4472 7103 4506
rect 7137 4472 7169 4506
rect 7070 4441 7169 4472
rect 5881 4410 6044 4441
rect 6116 4410 7169 4441
rect 5881 4376 5939 4410
rect 5973 4376 6029 4410
rect 6116 4376 6119 4410
rect 6153 4376 6209 4410
rect 6243 4376 6299 4410
rect 6333 4376 6389 4410
rect 6423 4376 6479 4410
rect 6513 4376 6569 4410
rect 6603 4376 6659 4410
rect 6693 4376 6749 4410
rect 6783 4376 6839 4410
rect 6873 4376 6929 4410
rect 6963 4376 7019 4410
rect 7053 4376 7169 4410
rect 5881 4342 6044 4376
rect 6116 4342 7169 4376
rect 329 4209 1382 4242
rect 1454 4209 1617 4242
rect 329 4175 387 4209
rect 421 4175 477 4209
rect 511 4175 567 4209
rect 601 4175 657 4209
rect 691 4175 747 4209
rect 781 4175 837 4209
rect 871 4175 927 4209
rect 961 4175 1017 4209
rect 1051 4175 1107 4209
rect 1141 4175 1197 4209
rect 1231 4175 1287 4209
rect 1321 4175 1377 4209
rect 1454 4175 1467 4209
rect 1501 4175 1617 4209
rect 329 4143 1382 4175
rect 1454 4143 1617 4175
rect 329 4108 428 4143
rect 329 4074 364 4108
rect 398 4074 428 4108
rect 1518 4108 1617 4143
rect 329 4018 428 4074
rect 329 3984 364 4018
rect 398 3984 428 4018
rect 329 3928 428 3984
rect 329 3894 364 3928
rect 398 3894 428 3928
rect 329 3838 428 3894
rect 329 3804 364 3838
rect 398 3804 428 3838
rect 329 3748 428 3804
rect 329 3714 364 3748
rect 398 3714 428 3748
rect 329 3658 428 3714
rect 329 3624 364 3658
rect 398 3624 428 3658
rect 329 3568 428 3624
rect 329 3534 364 3568
rect 398 3534 428 3568
rect 329 3478 428 3534
rect 329 3444 364 3478
rect 398 3444 428 3478
rect 329 3388 428 3444
rect 329 3354 364 3388
rect 398 3354 428 3388
rect 329 3298 428 3354
rect 329 3264 364 3298
rect 398 3264 428 3298
rect 329 3208 428 3264
rect 329 3174 364 3208
rect 398 3174 428 3208
rect 329 3118 428 3174
rect 329 3084 364 3118
rect 398 3084 428 3118
rect 492 4060 1382 4079
rect 492 4026 587 4060
rect 621 4026 677 4060
rect 711 4026 767 4060
rect 801 4026 857 4060
rect 891 4026 947 4060
rect 981 4026 1037 4060
rect 1071 4026 1127 4060
rect 1161 4026 1217 4060
rect 1251 4026 1307 4060
rect 1341 4026 1382 4060
rect 492 4007 1382 4026
rect 492 4002 564 4007
rect 492 3968 511 4002
rect 545 3968 564 4002
rect 492 3912 564 3968
rect 1382 3968 1454 4007
rect 492 3878 511 3912
rect 545 3878 564 3912
rect 492 3822 564 3878
rect 492 3788 511 3822
rect 545 3788 564 3822
rect 492 3732 564 3788
rect 492 3698 511 3732
rect 545 3698 564 3732
rect 492 3642 564 3698
rect 492 3608 511 3642
rect 545 3608 564 3642
rect 492 3552 564 3608
rect 492 3518 511 3552
rect 545 3518 564 3552
rect 492 3462 564 3518
rect 492 3428 511 3462
rect 545 3428 564 3462
rect 492 3372 564 3428
rect 492 3338 511 3372
rect 545 3338 564 3372
rect 492 3282 564 3338
rect 492 3248 511 3282
rect 545 3248 564 3282
rect 626 3886 1320 3945
rect 626 3852 685 3886
rect 719 3858 775 3886
rect 747 3852 775 3858
rect 809 3858 865 3886
rect 809 3852 813 3858
rect 626 3824 713 3852
rect 747 3824 813 3852
rect 847 3852 865 3858
rect 899 3858 955 3886
rect 899 3852 913 3858
rect 847 3824 913 3852
rect 947 3852 955 3858
rect 989 3858 1045 3886
rect 1079 3858 1135 3886
rect 1169 3858 1225 3886
rect 989 3852 1013 3858
rect 1079 3852 1113 3858
rect 1169 3852 1213 3858
rect 1259 3852 1320 3886
rect 947 3824 1013 3852
rect 1047 3824 1113 3852
rect 1147 3824 1213 3852
rect 1247 3824 1320 3852
rect 626 3796 1320 3824
rect 626 3762 685 3796
rect 719 3762 775 3796
rect 809 3762 865 3796
rect 899 3762 955 3796
rect 989 3762 1045 3796
rect 1079 3762 1135 3796
rect 1169 3762 1225 3796
rect 1259 3762 1320 3796
rect 626 3758 1320 3762
rect 626 3724 713 3758
rect 747 3724 813 3758
rect 847 3724 913 3758
rect 947 3724 1013 3758
rect 1047 3724 1113 3758
rect 1147 3724 1213 3758
rect 1247 3724 1320 3758
rect 626 3706 1320 3724
rect 626 3672 685 3706
rect 719 3672 775 3706
rect 809 3672 865 3706
rect 899 3672 955 3706
rect 989 3672 1045 3706
rect 1079 3672 1135 3706
rect 1169 3672 1225 3706
rect 1259 3672 1320 3706
rect 626 3658 1320 3672
rect 626 3624 713 3658
rect 747 3624 813 3658
rect 847 3624 913 3658
rect 947 3624 1013 3658
rect 1047 3624 1113 3658
rect 1147 3624 1213 3658
rect 1247 3624 1320 3658
rect 626 3616 1320 3624
rect 626 3582 685 3616
rect 719 3582 775 3616
rect 809 3582 865 3616
rect 899 3582 955 3616
rect 989 3582 1045 3616
rect 1079 3582 1135 3616
rect 1169 3582 1225 3616
rect 1259 3582 1320 3616
rect 626 3558 1320 3582
rect 626 3526 713 3558
rect 747 3526 813 3558
rect 626 3492 685 3526
rect 747 3524 775 3526
rect 719 3492 775 3524
rect 809 3524 813 3526
rect 847 3526 913 3558
rect 847 3524 865 3526
rect 809 3492 865 3524
rect 899 3524 913 3526
rect 947 3526 1013 3558
rect 1047 3526 1113 3558
rect 1147 3526 1213 3558
rect 1247 3526 1320 3558
rect 947 3524 955 3526
rect 899 3492 955 3524
rect 989 3524 1013 3526
rect 1079 3524 1113 3526
rect 1169 3524 1213 3526
rect 989 3492 1045 3524
rect 1079 3492 1135 3524
rect 1169 3492 1225 3524
rect 1259 3492 1320 3526
rect 626 3458 1320 3492
rect 626 3436 713 3458
rect 747 3436 813 3458
rect 626 3402 685 3436
rect 747 3424 775 3436
rect 719 3402 775 3424
rect 809 3424 813 3436
rect 847 3436 913 3458
rect 847 3424 865 3436
rect 809 3402 865 3424
rect 899 3424 913 3436
rect 947 3436 1013 3458
rect 1047 3436 1113 3458
rect 1147 3436 1213 3458
rect 1247 3436 1320 3458
rect 947 3424 955 3436
rect 899 3402 955 3424
rect 989 3424 1013 3436
rect 1079 3424 1113 3436
rect 1169 3424 1213 3436
rect 989 3402 1045 3424
rect 1079 3402 1135 3424
rect 1169 3402 1225 3424
rect 1259 3402 1320 3436
rect 626 3358 1320 3402
rect 626 3346 713 3358
rect 747 3346 813 3358
rect 626 3312 685 3346
rect 747 3324 775 3346
rect 719 3312 775 3324
rect 809 3324 813 3346
rect 847 3346 913 3358
rect 847 3324 865 3346
rect 809 3312 865 3324
rect 899 3324 913 3346
rect 947 3346 1013 3358
rect 1047 3346 1113 3358
rect 1147 3346 1213 3358
rect 1247 3346 1320 3358
rect 947 3324 955 3346
rect 899 3312 955 3324
rect 989 3324 1013 3346
rect 1079 3324 1113 3346
rect 1169 3324 1213 3346
rect 989 3312 1045 3324
rect 1079 3312 1135 3324
rect 1169 3312 1225 3324
rect 1259 3312 1320 3346
rect 626 3251 1320 3312
rect 1382 3934 1401 3968
rect 1435 3934 1454 3968
rect 1382 3878 1454 3934
rect 1382 3844 1401 3878
rect 1435 3844 1454 3878
rect 1382 3788 1454 3844
rect 1382 3754 1401 3788
rect 1435 3754 1454 3788
rect 1382 3698 1454 3754
rect 1382 3664 1401 3698
rect 1435 3664 1454 3698
rect 1382 3608 1454 3664
rect 1382 3574 1401 3608
rect 1435 3574 1454 3608
rect 1382 3518 1454 3574
rect 1382 3484 1401 3518
rect 1435 3484 1454 3518
rect 1382 3428 1454 3484
rect 1382 3394 1401 3428
rect 1435 3394 1454 3428
rect 1382 3338 1454 3394
rect 1382 3304 1401 3338
rect 1435 3304 1454 3338
rect 492 3189 564 3248
rect 1382 3248 1454 3304
rect 1382 3214 1401 3248
rect 1435 3214 1454 3248
rect 1382 3189 1454 3214
rect 492 3170 1382 3189
rect 492 3136 568 3170
rect 602 3136 658 3170
rect 692 3136 748 3170
rect 782 3136 838 3170
rect 872 3136 928 3170
rect 962 3136 1018 3170
rect 1052 3136 1108 3170
rect 1142 3136 1198 3170
rect 1232 3136 1288 3170
rect 1322 3136 1382 3170
rect 492 3117 1382 3136
rect 1518 4074 1551 4108
rect 1585 4074 1617 4108
rect 1518 4018 1617 4074
rect 1518 3984 1551 4018
rect 1585 3984 1617 4018
rect 1518 3928 1617 3984
rect 1518 3894 1551 3928
rect 1585 3894 1617 3928
rect 1518 3838 1617 3894
rect 1518 3804 1551 3838
rect 1585 3804 1617 3838
rect 1518 3748 1617 3804
rect 1518 3714 1551 3748
rect 1585 3714 1617 3748
rect 1518 3658 1617 3714
rect 1518 3624 1551 3658
rect 1585 3624 1617 3658
rect 1518 3568 1617 3624
rect 1518 3534 1551 3568
rect 1585 3534 1617 3568
rect 1518 3478 1617 3534
rect 1518 3444 1551 3478
rect 1585 3444 1617 3478
rect 1518 3388 1617 3444
rect 1518 3354 1551 3388
rect 1585 3354 1617 3388
rect 1518 3298 1617 3354
rect 1518 3264 1551 3298
rect 1585 3264 1617 3298
rect 1518 3208 1617 3264
rect 1518 3174 1551 3208
rect 1585 3174 1617 3208
rect 1518 3118 1617 3174
rect 329 3053 428 3084
rect 1518 3084 1551 3118
rect 1585 3084 1617 3118
rect 1518 3053 1617 3084
rect 329 3022 1382 3053
rect 1454 3022 1617 3053
rect 329 2988 387 3022
rect 421 2988 477 3022
rect 511 2988 567 3022
rect 601 2988 657 3022
rect 691 2988 747 3022
rect 781 2988 837 3022
rect 871 2988 927 3022
rect 961 2988 1017 3022
rect 1051 2988 1107 3022
rect 1141 2988 1197 3022
rect 1231 2988 1287 3022
rect 1321 2988 1377 3022
rect 1454 2988 1467 3022
rect 1501 2988 1617 3022
rect 329 2954 1382 2988
rect 1454 2954 1617 2988
rect 1717 4209 2770 4242
rect 2842 4209 3005 4242
rect 1717 4175 1775 4209
rect 1809 4175 1865 4209
rect 1899 4175 1955 4209
rect 1989 4175 2045 4209
rect 2079 4175 2135 4209
rect 2169 4175 2225 4209
rect 2259 4175 2315 4209
rect 2349 4175 2405 4209
rect 2439 4175 2495 4209
rect 2529 4175 2585 4209
rect 2619 4175 2675 4209
rect 2709 4175 2765 4209
rect 2842 4175 2855 4209
rect 2889 4175 3005 4209
rect 1717 4143 2770 4175
rect 2842 4143 3005 4175
rect 1717 4108 1816 4143
rect 1717 4074 1752 4108
rect 1786 4074 1816 4108
rect 2906 4108 3005 4143
rect 2906 4079 2939 4108
rect 2973 4079 3005 4108
rect 1717 4018 1816 4074
rect 1717 3984 1752 4018
rect 1786 3984 1816 4018
rect 1717 3928 1816 3984
rect 1717 3894 1752 3928
rect 1786 3894 1816 3928
rect 1717 3838 1816 3894
rect 1717 3804 1752 3838
rect 1786 3804 1816 3838
rect 1717 3748 1816 3804
rect 1717 3714 1752 3748
rect 1786 3714 1816 3748
rect 1717 3658 1816 3714
rect 1717 3624 1752 3658
rect 1786 3624 1816 3658
rect 1717 3568 1816 3624
rect 1717 3534 1752 3568
rect 1786 3534 1816 3568
rect 1717 3478 1816 3534
rect 1717 3444 1752 3478
rect 1786 3444 1816 3478
rect 1717 3388 1816 3444
rect 1717 3354 1752 3388
rect 1786 3354 1816 3388
rect 1717 3298 1816 3354
rect 1717 3264 1752 3298
rect 1786 3264 1816 3298
rect 1717 3208 1816 3264
rect 1717 3174 1752 3208
rect 1786 3174 1816 3208
rect 1717 3118 1816 3174
rect 1717 3084 1752 3118
rect 1786 3084 1816 3118
rect 1880 4060 2770 4079
rect 1880 4026 1975 4060
rect 2009 4026 2065 4060
rect 2099 4026 2155 4060
rect 2189 4026 2245 4060
rect 2279 4026 2335 4060
rect 2369 4026 2425 4060
rect 2459 4026 2515 4060
rect 2549 4026 2605 4060
rect 2639 4026 2695 4060
rect 2729 4026 2770 4060
rect 1880 4007 2770 4026
rect 1880 4002 1952 4007
rect 1880 3968 1899 4002
rect 1933 3968 1952 4002
rect 1880 3912 1952 3968
rect 2770 3968 2842 4007
rect 1880 3878 1899 3912
rect 1933 3878 1952 3912
rect 1880 3822 1952 3878
rect 1880 3788 1899 3822
rect 1933 3788 1952 3822
rect 1880 3732 1952 3788
rect 1880 3698 1899 3732
rect 1933 3698 1952 3732
rect 1880 3642 1952 3698
rect 1880 3608 1899 3642
rect 1933 3608 1952 3642
rect 1880 3552 1952 3608
rect 1880 3518 1899 3552
rect 1933 3518 1952 3552
rect 1880 3462 1952 3518
rect 1880 3428 1899 3462
rect 1933 3428 1952 3462
rect 1880 3372 1952 3428
rect 1880 3338 1899 3372
rect 1933 3338 1952 3372
rect 1880 3282 1952 3338
rect 1880 3248 1899 3282
rect 1933 3248 1952 3282
rect 2014 3886 2708 3945
rect 2014 3852 2073 3886
rect 2107 3858 2163 3886
rect 2135 3852 2163 3858
rect 2197 3858 2253 3886
rect 2197 3852 2201 3858
rect 2014 3824 2101 3852
rect 2135 3824 2201 3852
rect 2235 3852 2253 3858
rect 2287 3858 2343 3886
rect 2287 3852 2301 3858
rect 2235 3824 2301 3852
rect 2335 3852 2343 3858
rect 2377 3858 2433 3886
rect 2467 3858 2523 3886
rect 2557 3858 2613 3886
rect 2377 3852 2401 3858
rect 2467 3852 2501 3858
rect 2557 3852 2601 3858
rect 2647 3852 2708 3886
rect 2335 3824 2401 3852
rect 2435 3824 2501 3852
rect 2535 3824 2601 3852
rect 2635 3824 2708 3852
rect 2014 3796 2708 3824
rect 2014 3762 2073 3796
rect 2107 3762 2163 3796
rect 2197 3762 2253 3796
rect 2287 3762 2343 3796
rect 2377 3762 2433 3796
rect 2467 3762 2523 3796
rect 2557 3762 2613 3796
rect 2647 3762 2708 3796
rect 2014 3758 2708 3762
rect 2014 3724 2101 3758
rect 2135 3724 2201 3758
rect 2235 3724 2301 3758
rect 2335 3724 2401 3758
rect 2435 3724 2501 3758
rect 2535 3724 2601 3758
rect 2635 3724 2708 3758
rect 2014 3706 2708 3724
rect 2014 3672 2073 3706
rect 2107 3672 2163 3706
rect 2197 3672 2253 3706
rect 2287 3672 2343 3706
rect 2377 3672 2433 3706
rect 2467 3672 2523 3706
rect 2557 3672 2613 3706
rect 2647 3672 2708 3706
rect 2014 3658 2708 3672
rect 2014 3624 2101 3658
rect 2135 3624 2201 3658
rect 2235 3624 2301 3658
rect 2335 3624 2401 3658
rect 2435 3624 2501 3658
rect 2535 3624 2601 3658
rect 2635 3624 2708 3658
rect 2014 3616 2708 3624
rect 2014 3582 2073 3616
rect 2107 3582 2163 3616
rect 2197 3582 2253 3616
rect 2287 3582 2343 3616
rect 2377 3582 2433 3616
rect 2467 3582 2523 3616
rect 2557 3582 2613 3616
rect 2647 3582 2708 3616
rect 2014 3558 2708 3582
rect 2014 3526 2101 3558
rect 2135 3526 2201 3558
rect 2014 3492 2073 3526
rect 2135 3524 2163 3526
rect 2107 3492 2163 3524
rect 2197 3524 2201 3526
rect 2235 3526 2301 3558
rect 2235 3524 2253 3526
rect 2197 3492 2253 3524
rect 2287 3524 2301 3526
rect 2335 3526 2401 3558
rect 2435 3526 2501 3558
rect 2535 3526 2601 3558
rect 2635 3526 2708 3558
rect 2335 3524 2343 3526
rect 2287 3492 2343 3524
rect 2377 3524 2401 3526
rect 2467 3524 2501 3526
rect 2557 3524 2601 3526
rect 2377 3492 2433 3524
rect 2467 3492 2523 3524
rect 2557 3492 2613 3524
rect 2647 3492 2708 3526
rect 2014 3458 2708 3492
rect 2014 3436 2101 3458
rect 2135 3436 2201 3458
rect 2014 3402 2073 3436
rect 2135 3424 2163 3436
rect 2107 3402 2163 3424
rect 2197 3424 2201 3436
rect 2235 3436 2301 3458
rect 2235 3424 2253 3436
rect 2197 3402 2253 3424
rect 2287 3424 2301 3436
rect 2335 3436 2401 3458
rect 2435 3436 2501 3458
rect 2535 3436 2601 3458
rect 2635 3436 2708 3458
rect 2335 3424 2343 3436
rect 2287 3402 2343 3424
rect 2377 3424 2401 3436
rect 2467 3424 2501 3436
rect 2557 3424 2601 3436
rect 2377 3402 2433 3424
rect 2467 3402 2523 3424
rect 2557 3402 2613 3424
rect 2647 3402 2708 3436
rect 2014 3358 2708 3402
rect 2014 3346 2101 3358
rect 2135 3346 2201 3358
rect 2014 3312 2073 3346
rect 2135 3324 2163 3346
rect 2107 3312 2163 3324
rect 2197 3324 2201 3346
rect 2235 3346 2301 3358
rect 2235 3324 2253 3346
rect 2197 3312 2253 3324
rect 2287 3324 2301 3346
rect 2335 3346 2401 3358
rect 2435 3346 2501 3358
rect 2535 3346 2601 3358
rect 2635 3346 2708 3358
rect 2335 3324 2343 3346
rect 2287 3312 2343 3324
rect 2377 3324 2401 3346
rect 2467 3324 2501 3346
rect 2557 3324 2601 3346
rect 2377 3312 2433 3324
rect 2467 3312 2523 3324
rect 2557 3312 2613 3324
rect 2647 3312 2708 3346
rect 2014 3251 2708 3312
rect 2770 3934 2789 3968
rect 2823 3934 2842 3968
rect 2770 3878 2842 3934
rect 2770 3844 2789 3878
rect 2823 3844 2842 3878
rect 2770 3788 2842 3844
rect 2770 3754 2789 3788
rect 2823 3754 2842 3788
rect 2770 3698 2842 3754
rect 2770 3664 2789 3698
rect 2823 3664 2842 3698
rect 2770 3608 2842 3664
rect 2770 3574 2789 3608
rect 2823 3574 2842 3608
rect 2770 3518 2842 3574
rect 2770 3484 2789 3518
rect 2823 3484 2842 3518
rect 2770 3428 2842 3484
rect 2770 3394 2789 3428
rect 2823 3394 2842 3428
rect 2770 3338 2842 3394
rect 2770 3304 2789 3338
rect 2823 3304 2842 3338
rect 1880 3189 1952 3248
rect 2770 3248 2842 3304
rect 2770 3214 2789 3248
rect 2823 3214 2842 3248
rect 2770 3189 2842 3214
rect 1880 3170 2842 3189
rect 1880 3136 1956 3170
rect 1990 3136 2046 3170
rect 2080 3136 2136 3170
rect 2170 3136 2226 3170
rect 2260 3136 2316 3170
rect 2350 3136 2406 3170
rect 2440 3136 2496 3170
rect 2530 3136 2586 3170
rect 2620 3136 2676 3170
rect 2710 3136 2842 3170
rect 1880 3117 2842 3136
rect 2906 3984 2939 4007
rect 2973 3984 3005 4007
rect 2906 3928 3005 3984
rect 2906 3894 2939 3928
rect 2973 3894 3005 3928
rect 2906 3838 3005 3894
rect 2906 3804 2939 3838
rect 2973 3804 3005 3838
rect 2906 3748 3005 3804
rect 2906 3714 2939 3748
rect 2973 3714 3005 3748
rect 2906 3658 3005 3714
rect 2906 3624 2939 3658
rect 2973 3624 3005 3658
rect 2906 3568 3005 3624
rect 2906 3534 2939 3568
rect 2973 3534 3005 3568
rect 2906 3478 3005 3534
rect 2906 3444 2939 3478
rect 2973 3444 3005 3478
rect 2906 3388 3005 3444
rect 2906 3354 2939 3388
rect 2973 3354 3005 3388
rect 2906 3298 3005 3354
rect 2906 3264 2939 3298
rect 2973 3264 3005 3298
rect 2906 3208 3005 3264
rect 2906 3174 2939 3208
rect 2973 3174 3005 3208
rect 2906 3118 3005 3174
rect 1717 3053 1816 3084
rect 2906 3084 2939 3118
rect 2973 3084 3005 3118
rect 2906 3053 3005 3084
rect 1717 3022 3005 3053
rect 1717 2988 1775 3022
rect 1809 2988 1865 3022
rect 1899 2988 1955 3022
rect 1989 2988 2045 3022
rect 2079 2988 2135 3022
rect 2169 2988 2225 3022
rect 2259 2988 2315 3022
rect 2349 2988 2405 3022
rect 2439 2988 2495 3022
rect 2529 2988 2585 3022
rect 2619 2988 2675 3022
rect 2709 2988 2765 3022
rect 2799 2988 2855 3022
rect 2889 2988 3005 3022
rect 1717 2954 3005 2988
rect 3105 4209 4393 4242
rect 3105 4175 3163 4209
rect 3197 4175 3253 4209
rect 3287 4175 3343 4209
rect 3377 4175 3433 4209
rect 3467 4175 3523 4209
rect 3557 4175 3613 4209
rect 3647 4175 3703 4209
rect 3737 4175 3793 4209
rect 3827 4175 3883 4209
rect 3917 4175 3973 4209
rect 4007 4175 4063 4209
rect 4097 4175 4153 4209
rect 4187 4175 4243 4209
rect 4277 4175 4393 4209
rect 3105 4143 4393 4175
rect 3105 4108 3204 4143
rect 3105 4079 3140 4108
rect 3174 4079 3204 4108
rect 4294 4108 4393 4143
rect 4294 4079 4327 4108
rect 4361 4079 4393 4108
rect 3105 3984 3140 4007
rect 3174 3984 3204 4007
rect 3105 3928 3204 3984
rect 3105 3894 3140 3928
rect 3174 3894 3204 3928
rect 3105 3838 3204 3894
rect 3105 3804 3140 3838
rect 3174 3804 3204 3838
rect 3105 3748 3204 3804
rect 3105 3714 3140 3748
rect 3174 3714 3204 3748
rect 3105 3658 3204 3714
rect 3105 3624 3140 3658
rect 3174 3624 3204 3658
rect 3105 3568 3204 3624
rect 3105 3534 3140 3568
rect 3174 3534 3204 3568
rect 3105 3478 3204 3534
rect 3105 3444 3140 3478
rect 3174 3444 3204 3478
rect 3105 3388 3204 3444
rect 3105 3354 3140 3388
rect 3174 3354 3204 3388
rect 3105 3298 3204 3354
rect 3105 3264 3140 3298
rect 3174 3264 3204 3298
rect 3105 3208 3204 3264
rect 3105 3174 3140 3208
rect 3174 3174 3204 3208
rect 3105 3118 3204 3174
rect 3105 3084 3140 3118
rect 3174 3084 3204 3118
rect 3340 4060 4158 4079
rect 3340 4026 3363 4060
rect 3397 4026 3453 4060
rect 3487 4026 3543 4060
rect 3577 4026 3633 4060
rect 3667 4026 3723 4060
rect 3757 4026 3813 4060
rect 3847 4026 3903 4060
rect 3937 4026 3993 4060
rect 4027 4026 4083 4060
rect 4117 4026 4158 4060
rect 3340 4007 4158 4026
rect 3268 4002 3340 4007
rect 3268 3968 3287 4002
rect 3321 3968 3340 4002
rect 3268 3912 3340 3968
rect 4158 3968 4230 4007
rect 3268 3878 3287 3912
rect 3321 3878 3340 3912
rect 3268 3822 3340 3878
rect 3268 3788 3287 3822
rect 3321 3788 3340 3822
rect 3268 3732 3340 3788
rect 3268 3698 3287 3732
rect 3321 3698 3340 3732
rect 3268 3642 3340 3698
rect 3268 3608 3287 3642
rect 3321 3608 3340 3642
rect 3268 3552 3340 3608
rect 3268 3518 3287 3552
rect 3321 3518 3340 3552
rect 3268 3462 3340 3518
rect 3268 3428 3287 3462
rect 3321 3428 3340 3462
rect 3268 3372 3340 3428
rect 3268 3338 3287 3372
rect 3321 3338 3340 3372
rect 3268 3282 3340 3338
rect 3268 3248 3287 3282
rect 3321 3248 3340 3282
rect 3402 3886 4096 3945
rect 3402 3852 3461 3886
rect 3495 3858 3551 3886
rect 3523 3852 3551 3858
rect 3585 3858 3641 3886
rect 3585 3852 3589 3858
rect 3402 3824 3489 3852
rect 3523 3824 3589 3852
rect 3623 3852 3641 3858
rect 3675 3858 3731 3886
rect 3675 3852 3689 3858
rect 3623 3824 3689 3852
rect 3723 3852 3731 3858
rect 3765 3858 3821 3886
rect 3855 3858 3911 3886
rect 3945 3858 4001 3886
rect 3765 3852 3789 3858
rect 3855 3852 3889 3858
rect 3945 3852 3989 3858
rect 4035 3852 4096 3886
rect 3723 3824 3789 3852
rect 3823 3824 3889 3852
rect 3923 3824 3989 3852
rect 4023 3824 4096 3852
rect 3402 3796 4096 3824
rect 3402 3762 3461 3796
rect 3495 3762 3551 3796
rect 3585 3762 3641 3796
rect 3675 3762 3731 3796
rect 3765 3762 3821 3796
rect 3855 3762 3911 3796
rect 3945 3762 4001 3796
rect 4035 3762 4096 3796
rect 3402 3758 4096 3762
rect 3402 3724 3489 3758
rect 3523 3724 3589 3758
rect 3623 3724 3689 3758
rect 3723 3724 3789 3758
rect 3823 3724 3889 3758
rect 3923 3724 3989 3758
rect 4023 3724 4096 3758
rect 3402 3706 4096 3724
rect 3402 3672 3461 3706
rect 3495 3672 3551 3706
rect 3585 3672 3641 3706
rect 3675 3672 3731 3706
rect 3765 3672 3821 3706
rect 3855 3672 3911 3706
rect 3945 3672 4001 3706
rect 4035 3672 4096 3706
rect 3402 3658 4096 3672
rect 3402 3624 3489 3658
rect 3523 3624 3589 3658
rect 3623 3624 3689 3658
rect 3723 3624 3789 3658
rect 3823 3624 3889 3658
rect 3923 3624 3989 3658
rect 4023 3624 4096 3658
rect 3402 3616 4096 3624
rect 3402 3582 3461 3616
rect 3495 3582 3551 3616
rect 3585 3582 3641 3616
rect 3675 3582 3731 3616
rect 3765 3582 3821 3616
rect 3855 3582 3911 3616
rect 3945 3582 4001 3616
rect 4035 3582 4096 3616
rect 3402 3558 4096 3582
rect 3402 3526 3489 3558
rect 3523 3526 3589 3558
rect 3402 3492 3461 3526
rect 3523 3524 3551 3526
rect 3495 3492 3551 3524
rect 3585 3524 3589 3526
rect 3623 3526 3689 3558
rect 3623 3524 3641 3526
rect 3585 3492 3641 3524
rect 3675 3524 3689 3526
rect 3723 3526 3789 3558
rect 3823 3526 3889 3558
rect 3923 3526 3989 3558
rect 4023 3526 4096 3558
rect 3723 3524 3731 3526
rect 3675 3492 3731 3524
rect 3765 3524 3789 3526
rect 3855 3524 3889 3526
rect 3945 3524 3989 3526
rect 3765 3492 3821 3524
rect 3855 3492 3911 3524
rect 3945 3492 4001 3524
rect 4035 3492 4096 3526
rect 3402 3458 4096 3492
rect 3402 3436 3489 3458
rect 3523 3436 3589 3458
rect 3402 3402 3461 3436
rect 3523 3424 3551 3436
rect 3495 3402 3551 3424
rect 3585 3424 3589 3436
rect 3623 3436 3689 3458
rect 3623 3424 3641 3436
rect 3585 3402 3641 3424
rect 3675 3424 3689 3436
rect 3723 3436 3789 3458
rect 3823 3436 3889 3458
rect 3923 3436 3989 3458
rect 4023 3436 4096 3458
rect 3723 3424 3731 3436
rect 3675 3402 3731 3424
rect 3765 3424 3789 3436
rect 3855 3424 3889 3436
rect 3945 3424 3989 3436
rect 3765 3402 3821 3424
rect 3855 3402 3911 3424
rect 3945 3402 4001 3424
rect 4035 3402 4096 3436
rect 3402 3358 4096 3402
rect 3402 3346 3489 3358
rect 3523 3346 3589 3358
rect 3402 3312 3461 3346
rect 3523 3324 3551 3346
rect 3495 3312 3551 3324
rect 3585 3324 3589 3346
rect 3623 3346 3689 3358
rect 3623 3324 3641 3346
rect 3585 3312 3641 3324
rect 3675 3324 3689 3346
rect 3723 3346 3789 3358
rect 3823 3346 3889 3358
rect 3923 3346 3989 3358
rect 4023 3346 4096 3358
rect 3723 3324 3731 3346
rect 3675 3312 3731 3324
rect 3765 3324 3789 3346
rect 3855 3324 3889 3346
rect 3945 3324 3989 3346
rect 3765 3312 3821 3324
rect 3855 3312 3911 3324
rect 3945 3312 4001 3324
rect 4035 3312 4096 3346
rect 3402 3251 4096 3312
rect 4158 3934 4177 3968
rect 4211 3934 4230 3968
rect 4158 3878 4230 3934
rect 4158 3844 4177 3878
rect 4211 3844 4230 3878
rect 4158 3788 4230 3844
rect 4158 3754 4177 3788
rect 4211 3754 4230 3788
rect 4158 3698 4230 3754
rect 4158 3664 4177 3698
rect 4211 3664 4230 3698
rect 4158 3608 4230 3664
rect 4158 3574 4177 3608
rect 4211 3574 4230 3608
rect 4158 3518 4230 3574
rect 4158 3484 4177 3518
rect 4211 3484 4230 3518
rect 4158 3428 4230 3484
rect 4158 3394 4177 3428
rect 4211 3394 4230 3428
rect 4158 3338 4230 3394
rect 4158 3304 4177 3338
rect 4211 3304 4230 3338
rect 3268 3189 3340 3248
rect 4158 3248 4230 3304
rect 4158 3214 4177 3248
rect 4211 3214 4230 3248
rect 4158 3189 4230 3214
rect 3268 3170 4230 3189
rect 3268 3136 3344 3170
rect 3378 3136 3434 3170
rect 3468 3136 3524 3170
rect 3558 3136 3614 3170
rect 3648 3136 3704 3170
rect 3738 3136 3794 3170
rect 3828 3136 3884 3170
rect 3918 3136 3974 3170
rect 4008 3136 4064 3170
rect 4098 3136 4230 3170
rect 3268 3117 4230 3136
rect 4294 3984 4327 4007
rect 4361 3984 4393 4007
rect 4294 3928 4393 3984
rect 4294 3894 4327 3928
rect 4361 3894 4393 3928
rect 4294 3838 4393 3894
rect 4294 3804 4327 3838
rect 4361 3804 4393 3838
rect 4294 3748 4393 3804
rect 4294 3714 4327 3748
rect 4361 3714 4393 3748
rect 4294 3658 4393 3714
rect 4294 3624 4327 3658
rect 4361 3624 4393 3658
rect 4294 3568 4393 3624
rect 4294 3534 4327 3568
rect 4361 3534 4393 3568
rect 4294 3478 4393 3534
rect 4294 3444 4327 3478
rect 4361 3444 4393 3478
rect 4294 3388 4393 3444
rect 4294 3354 4327 3388
rect 4361 3354 4393 3388
rect 4294 3298 4393 3354
rect 4294 3264 4327 3298
rect 4361 3264 4393 3298
rect 4294 3208 4393 3264
rect 4294 3174 4327 3208
rect 4361 3174 4393 3208
rect 4294 3118 4393 3174
rect 3105 3053 3204 3084
rect 4294 3084 4327 3118
rect 4361 3084 4393 3118
rect 4294 3053 4393 3084
rect 3105 3022 4393 3053
rect 3105 2988 3163 3022
rect 3197 2988 3253 3022
rect 3287 2988 3343 3022
rect 3377 2988 3433 3022
rect 3467 2988 3523 3022
rect 3557 2988 3613 3022
rect 3647 2988 3703 3022
rect 3737 2988 3793 3022
rect 3827 2988 3883 3022
rect 3917 2988 3973 3022
rect 4007 2988 4063 3022
rect 4097 2988 4153 3022
rect 4187 2988 4243 3022
rect 4277 2988 4393 3022
rect 3105 2954 4393 2988
rect 4493 4209 4656 4242
rect 4728 4209 5781 4242
rect 4493 4175 4551 4209
rect 4585 4175 4641 4209
rect 4728 4175 4731 4209
rect 4765 4175 4821 4209
rect 4855 4175 4911 4209
rect 4945 4175 5001 4209
rect 5035 4175 5091 4209
rect 5125 4175 5181 4209
rect 5215 4175 5271 4209
rect 5305 4175 5361 4209
rect 5395 4175 5451 4209
rect 5485 4175 5541 4209
rect 5575 4175 5631 4209
rect 5665 4175 5781 4209
rect 4493 4143 4656 4175
rect 4728 4143 5781 4175
rect 4493 4108 4592 4143
rect 4493 4079 4528 4108
rect 4562 4079 4592 4108
rect 5682 4108 5781 4143
rect 4493 3984 4528 4007
rect 4562 3984 4592 4007
rect 4493 3928 4592 3984
rect 4493 3894 4528 3928
rect 4562 3894 4592 3928
rect 4493 3838 4592 3894
rect 4493 3804 4528 3838
rect 4562 3804 4592 3838
rect 4493 3748 4592 3804
rect 4493 3714 4528 3748
rect 4562 3714 4592 3748
rect 4493 3658 4592 3714
rect 4493 3624 4528 3658
rect 4562 3624 4592 3658
rect 4493 3568 4592 3624
rect 4493 3534 4528 3568
rect 4562 3534 4592 3568
rect 4493 3478 4592 3534
rect 4493 3444 4528 3478
rect 4562 3444 4592 3478
rect 4493 3388 4592 3444
rect 4493 3354 4528 3388
rect 4562 3354 4592 3388
rect 4493 3298 4592 3354
rect 4493 3264 4528 3298
rect 4562 3264 4592 3298
rect 4493 3208 4592 3264
rect 4493 3174 4528 3208
rect 4562 3174 4592 3208
rect 4493 3118 4592 3174
rect 4493 3084 4528 3118
rect 4562 3084 4592 3118
rect 4728 4060 5618 4079
rect 4728 4026 4751 4060
rect 4785 4026 4841 4060
rect 4875 4026 4931 4060
rect 4965 4026 5021 4060
rect 5055 4026 5111 4060
rect 5145 4026 5201 4060
rect 5235 4026 5291 4060
rect 5325 4026 5381 4060
rect 5415 4026 5471 4060
rect 5505 4026 5618 4060
rect 4728 4007 5618 4026
rect 4656 4002 4728 4007
rect 4656 3968 4675 4002
rect 4709 3968 4728 4002
rect 4656 3912 4728 3968
rect 5546 3968 5618 4007
rect 4656 3878 4675 3912
rect 4709 3878 4728 3912
rect 4656 3822 4728 3878
rect 4656 3788 4675 3822
rect 4709 3788 4728 3822
rect 4656 3732 4728 3788
rect 4656 3698 4675 3732
rect 4709 3698 4728 3732
rect 4656 3642 4728 3698
rect 4656 3608 4675 3642
rect 4709 3608 4728 3642
rect 4656 3552 4728 3608
rect 4656 3518 4675 3552
rect 4709 3518 4728 3552
rect 4656 3462 4728 3518
rect 4656 3428 4675 3462
rect 4709 3428 4728 3462
rect 4656 3372 4728 3428
rect 4656 3338 4675 3372
rect 4709 3338 4728 3372
rect 4656 3282 4728 3338
rect 4656 3248 4675 3282
rect 4709 3248 4728 3282
rect 4790 3886 5484 3945
rect 4790 3852 4849 3886
rect 4883 3858 4939 3886
rect 4911 3852 4939 3858
rect 4973 3858 5029 3886
rect 4973 3852 4977 3858
rect 4790 3824 4877 3852
rect 4911 3824 4977 3852
rect 5011 3852 5029 3858
rect 5063 3858 5119 3886
rect 5063 3852 5077 3858
rect 5011 3824 5077 3852
rect 5111 3852 5119 3858
rect 5153 3858 5209 3886
rect 5243 3858 5299 3886
rect 5333 3858 5389 3886
rect 5153 3852 5177 3858
rect 5243 3852 5277 3858
rect 5333 3852 5377 3858
rect 5423 3852 5484 3886
rect 5111 3824 5177 3852
rect 5211 3824 5277 3852
rect 5311 3824 5377 3852
rect 5411 3824 5484 3852
rect 4790 3796 5484 3824
rect 4790 3762 4849 3796
rect 4883 3762 4939 3796
rect 4973 3762 5029 3796
rect 5063 3762 5119 3796
rect 5153 3762 5209 3796
rect 5243 3762 5299 3796
rect 5333 3762 5389 3796
rect 5423 3762 5484 3796
rect 4790 3758 5484 3762
rect 4790 3724 4877 3758
rect 4911 3724 4977 3758
rect 5011 3724 5077 3758
rect 5111 3724 5177 3758
rect 5211 3724 5277 3758
rect 5311 3724 5377 3758
rect 5411 3724 5484 3758
rect 4790 3706 5484 3724
rect 4790 3672 4849 3706
rect 4883 3672 4939 3706
rect 4973 3672 5029 3706
rect 5063 3672 5119 3706
rect 5153 3672 5209 3706
rect 5243 3672 5299 3706
rect 5333 3672 5389 3706
rect 5423 3672 5484 3706
rect 4790 3658 5484 3672
rect 4790 3624 4877 3658
rect 4911 3624 4977 3658
rect 5011 3624 5077 3658
rect 5111 3624 5177 3658
rect 5211 3624 5277 3658
rect 5311 3624 5377 3658
rect 5411 3624 5484 3658
rect 4790 3616 5484 3624
rect 4790 3582 4849 3616
rect 4883 3582 4939 3616
rect 4973 3582 5029 3616
rect 5063 3582 5119 3616
rect 5153 3582 5209 3616
rect 5243 3582 5299 3616
rect 5333 3582 5389 3616
rect 5423 3582 5484 3616
rect 4790 3558 5484 3582
rect 4790 3526 4877 3558
rect 4911 3526 4977 3558
rect 4790 3492 4849 3526
rect 4911 3524 4939 3526
rect 4883 3492 4939 3524
rect 4973 3524 4977 3526
rect 5011 3526 5077 3558
rect 5011 3524 5029 3526
rect 4973 3492 5029 3524
rect 5063 3524 5077 3526
rect 5111 3526 5177 3558
rect 5211 3526 5277 3558
rect 5311 3526 5377 3558
rect 5411 3526 5484 3558
rect 5111 3524 5119 3526
rect 5063 3492 5119 3524
rect 5153 3524 5177 3526
rect 5243 3524 5277 3526
rect 5333 3524 5377 3526
rect 5153 3492 5209 3524
rect 5243 3492 5299 3524
rect 5333 3492 5389 3524
rect 5423 3492 5484 3526
rect 4790 3458 5484 3492
rect 4790 3436 4877 3458
rect 4911 3436 4977 3458
rect 4790 3402 4849 3436
rect 4911 3424 4939 3436
rect 4883 3402 4939 3424
rect 4973 3424 4977 3436
rect 5011 3436 5077 3458
rect 5011 3424 5029 3436
rect 4973 3402 5029 3424
rect 5063 3424 5077 3436
rect 5111 3436 5177 3458
rect 5211 3436 5277 3458
rect 5311 3436 5377 3458
rect 5411 3436 5484 3458
rect 5111 3424 5119 3436
rect 5063 3402 5119 3424
rect 5153 3424 5177 3436
rect 5243 3424 5277 3436
rect 5333 3424 5377 3436
rect 5153 3402 5209 3424
rect 5243 3402 5299 3424
rect 5333 3402 5389 3424
rect 5423 3402 5484 3436
rect 4790 3358 5484 3402
rect 4790 3346 4877 3358
rect 4911 3346 4977 3358
rect 4790 3312 4849 3346
rect 4911 3324 4939 3346
rect 4883 3312 4939 3324
rect 4973 3324 4977 3346
rect 5011 3346 5077 3358
rect 5011 3324 5029 3346
rect 4973 3312 5029 3324
rect 5063 3324 5077 3346
rect 5111 3346 5177 3358
rect 5211 3346 5277 3358
rect 5311 3346 5377 3358
rect 5411 3346 5484 3358
rect 5111 3324 5119 3346
rect 5063 3312 5119 3324
rect 5153 3324 5177 3346
rect 5243 3324 5277 3346
rect 5333 3324 5377 3346
rect 5153 3312 5209 3324
rect 5243 3312 5299 3324
rect 5333 3312 5389 3324
rect 5423 3312 5484 3346
rect 4790 3251 5484 3312
rect 5546 3934 5565 3968
rect 5599 3934 5618 3968
rect 5546 3878 5618 3934
rect 5546 3844 5565 3878
rect 5599 3844 5618 3878
rect 5546 3788 5618 3844
rect 5546 3754 5565 3788
rect 5599 3754 5618 3788
rect 5546 3698 5618 3754
rect 5546 3664 5565 3698
rect 5599 3664 5618 3698
rect 5546 3608 5618 3664
rect 5546 3574 5565 3608
rect 5599 3574 5618 3608
rect 5546 3518 5618 3574
rect 5546 3484 5565 3518
rect 5599 3484 5618 3518
rect 5546 3428 5618 3484
rect 5546 3394 5565 3428
rect 5599 3394 5618 3428
rect 5546 3338 5618 3394
rect 5546 3304 5565 3338
rect 5599 3304 5618 3338
rect 4656 3189 4728 3248
rect 5546 3248 5618 3304
rect 5546 3214 5565 3248
rect 5599 3214 5618 3248
rect 5546 3189 5618 3214
rect 4656 3170 5618 3189
rect 4656 3136 4732 3170
rect 4766 3136 4822 3170
rect 4856 3136 4912 3170
rect 4946 3136 5002 3170
rect 5036 3136 5092 3170
rect 5126 3136 5182 3170
rect 5216 3136 5272 3170
rect 5306 3136 5362 3170
rect 5396 3136 5452 3170
rect 5486 3136 5618 3170
rect 4656 3117 5618 3136
rect 5682 4074 5715 4108
rect 5749 4074 5781 4108
rect 5682 4018 5781 4074
rect 5682 3984 5715 4018
rect 5749 3984 5781 4018
rect 5682 3928 5781 3984
rect 5682 3894 5715 3928
rect 5749 3894 5781 3928
rect 5682 3838 5781 3894
rect 5682 3804 5715 3838
rect 5749 3804 5781 3838
rect 5682 3748 5781 3804
rect 5682 3714 5715 3748
rect 5749 3714 5781 3748
rect 5682 3658 5781 3714
rect 5682 3624 5715 3658
rect 5749 3624 5781 3658
rect 5682 3568 5781 3624
rect 5682 3534 5715 3568
rect 5749 3534 5781 3568
rect 5682 3478 5781 3534
rect 5682 3444 5715 3478
rect 5749 3444 5781 3478
rect 5682 3388 5781 3444
rect 5682 3354 5715 3388
rect 5749 3354 5781 3388
rect 5682 3298 5781 3354
rect 5682 3264 5715 3298
rect 5749 3264 5781 3298
rect 5682 3208 5781 3264
rect 5682 3174 5715 3208
rect 5749 3174 5781 3208
rect 5682 3118 5781 3174
rect 4493 3053 4592 3084
rect 5682 3084 5715 3118
rect 5749 3084 5781 3118
rect 5682 3053 5781 3084
rect 4493 3022 5781 3053
rect 4493 2988 4551 3022
rect 4585 2988 4641 3022
rect 4675 2988 4731 3022
rect 4765 2988 4821 3022
rect 4855 2988 4911 3022
rect 4945 2988 5001 3022
rect 5035 2988 5091 3022
rect 5125 2988 5181 3022
rect 5215 2988 5271 3022
rect 5305 2988 5361 3022
rect 5395 2988 5451 3022
rect 5485 2988 5541 3022
rect 5575 2988 5631 3022
rect 5665 2988 5781 3022
rect 4493 2954 5781 2988
rect 5881 4209 6044 4242
rect 6116 4209 7169 4242
rect 5881 4175 5939 4209
rect 5973 4175 6029 4209
rect 6116 4175 6119 4209
rect 6153 4175 6209 4209
rect 6243 4175 6299 4209
rect 6333 4175 6389 4209
rect 6423 4175 6479 4209
rect 6513 4175 6569 4209
rect 6603 4175 6659 4209
rect 6693 4175 6749 4209
rect 6783 4175 6839 4209
rect 6873 4175 6929 4209
rect 6963 4175 7019 4209
rect 7053 4175 7169 4209
rect 5881 4143 6044 4175
rect 6116 4143 7169 4175
rect 5881 4108 5980 4143
rect 5881 4074 5916 4108
rect 5950 4074 5980 4108
rect 7070 4108 7169 4143
rect 5881 4018 5980 4074
rect 5881 3984 5916 4018
rect 5950 3984 5980 4018
rect 5881 3928 5980 3984
rect 5881 3894 5916 3928
rect 5950 3894 5980 3928
rect 5881 3838 5980 3894
rect 5881 3804 5916 3838
rect 5950 3804 5980 3838
rect 5881 3748 5980 3804
rect 5881 3714 5916 3748
rect 5950 3714 5980 3748
rect 5881 3658 5980 3714
rect 5881 3624 5916 3658
rect 5950 3624 5980 3658
rect 5881 3568 5980 3624
rect 5881 3534 5916 3568
rect 5950 3534 5980 3568
rect 5881 3478 5980 3534
rect 5881 3444 5916 3478
rect 5950 3444 5980 3478
rect 5881 3388 5980 3444
rect 5881 3354 5916 3388
rect 5950 3354 5980 3388
rect 5881 3298 5980 3354
rect 5881 3264 5916 3298
rect 5950 3264 5980 3298
rect 5881 3208 5980 3264
rect 5881 3174 5916 3208
rect 5950 3174 5980 3208
rect 5881 3118 5980 3174
rect 5881 3084 5916 3118
rect 5950 3084 5980 3118
rect 6116 4060 7006 4079
rect 6116 4026 6139 4060
rect 6173 4026 6229 4060
rect 6263 4026 6319 4060
rect 6353 4026 6409 4060
rect 6443 4026 6499 4060
rect 6533 4026 6589 4060
rect 6623 4026 6679 4060
rect 6713 4026 6769 4060
rect 6803 4026 6859 4060
rect 6893 4026 7006 4060
rect 6116 4007 7006 4026
rect 6044 4002 6116 4007
rect 6044 3968 6063 4002
rect 6097 3968 6116 4002
rect 6044 3912 6116 3968
rect 6934 3968 7006 4007
rect 6044 3878 6063 3912
rect 6097 3878 6116 3912
rect 6044 3822 6116 3878
rect 6044 3788 6063 3822
rect 6097 3788 6116 3822
rect 6044 3732 6116 3788
rect 6044 3698 6063 3732
rect 6097 3698 6116 3732
rect 6044 3642 6116 3698
rect 6044 3608 6063 3642
rect 6097 3608 6116 3642
rect 6044 3552 6116 3608
rect 6044 3518 6063 3552
rect 6097 3518 6116 3552
rect 6044 3462 6116 3518
rect 6044 3428 6063 3462
rect 6097 3428 6116 3462
rect 6044 3372 6116 3428
rect 6044 3338 6063 3372
rect 6097 3338 6116 3372
rect 6044 3282 6116 3338
rect 6044 3248 6063 3282
rect 6097 3248 6116 3282
rect 6178 3886 6872 3945
rect 6178 3852 6237 3886
rect 6271 3858 6327 3886
rect 6299 3852 6327 3858
rect 6361 3858 6417 3886
rect 6361 3852 6365 3858
rect 6178 3824 6265 3852
rect 6299 3824 6365 3852
rect 6399 3852 6417 3858
rect 6451 3858 6507 3886
rect 6451 3852 6465 3858
rect 6399 3824 6465 3852
rect 6499 3852 6507 3858
rect 6541 3858 6597 3886
rect 6631 3858 6687 3886
rect 6721 3858 6777 3886
rect 6541 3852 6565 3858
rect 6631 3852 6665 3858
rect 6721 3852 6765 3858
rect 6811 3852 6872 3886
rect 6499 3824 6565 3852
rect 6599 3824 6665 3852
rect 6699 3824 6765 3852
rect 6799 3824 6872 3852
rect 6178 3796 6872 3824
rect 6178 3762 6237 3796
rect 6271 3762 6327 3796
rect 6361 3762 6417 3796
rect 6451 3762 6507 3796
rect 6541 3762 6597 3796
rect 6631 3762 6687 3796
rect 6721 3762 6777 3796
rect 6811 3762 6872 3796
rect 6178 3758 6872 3762
rect 6178 3724 6265 3758
rect 6299 3724 6365 3758
rect 6399 3724 6465 3758
rect 6499 3724 6565 3758
rect 6599 3724 6665 3758
rect 6699 3724 6765 3758
rect 6799 3724 6872 3758
rect 6178 3706 6872 3724
rect 6178 3672 6237 3706
rect 6271 3672 6327 3706
rect 6361 3672 6417 3706
rect 6451 3672 6507 3706
rect 6541 3672 6597 3706
rect 6631 3672 6687 3706
rect 6721 3672 6777 3706
rect 6811 3672 6872 3706
rect 6178 3658 6872 3672
rect 6178 3624 6265 3658
rect 6299 3624 6365 3658
rect 6399 3624 6465 3658
rect 6499 3624 6565 3658
rect 6599 3624 6665 3658
rect 6699 3624 6765 3658
rect 6799 3624 6872 3658
rect 6178 3616 6872 3624
rect 6178 3582 6237 3616
rect 6271 3582 6327 3616
rect 6361 3582 6417 3616
rect 6451 3582 6507 3616
rect 6541 3582 6597 3616
rect 6631 3582 6687 3616
rect 6721 3582 6777 3616
rect 6811 3582 6872 3616
rect 6178 3558 6872 3582
rect 6178 3526 6265 3558
rect 6299 3526 6365 3558
rect 6178 3492 6237 3526
rect 6299 3524 6327 3526
rect 6271 3492 6327 3524
rect 6361 3524 6365 3526
rect 6399 3526 6465 3558
rect 6399 3524 6417 3526
rect 6361 3492 6417 3524
rect 6451 3524 6465 3526
rect 6499 3526 6565 3558
rect 6599 3526 6665 3558
rect 6699 3526 6765 3558
rect 6799 3526 6872 3558
rect 6499 3524 6507 3526
rect 6451 3492 6507 3524
rect 6541 3524 6565 3526
rect 6631 3524 6665 3526
rect 6721 3524 6765 3526
rect 6541 3492 6597 3524
rect 6631 3492 6687 3524
rect 6721 3492 6777 3524
rect 6811 3492 6872 3526
rect 6178 3458 6872 3492
rect 6178 3436 6265 3458
rect 6299 3436 6365 3458
rect 6178 3402 6237 3436
rect 6299 3424 6327 3436
rect 6271 3402 6327 3424
rect 6361 3424 6365 3436
rect 6399 3436 6465 3458
rect 6399 3424 6417 3436
rect 6361 3402 6417 3424
rect 6451 3424 6465 3436
rect 6499 3436 6565 3458
rect 6599 3436 6665 3458
rect 6699 3436 6765 3458
rect 6799 3436 6872 3458
rect 6499 3424 6507 3436
rect 6451 3402 6507 3424
rect 6541 3424 6565 3436
rect 6631 3424 6665 3436
rect 6721 3424 6765 3436
rect 6541 3402 6597 3424
rect 6631 3402 6687 3424
rect 6721 3402 6777 3424
rect 6811 3402 6872 3436
rect 6178 3358 6872 3402
rect 6178 3346 6265 3358
rect 6299 3346 6365 3358
rect 6178 3312 6237 3346
rect 6299 3324 6327 3346
rect 6271 3312 6327 3324
rect 6361 3324 6365 3346
rect 6399 3346 6465 3358
rect 6399 3324 6417 3346
rect 6361 3312 6417 3324
rect 6451 3324 6465 3346
rect 6499 3346 6565 3358
rect 6599 3346 6665 3358
rect 6699 3346 6765 3358
rect 6799 3346 6872 3358
rect 6499 3324 6507 3346
rect 6451 3312 6507 3324
rect 6541 3324 6565 3346
rect 6631 3324 6665 3346
rect 6721 3324 6765 3346
rect 6541 3312 6597 3324
rect 6631 3312 6687 3324
rect 6721 3312 6777 3324
rect 6811 3312 6872 3346
rect 6178 3251 6872 3312
rect 6934 3934 6953 3968
rect 6987 3934 7006 3968
rect 6934 3878 7006 3934
rect 6934 3844 6953 3878
rect 6987 3844 7006 3878
rect 6934 3788 7006 3844
rect 6934 3754 6953 3788
rect 6987 3754 7006 3788
rect 6934 3698 7006 3754
rect 6934 3664 6953 3698
rect 6987 3664 7006 3698
rect 6934 3608 7006 3664
rect 6934 3574 6953 3608
rect 6987 3574 7006 3608
rect 6934 3518 7006 3574
rect 6934 3484 6953 3518
rect 6987 3484 7006 3518
rect 6934 3428 7006 3484
rect 6934 3394 6953 3428
rect 6987 3394 7006 3428
rect 6934 3338 7006 3394
rect 6934 3304 6953 3338
rect 6987 3304 7006 3338
rect 6044 3189 6116 3248
rect 6934 3248 7006 3304
rect 6934 3214 6953 3248
rect 6987 3214 7006 3248
rect 6934 3189 7006 3214
rect 6116 3170 7006 3189
rect 6116 3136 6120 3170
rect 6154 3136 6210 3170
rect 6244 3136 6300 3170
rect 6334 3136 6390 3170
rect 6424 3136 6480 3170
rect 6514 3136 6570 3170
rect 6604 3136 6660 3170
rect 6694 3136 6750 3170
rect 6784 3136 6840 3170
rect 6874 3136 7006 3170
rect 6116 3117 7006 3136
rect 7070 4074 7103 4108
rect 7137 4074 7169 4108
rect 7070 4018 7169 4074
rect 7070 3984 7103 4018
rect 7137 3984 7169 4018
rect 7070 3928 7169 3984
rect 7070 3894 7103 3928
rect 7137 3894 7169 3928
rect 7070 3838 7169 3894
rect 7070 3804 7103 3838
rect 7137 3804 7169 3838
rect 7070 3748 7169 3804
rect 7070 3714 7103 3748
rect 7137 3714 7169 3748
rect 7070 3658 7169 3714
rect 7070 3624 7103 3658
rect 7137 3624 7169 3658
rect 7070 3568 7169 3624
rect 7070 3534 7103 3568
rect 7137 3534 7169 3568
rect 7070 3478 7169 3534
rect 7070 3444 7103 3478
rect 7137 3444 7169 3478
rect 7070 3388 7169 3444
rect 7070 3354 7103 3388
rect 7137 3354 7169 3388
rect 7070 3298 7169 3354
rect 7070 3264 7103 3298
rect 7137 3264 7169 3298
rect 7070 3208 7169 3264
rect 7070 3174 7103 3208
rect 7137 3174 7169 3208
rect 7070 3118 7169 3174
rect 5881 3053 5980 3084
rect 7070 3084 7103 3118
rect 7137 3084 7169 3118
rect 7070 3053 7169 3084
rect 5881 3022 6044 3053
rect 6116 3022 7169 3053
rect 5881 2988 5939 3022
rect 5973 2988 6029 3022
rect 6116 2988 6119 3022
rect 6153 2988 6209 3022
rect 6243 2988 6299 3022
rect 6333 2988 6389 3022
rect 6423 2988 6479 3022
rect 6513 2988 6569 3022
rect 6603 2988 6659 3022
rect 6693 2988 6749 3022
rect 6783 2988 6839 3022
rect 6873 2988 6929 3022
rect 6963 2988 7019 3022
rect 7053 2988 7169 3022
rect 5881 2954 6044 2988
rect 6116 2954 7169 2988
rect 329 2821 1382 2854
rect 1454 2821 1617 2854
rect 329 2787 387 2821
rect 421 2787 477 2821
rect 511 2787 567 2821
rect 601 2787 657 2821
rect 691 2787 747 2821
rect 781 2787 837 2821
rect 871 2787 927 2821
rect 961 2787 1017 2821
rect 1051 2787 1107 2821
rect 1141 2787 1197 2821
rect 1231 2787 1287 2821
rect 1321 2787 1377 2821
rect 1454 2787 1467 2821
rect 1501 2787 1617 2821
rect 329 2755 1382 2787
rect 1454 2755 1617 2787
rect 329 2720 428 2755
rect 329 2686 364 2720
rect 398 2686 428 2720
rect 1518 2720 1617 2755
rect 1518 2691 1551 2720
rect 1585 2691 1617 2720
rect 329 2630 428 2686
rect 329 2596 364 2630
rect 398 2596 428 2630
rect 329 2540 428 2596
rect 329 2506 364 2540
rect 398 2506 428 2540
rect 329 2450 428 2506
rect 329 2416 364 2450
rect 398 2416 428 2450
rect 329 2360 428 2416
rect 329 2326 364 2360
rect 398 2326 428 2360
rect 329 2270 428 2326
rect 329 2236 364 2270
rect 398 2236 428 2270
rect 329 2180 428 2236
rect 329 2146 364 2180
rect 398 2146 428 2180
rect 329 2090 428 2146
rect 329 2056 364 2090
rect 398 2056 428 2090
rect 329 2000 428 2056
rect 329 1966 364 2000
rect 398 1966 428 2000
rect 329 1910 428 1966
rect 329 1876 364 1910
rect 398 1876 428 1910
rect 329 1820 428 1876
rect 329 1786 364 1820
rect 398 1786 428 1820
rect 329 1730 428 1786
rect 329 1696 364 1730
rect 398 1696 428 1730
rect 492 2672 1382 2691
rect 492 2638 587 2672
rect 621 2638 677 2672
rect 711 2638 767 2672
rect 801 2638 857 2672
rect 891 2638 947 2672
rect 981 2638 1037 2672
rect 1071 2638 1127 2672
rect 1161 2638 1217 2672
rect 1251 2638 1307 2672
rect 1341 2638 1382 2672
rect 492 2619 1382 2638
rect 492 2614 564 2619
rect 492 2580 511 2614
rect 545 2580 564 2614
rect 492 2524 564 2580
rect 1382 2580 1454 2619
rect 492 2490 511 2524
rect 545 2490 564 2524
rect 492 2434 564 2490
rect 492 2400 511 2434
rect 545 2400 564 2434
rect 492 2344 564 2400
rect 492 2310 511 2344
rect 545 2310 564 2344
rect 492 2254 564 2310
rect 492 2220 511 2254
rect 545 2220 564 2254
rect 492 2164 564 2220
rect 492 2130 511 2164
rect 545 2130 564 2164
rect 492 2074 564 2130
rect 492 2040 511 2074
rect 545 2040 564 2074
rect 492 1984 564 2040
rect 492 1950 511 1984
rect 545 1950 564 1984
rect 492 1894 564 1950
rect 492 1860 511 1894
rect 545 1860 564 1894
rect 626 2498 1320 2557
rect 626 2464 685 2498
rect 719 2470 775 2498
rect 747 2464 775 2470
rect 809 2470 865 2498
rect 809 2464 813 2470
rect 626 2436 713 2464
rect 747 2436 813 2464
rect 847 2464 865 2470
rect 899 2470 955 2498
rect 899 2464 913 2470
rect 847 2436 913 2464
rect 947 2464 955 2470
rect 989 2470 1045 2498
rect 1079 2470 1135 2498
rect 1169 2470 1225 2498
rect 989 2464 1013 2470
rect 1079 2464 1113 2470
rect 1169 2464 1213 2470
rect 1259 2464 1320 2498
rect 947 2436 1013 2464
rect 1047 2436 1113 2464
rect 1147 2436 1213 2464
rect 1247 2436 1320 2464
rect 626 2408 1320 2436
rect 626 2374 685 2408
rect 719 2374 775 2408
rect 809 2374 865 2408
rect 899 2374 955 2408
rect 989 2374 1045 2408
rect 1079 2374 1135 2408
rect 1169 2374 1225 2408
rect 1259 2374 1320 2408
rect 626 2370 1320 2374
rect 626 2336 713 2370
rect 747 2336 813 2370
rect 847 2336 913 2370
rect 947 2336 1013 2370
rect 1047 2336 1113 2370
rect 1147 2336 1213 2370
rect 1247 2336 1320 2370
rect 626 2318 1320 2336
rect 626 2284 685 2318
rect 719 2284 775 2318
rect 809 2284 865 2318
rect 899 2284 955 2318
rect 989 2284 1045 2318
rect 1079 2284 1135 2318
rect 1169 2284 1225 2318
rect 1259 2284 1320 2318
rect 626 2270 1320 2284
rect 626 2236 713 2270
rect 747 2236 813 2270
rect 847 2236 913 2270
rect 947 2236 1013 2270
rect 1047 2236 1113 2270
rect 1147 2236 1213 2270
rect 1247 2236 1320 2270
rect 626 2228 1320 2236
rect 626 2194 685 2228
rect 719 2194 775 2228
rect 809 2194 865 2228
rect 899 2194 955 2228
rect 989 2194 1045 2228
rect 1079 2194 1135 2228
rect 1169 2194 1225 2228
rect 1259 2194 1320 2228
rect 626 2170 1320 2194
rect 626 2138 713 2170
rect 747 2138 813 2170
rect 626 2104 685 2138
rect 747 2136 775 2138
rect 719 2104 775 2136
rect 809 2136 813 2138
rect 847 2138 913 2170
rect 847 2136 865 2138
rect 809 2104 865 2136
rect 899 2136 913 2138
rect 947 2138 1013 2170
rect 1047 2138 1113 2170
rect 1147 2138 1213 2170
rect 1247 2138 1320 2170
rect 947 2136 955 2138
rect 899 2104 955 2136
rect 989 2136 1013 2138
rect 1079 2136 1113 2138
rect 1169 2136 1213 2138
rect 989 2104 1045 2136
rect 1079 2104 1135 2136
rect 1169 2104 1225 2136
rect 1259 2104 1320 2138
rect 626 2070 1320 2104
rect 626 2048 713 2070
rect 747 2048 813 2070
rect 626 2014 685 2048
rect 747 2036 775 2048
rect 719 2014 775 2036
rect 809 2036 813 2048
rect 847 2048 913 2070
rect 847 2036 865 2048
rect 809 2014 865 2036
rect 899 2036 913 2048
rect 947 2048 1013 2070
rect 1047 2048 1113 2070
rect 1147 2048 1213 2070
rect 1247 2048 1320 2070
rect 947 2036 955 2048
rect 899 2014 955 2036
rect 989 2036 1013 2048
rect 1079 2036 1113 2048
rect 1169 2036 1213 2048
rect 989 2014 1045 2036
rect 1079 2014 1135 2036
rect 1169 2014 1225 2036
rect 1259 2014 1320 2048
rect 626 1970 1320 2014
rect 626 1958 713 1970
rect 747 1958 813 1970
rect 626 1924 685 1958
rect 747 1936 775 1958
rect 719 1924 775 1936
rect 809 1936 813 1958
rect 847 1958 913 1970
rect 847 1936 865 1958
rect 809 1924 865 1936
rect 899 1936 913 1958
rect 947 1958 1013 1970
rect 1047 1958 1113 1970
rect 1147 1958 1213 1970
rect 1247 1958 1320 1970
rect 947 1936 955 1958
rect 899 1924 955 1936
rect 989 1936 1013 1958
rect 1079 1936 1113 1958
rect 1169 1936 1213 1958
rect 989 1924 1045 1936
rect 1079 1924 1135 1936
rect 1169 1924 1225 1936
rect 1259 1924 1320 1958
rect 626 1863 1320 1924
rect 1382 2546 1401 2580
rect 1435 2546 1454 2580
rect 1382 2490 1454 2546
rect 1382 2456 1401 2490
rect 1435 2456 1454 2490
rect 1382 2400 1454 2456
rect 1382 2366 1401 2400
rect 1435 2366 1454 2400
rect 1382 2310 1454 2366
rect 1382 2276 1401 2310
rect 1435 2276 1454 2310
rect 1382 2220 1454 2276
rect 1382 2186 1401 2220
rect 1435 2186 1454 2220
rect 1382 2130 1454 2186
rect 1382 2096 1401 2130
rect 1435 2096 1454 2130
rect 1382 2040 1454 2096
rect 1382 2006 1401 2040
rect 1435 2006 1454 2040
rect 1382 1950 1454 2006
rect 1382 1916 1401 1950
rect 1435 1916 1454 1950
rect 492 1801 564 1860
rect 1382 1860 1454 1916
rect 1382 1826 1401 1860
rect 1435 1826 1454 1860
rect 1382 1801 1454 1826
rect 492 1782 1454 1801
rect 492 1748 568 1782
rect 602 1748 658 1782
rect 692 1748 748 1782
rect 782 1748 838 1782
rect 872 1748 928 1782
rect 962 1748 1018 1782
rect 1052 1748 1108 1782
rect 1142 1748 1198 1782
rect 1232 1748 1288 1782
rect 1322 1748 1454 1782
rect 492 1729 1454 1748
rect 1518 2596 1551 2619
rect 1585 2596 1617 2619
rect 1518 2540 1617 2596
rect 1518 2506 1551 2540
rect 1585 2506 1617 2540
rect 1518 2450 1617 2506
rect 1518 2416 1551 2450
rect 1585 2416 1617 2450
rect 1518 2360 1617 2416
rect 1518 2326 1551 2360
rect 1585 2326 1617 2360
rect 1518 2270 1617 2326
rect 1518 2236 1551 2270
rect 1585 2236 1617 2270
rect 1518 2180 1617 2236
rect 1518 2146 1551 2180
rect 1585 2146 1617 2180
rect 1518 2090 1617 2146
rect 1518 2056 1551 2090
rect 1585 2056 1617 2090
rect 1518 2000 1617 2056
rect 1518 1966 1551 2000
rect 1585 1966 1617 2000
rect 1518 1910 1617 1966
rect 1518 1876 1551 1910
rect 1585 1876 1617 1910
rect 1518 1820 1617 1876
rect 1518 1786 1551 1820
rect 1585 1786 1617 1820
rect 1518 1730 1617 1786
rect 329 1665 428 1696
rect 1518 1696 1551 1730
rect 1585 1696 1617 1730
rect 1518 1665 1617 1696
rect 329 1634 1617 1665
rect 329 1600 387 1634
rect 421 1600 477 1634
rect 511 1600 567 1634
rect 601 1600 657 1634
rect 691 1600 747 1634
rect 781 1600 837 1634
rect 871 1600 927 1634
rect 961 1600 1017 1634
rect 1051 1600 1107 1634
rect 1141 1600 1197 1634
rect 1231 1600 1287 1634
rect 1321 1600 1377 1634
rect 1411 1600 1467 1634
rect 1501 1600 1617 1634
rect 329 1566 1617 1600
rect 1717 2821 3005 2854
rect 1717 2787 1775 2821
rect 1809 2787 1865 2821
rect 1899 2787 1955 2821
rect 1989 2787 2045 2821
rect 2079 2787 2135 2821
rect 2169 2787 2225 2821
rect 2259 2787 2315 2821
rect 2349 2787 2405 2821
rect 2439 2787 2495 2821
rect 2529 2787 2585 2821
rect 2619 2787 2675 2821
rect 2709 2787 2765 2821
rect 2799 2787 2855 2821
rect 2889 2787 3005 2821
rect 1717 2755 3005 2787
rect 1717 2720 1816 2755
rect 1717 2691 1752 2720
rect 1786 2691 1816 2720
rect 2906 2720 3005 2755
rect 2906 2691 2939 2720
rect 2973 2691 3005 2720
rect 1717 2596 1752 2619
rect 1786 2596 1816 2619
rect 1717 2540 1816 2596
rect 1717 2506 1752 2540
rect 1786 2506 1816 2540
rect 1717 2450 1816 2506
rect 1717 2416 1752 2450
rect 1786 2416 1816 2450
rect 1717 2360 1816 2416
rect 1717 2326 1752 2360
rect 1786 2326 1816 2360
rect 1717 2270 1816 2326
rect 1717 2236 1752 2270
rect 1786 2236 1816 2270
rect 1717 2180 1816 2236
rect 1717 2146 1752 2180
rect 1786 2146 1816 2180
rect 1717 2090 1816 2146
rect 1717 2056 1752 2090
rect 1786 2056 1816 2090
rect 1717 2000 1816 2056
rect 1717 1966 1752 2000
rect 1786 1966 1816 2000
rect 1717 1910 1816 1966
rect 1717 1876 1752 1910
rect 1786 1876 1816 1910
rect 1717 1820 1816 1876
rect 1717 1786 1752 1820
rect 1786 1786 1816 1820
rect 1717 1730 1816 1786
rect 1717 1696 1752 1730
rect 1786 1696 1816 1730
rect 1952 2672 2770 2691
rect 1952 2638 1975 2672
rect 2009 2638 2065 2672
rect 2099 2638 2155 2672
rect 2189 2638 2245 2672
rect 2279 2638 2335 2672
rect 2369 2638 2425 2672
rect 2459 2638 2515 2672
rect 2549 2638 2605 2672
rect 2639 2638 2695 2672
rect 2729 2638 2770 2672
rect 1952 2619 2770 2638
rect 1880 2614 1952 2619
rect 1880 2580 1899 2614
rect 1933 2580 1952 2614
rect 1880 2524 1952 2580
rect 2770 2580 2842 2619
rect 1880 2490 1899 2524
rect 1933 2490 1952 2524
rect 1880 2434 1952 2490
rect 1880 2400 1899 2434
rect 1933 2400 1952 2434
rect 1880 2344 1952 2400
rect 1880 2310 1899 2344
rect 1933 2310 1952 2344
rect 1880 2254 1952 2310
rect 1880 2220 1899 2254
rect 1933 2220 1952 2254
rect 1880 2164 1952 2220
rect 1880 2130 1899 2164
rect 1933 2130 1952 2164
rect 1880 2074 1952 2130
rect 1880 2040 1899 2074
rect 1933 2040 1952 2074
rect 1880 1984 1952 2040
rect 1880 1950 1899 1984
rect 1933 1950 1952 1984
rect 1880 1894 1952 1950
rect 1880 1860 1899 1894
rect 1933 1860 1952 1894
rect 2014 2498 2708 2557
rect 2014 2464 2073 2498
rect 2107 2470 2163 2498
rect 2135 2464 2163 2470
rect 2197 2470 2253 2498
rect 2197 2464 2201 2470
rect 2014 2436 2101 2464
rect 2135 2436 2201 2464
rect 2235 2464 2253 2470
rect 2287 2470 2343 2498
rect 2287 2464 2301 2470
rect 2235 2436 2301 2464
rect 2335 2464 2343 2470
rect 2377 2470 2433 2498
rect 2467 2470 2523 2498
rect 2557 2470 2613 2498
rect 2377 2464 2401 2470
rect 2467 2464 2501 2470
rect 2557 2464 2601 2470
rect 2647 2464 2708 2498
rect 2335 2436 2401 2464
rect 2435 2436 2501 2464
rect 2535 2436 2601 2464
rect 2635 2436 2708 2464
rect 2014 2408 2708 2436
rect 2014 2374 2073 2408
rect 2107 2374 2163 2408
rect 2197 2374 2253 2408
rect 2287 2374 2343 2408
rect 2377 2374 2433 2408
rect 2467 2374 2523 2408
rect 2557 2374 2613 2408
rect 2647 2374 2708 2408
rect 2014 2370 2708 2374
rect 2014 2336 2101 2370
rect 2135 2336 2201 2370
rect 2235 2336 2301 2370
rect 2335 2336 2401 2370
rect 2435 2336 2501 2370
rect 2535 2336 2601 2370
rect 2635 2336 2708 2370
rect 2014 2318 2708 2336
rect 2014 2284 2073 2318
rect 2107 2284 2163 2318
rect 2197 2284 2253 2318
rect 2287 2284 2343 2318
rect 2377 2284 2433 2318
rect 2467 2284 2523 2318
rect 2557 2284 2613 2318
rect 2647 2284 2708 2318
rect 2014 2270 2708 2284
rect 2014 2236 2101 2270
rect 2135 2236 2201 2270
rect 2235 2236 2301 2270
rect 2335 2236 2401 2270
rect 2435 2236 2501 2270
rect 2535 2236 2601 2270
rect 2635 2236 2708 2270
rect 2014 2228 2708 2236
rect 2014 2194 2073 2228
rect 2107 2194 2163 2228
rect 2197 2194 2253 2228
rect 2287 2194 2343 2228
rect 2377 2194 2433 2228
rect 2467 2194 2523 2228
rect 2557 2194 2613 2228
rect 2647 2194 2708 2228
rect 2014 2170 2708 2194
rect 2014 2138 2101 2170
rect 2135 2138 2201 2170
rect 2014 2104 2073 2138
rect 2135 2136 2163 2138
rect 2107 2104 2163 2136
rect 2197 2136 2201 2138
rect 2235 2138 2301 2170
rect 2235 2136 2253 2138
rect 2197 2104 2253 2136
rect 2287 2136 2301 2138
rect 2335 2138 2401 2170
rect 2435 2138 2501 2170
rect 2535 2138 2601 2170
rect 2635 2138 2708 2170
rect 2335 2136 2343 2138
rect 2287 2104 2343 2136
rect 2377 2136 2401 2138
rect 2467 2136 2501 2138
rect 2557 2136 2601 2138
rect 2377 2104 2433 2136
rect 2467 2104 2523 2136
rect 2557 2104 2613 2136
rect 2647 2104 2708 2138
rect 2014 2070 2708 2104
rect 2014 2048 2101 2070
rect 2135 2048 2201 2070
rect 2014 2014 2073 2048
rect 2135 2036 2163 2048
rect 2107 2014 2163 2036
rect 2197 2036 2201 2048
rect 2235 2048 2301 2070
rect 2235 2036 2253 2048
rect 2197 2014 2253 2036
rect 2287 2036 2301 2048
rect 2335 2048 2401 2070
rect 2435 2048 2501 2070
rect 2535 2048 2601 2070
rect 2635 2048 2708 2070
rect 2335 2036 2343 2048
rect 2287 2014 2343 2036
rect 2377 2036 2401 2048
rect 2467 2036 2501 2048
rect 2557 2036 2601 2048
rect 2377 2014 2433 2036
rect 2467 2014 2523 2036
rect 2557 2014 2613 2036
rect 2647 2014 2708 2048
rect 2014 1970 2708 2014
rect 2014 1958 2101 1970
rect 2135 1958 2201 1970
rect 2014 1924 2073 1958
rect 2135 1936 2163 1958
rect 2107 1924 2163 1936
rect 2197 1936 2201 1958
rect 2235 1958 2301 1970
rect 2235 1936 2253 1958
rect 2197 1924 2253 1936
rect 2287 1936 2301 1958
rect 2335 1958 2401 1970
rect 2435 1958 2501 1970
rect 2535 1958 2601 1970
rect 2635 1958 2708 1970
rect 2335 1936 2343 1958
rect 2287 1924 2343 1936
rect 2377 1936 2401 1958
rect 2467 1936 2501 1958
rect 2557 1936 2601 1958
rect 2377 1924 2433 1936
rect 2467 1924 2523 1936
rect 2557 1924 2613 1936
rect 2647 1924 2708 1958
rect 2014 1863 2708 1924
rect 2770 2546 2789 2580
rect 2823 2546 2842 2580
rect 2770 2490 2842 2546
rect 2770 2456 2789 2490
rect 2823 2456 2842 2490
rect 2770 2400 2842 2456
rect 2770 2366 2789 2400
rect 2823 2366 2842 2400
rect 2770 2310 2842 2366
rect 2770 2276 2789 2310
rect 2823 2276 2842 2310
rect 2770 2220 2842 2276
rect 2770 2186 2789 2220
rect 2823 2186 2842 2220
rect 2770 2130 2842 2186
rect 2770 2096 2789 2130
rect 2823 2096 2842 2130
rect 2770 2040 2842 2096
rect 2770 2006 2789 2040
rect 2823 2006 2842 2040
rect 2770 1950 2842 2006
rect 2770 1916 2789 1950
rect 2823 1916 2842 1950
rect 1880 1801 1952 1860
rect 2770 1860 2842 1916
rect 2770 1826 2789 1860
rect 2823 1826 2842 1860
rect 2770 1801 2842 1826
rect 1880 1782 2842 1801
rect 1880 1748 1956 1782
rect 1990 1748 2046 1782
rect 2080 1748 2136 1782
rect 2170 1748 2226 1782
rect 2260 1748 2316 1782
rect 2350 1748 2406 1782
rect 2440 1748 2496 1782
rect 2530 1748 2586 1782
rect 2620 1748 2676 1782
rect 2710 1748 2842 1782
rect 1880 1729 2842 1748
rect 2906 2596 2939 2619
rect 2973 2596 3005 2619
rect 2906 2540 3005 2596
rect 2906 2506 2939 2540
rect 2973 2506 3005 2540
rect 2906 2450 3005 2506
rect 2906 2416 2939 2450
rect 2973 2416 3005 2450
rect 2906 2360 3005 2416
rect 2906 2326 2939 2360
rect 2973 2326 3005 2360
rect 2906 2270 3005 2326
rect 2906 2236 2939 2270
rect 2973 2236 3005 2270
rect 2906 2180 3005 2236
rect 2906 2146 2939 2180
rect 2973 2146 3005 2180
rect 2906 2090 3005 2146
rect 2906 2056 2939 2090
rect 2973 2056 3005 2090
rect 2906 2000 3005 2056
rect 2906 1966 2939 2000
rect 2973 1966 3005 2000
rect 2906 1910 3005 1966
rect 2906 1876 2939 1910
rect 2973 1876 3005 1910
rect 2906 1820 3005 1876
rect 2906 1786 2939 1820
rect 2973 1786 3005 1820
rect 2906 1730 3005 1786
rect 1717 1665 1816 1696
rect 2906 1696 2939 1730
rect 2973 1696 3005 1730
rect 2906 1665 3005 1696
rect 1717 1634 3005 1665
rect 1717 1600 1775 1634
rect 1809 1600 1865 1634
rect 1899 1600 1955 1634
rect 1989 1600 2045 1634
rect 2079 1600 2135 1634
rect 2169 1600 2225 1634
rect 2259 1600 2315 1634
rect 2349 1600 2405 1634
rect 2439 1600 2495 1634
rect 2529 1600 2585 1634
rect 2619 1600 2675 1634
rect 2709 1600 2765 1634
rect 2799 1600 2855 1634
rect 2889 1600 3005 1634
rect 1717 1566 3005 1600
rect 3105 2821 4393 2854
rect 3105 2787 3163 2821
rect 3197 2787 3253 2821
rect 3287 2787 3343 2821
rect 3377 2787 3433 2821
rect 3467 2787 3523 2821
rect 3557 2787 3613 2821
rect 3647 2787 3703 2821
rect 3737 2787 3793 2821
rect 3827 2787 3883 2821
rect 3917 2787 3973 2821
rect 4007 2787 4063 2821
rect 4097 2787 4153 2821
rect 4187 2787 4243 2821
rect 4277 2787 4393 2821
rect 3105 2755 4393 2787
rect 3105 2720 3204 2755
rect 3105 2691 3140 2720
rect 3174 2691 3204 2720
rect 4294 2720 4393 2755
rect 4294 2691 4327 2720
rect 4361 2691 4393 2720
rect 3105 2596 3140 2619
rect 3174 2596 3204 2619
rect 3105 2540 3204 2596
rect 3105 2506 3140 2540
rect 3174 2506 3204 2540
rect 3105 2450 3204 2506
rect 3105 2416 3140 2450
rect 3174 2416 3204 2450
rect 3105 2360 3204 2416
rect 3105 2326 3140 2360
rect 3174 2326 3204 2360
rect 3105 2270 3204 2326
rect 3105 2236 3140 2270
rect 3174 2236 3204 2270
rect 3105 2180 3204 2236
rect 3105 2146 3140 2180
rect 3174 2146 3204 2180
rect 3105 2090 3204 2146
rect 3105 2056 3140 2090
rect 3174 2056 3204 2090
rect 3105 2000 3204 2056
rect 3105 1966 3140 2000
rect 3174 1966 3204 2000
rect 3105 1910 3204 1966
rect 3105 1876 3140 1910
rect 3174 1876 3204 1910
rect 3105 1820 3204 1876
rect 3105 1786 3140 1820
rect 3174 1786 3204 1820
rect 3105 1730 3204 1786
rect 3105 1696 3140 1730
rect 3174 1696 3204 1730
rect 3340 2672 4158 2691
rect 3340 2638 3363 2672
rect 3397 2638 3453 2672
rect 3487 2638 3543 2672
rect 3577 2638 3633 2672
rect 3667 2638 3723 2672
rect 3757 2638 3813 2672
rect 3847 2638 3903 2672
rect 3937 2638 3993 2672
rect 4027 2638 4083 2672
rect 4117 2638 4158 2672
rect 3340 2619 4158 2638
rect 3268 2614 3340 2619
rect 3268 2580 3287 2614
rect 3321 2580 3340 2614
rect 3268 2524 3340 2580
rect 4158 2580 4230 2619
rect 3268 2490 3287 2524
rect 3321 2490 3340 2524
rect 3268 2434 3340 2490
rect 3268 2400 3287 2434
rect 3321 2400 3340 2434
rect 3268 2344 3340 2400
rect 3268 2310 3287 2344
rect 3321 2310 3340 2344
rect 3268 2254 3340 2310
rect 3268 2220 3287 2254
rect 3321 2220 3340 2254
rect 3268 2164 3340 2220
rect 3268 2130 3287 2164
rect 3321 2130 3340 2164
rect 3268 2074 3340 2130
rect 3268 2040 3287 2074
rect 3321 2040 3340 2074
rect 3268 1984 3340 2040
rect 3268 1950 3287 1984
rect 3321 1950 3340 1984
rect 3268 1894 3340 1950
rect 3268 1860 3287 1894
rect 3321 1860 3340 1894
rect 3402 2498 4096 2557
rect 3402 2464 3461 2498
rect 3495 2470 3551 2498
rect 3523 2464 3551 2470
rect 3585 2470 3641 2498
rect 3585 2464 3589 2470
rect 3402 2436 3489 2464
rect 3523 2436 3589 2464
rect 3623 2464 3641 2470
rect 3675 2470 3731 2498
rect 3675 2464 3689 2470
rect 3623 2436 3689 2464
rect 3723 2464 3731 2470
rect 3765 2470 3821 2498
rect 3855 2470 3911 2498
rect 3945 2470 4001 2498
rect 3765 2464 3789 2470
rect 3855 2464 3889 2470
rect 3945 2464 3989 2470
rect 4035 2464 4096 2498
rect 3723 2436 3789 2464
rect 3823 2436 3889 2464
rect 3923 2436 3989 2464
rect 4023 2436 4096 2464
rect 3402 2408 4096 2436
rect 3402 2374 3461 2408
rect 3495 2374 3551 2408
rect 3585 2374 3641 2408
rect 3675 2374 3731 2408
rect 3765 2374 3821 2408
rect 3855 2374 3911 2408
rect 3945 2374 4001 2408
rect 4035 2374 4096 2408
rect 3402 2370 4096 2374
rect 3402 2336 3489 2370
rect 3523 2336 3589 2370
rect 3623 2336 3689 2370
rect 3723 2336 3789 2370
rect 3823 2336 3889 2370
rect 3923 2336 3989 2370
rect 4023 2336 4096 2370
rect 3402 2318 4096 2336
rect 3402 2284 3461 2318
rect 3495 2284 3551 2318
rect 3585 2284 3641 2318
rect 3675 2284 3731 2318
rect 3765 2284 3821 2318
rect 3855 2284 3911 2318
rect 3945 2284 4001 2318
rect 4035 2284 4096 2318
rect 3402 2270 4096 2284
rect 3402 2236 3489 2270
rect 3523 2236 3589 2270
rect 3623 2236 3689 2270
rect 3723 2236 3789 2270
rect 3823 2236 3889 2270
rect 3923 2236 3989 2270
rect 4023 2236 4096 2270
rect 3402 2228 4096 2236
rect 3402 2194 3461 2228
rect 3495 2194 3551 2228
rect 3585 2194 3641 2228
rect 3675 2194 3731 2228
rect 3765 2194 3821 2228
rect 3855 2194 3911 2228
rect 3945 2194 4001 2228
rect 4035 2194 4096 2228
rect 3402 2170 4096 2194
rect 3402 2138 3489 2170
rect 3523 2138 3589 2170
rect 3402 2104 3461 2138
rect 3523 2136 3551 2138
rect 3495 2104 3551 2136
rect 3585 2136 3589 2138
rect 3623 2138 3689 2170
rect 3623 2136 3641 2138
rect 3585 2104 3641 2136
rect 3675 2136 3689 2138
rect 3723 2138 3789 2170
rect 3823 2138 3889 2170
rect 3923 2138 3989 2170
rect 4023 2138 4096 2170
rect 3723 2136 3731 2138
rect 3675 2104 3731 2136
rect 3765 2136 3789 2138
rect 3855 2136 3889 2138
rect 3945 2136 3989 2138
rect 3765 2104 3821 2136
rect 3855 2104 3911 2136
rect 3945 2104 4001 2136
rect 4035 2104 4096 2138
rect 3402 2070 4096 2104
rect 3402 2048 3489 2070
rect 3523 2048 3589 2070
rect 3402 2014 3461 2048
rect 3523 2036 3551 2048
rect 3495 2014 3551 2036
rect 3585 2036 3589 2048
rect 3623 2048 3689 2070
rect 3623 2036 3641 2048
rect 3585 2014 3641 2036
rect 3675 2036 3689 2048
rect 3723 2048 3789 2070
rect 3823 2048 3889 2070
rect 3923 2048 3989 2070
rect 4023 2048 4096 2070
rect 3723 2036 3731 2048
rect 3675 2014 3731 2036
rect 3765 2036 3789 2048
rect 3855 2036 3889 2048
rect 3945 2036 3989 2048
rect 3765 2014 3821 2036
rect 3855 2014 3911 2036
rect 3945 2014 4001 2036
rect 4035 2014 4096 2048
rect 3402 1970 4096 2014
rect 3402 1958 3489 1970
rect 3523 1958 3589 1970
rect 3402 1924 3461 1958
rect 3523 1936 3551 1958
rect 3495 1924 3551 1936
rect 3585 1936 3589 1958
rect 3623 1958 3689 1970
rect 3623 1936 3641 1958
rect 3585 1924 3641 1936
rect 3675 1936 3689 1958
rect 3723 1958 3789 1970
rect 3823 1958 3889 1970
rect 3923 1958 3989 1970
rect 4023 1958 4096 1970
rect 3723 1936 3731 1958
rect 3675 1924 3731 1936
rect 3765 1936 3789 1958
rect 3855 1936 3889 1958
rect 3945 1936 3989 1958
rect 3765 1924 3821 1936
rect 3855 1924 3911 1936
rect 3945 1924 4001 1936
rect 4035 1924 4096 1958
rect 3402 1863 4096 1924
rect 4158 2546 4177 2580
rect 4211 2546 4230 2580
rect 4158 2490 4230 2546
rect 4158 2456 4177 2490
rect 4211 2456 4230 2490
rect 4158 2400 4230 2456
rect 4158 2366 4177 2400
rect 4211 2366 4230 2400
rect 4158 2310 4230 2366
rect 4158 2276 4177 2310
rect 4211 2276 4230 2310
rect 4158 2220 4230 2276
rect 4158 2186 4177 2220
rect 4211 2186 4230 2220
rect 4158 2130 4230 2186
rect 4158 2096 4177 2130
rect 4211 2096 4230 2130
rect 4158 2040 4230 2096
rect 4158 2006 4177 2040
rect 4211 2006 4230 2040
rect 4158 1950 4230 2006
rect 4158 1916 4177 1950
rect 4211 1916 4230 1950
rect 3268 1801 3340 1860
rect 4158 1860 4230 1916
rect 4158 1826 4177 1860
rect 4211 1826 4230 1860
rect 4158 1801 4230 1826
rect 3268 1782 4230 1801
rect 3268 1748 3344 1782
rect 3378 1748 3434 1782
rect 3468 1748 3524 1782
rect 3558 1748 3614 1782
rect 3648 1748 3704 1782
rect 3738 1748 3794 1782
rect 3828 1748 3884 1782
rect 3918 1748 3974 1782
rect 4008 1748 4064 1782
rect 4098 1748 4230 1782
rect 3268 1729 4230 1748
rect 4294 2596 4327 2619
rect 4361 2596 4393 2619
rect 4294 2540 4393 2596
rect 4294 2506 4327 2540
rect 4361 2506 4393 2540
rect 4294 2450 4393 2506
rect 4294 2416 4327 2450
rect 4361 2416 4393 2450
rect 4294 2360 4393 2416
rect 4294 2326 4327 2360
rect 4361 2326 4393 2360
rect 4294 2270 4393 2326
rect 4294 2236 4327 2270
rect 4361 2236 4393 2270
rect 4294 2180 4393 2236
rect 4294 2146 4327 2180
rect 4361 2146 4393 2180
rect 4294 2090 4393 2146
rect 4294 2056 4327 2090
rect 4361 2056 4393 2090
rect 4294 2000 4393 2056
rect 4294 1966 4327 2000
rect 4361 1966 4393 2000
rect 4294 1910 4393 1966
rect 4294 1876 4327 1910
rect 4361 1876 4393 1910
rect 4294 1820 4393 1876
rect 4294 1786 4327 1820
rect 4361 1786 4393 1820
rect 4294 1730 4393 1786
rect 3105 1665 3204 1696
rect 4294 1696 4327 1730
rect 4361 1696 4393 1730
rect 4294 1665 4393 1696
rect 3105 1634 4393 1665
rect 3105 1600 3163 1634
rect 3197 1600 3253 1634
rect 3287 1600 3343 1634
rect 3377 1600 3433 1634
rect 3467 1600 3523 1634
rect 3557 1600 3613 1634
rect 3647 1600 3703 1634
rect 3737 1600 3793 1634
rect 3827 1600 3883 1634
rect 3917 1600 3973 1634
rect 4007 1600 4063 1634
rect 4097 1600 4153 1634
rect 4187 1600 4243 1634
rect 4277 1600 4393 1634
rect 3105 1566 4393 1600
rect 4493 2821 5781 2854
rect 4493 2787 4551 2821
rect 4585 2787 4641 2821
rect 4675 2787 4731 2821
rect 4765 2787 4821 2821
rect 4855 2787 4911 2821
rect 4945 2787 5001 2821
rect 5035 2787 5091 2821
rect 5125 2787 5181 2821
rect 5215 2787 5271 2821
rect 5305 2787 5361 2821
rect 5395 2787 5451 2821
rect 5485 2787 5541 2821
rect 5575 2787 5631 2821
rect 5665 2787 5781 2821
rect 4493 2755 5781 2787
rect 4493 2720 4592 2755
rect 4493 2691 4528 2720
rect 4562 2691 4592 2720
rect 5682 2720 5781 2755
rect 5682 2691 5715 2720
rect 5749 2691 5781 2720
rect 5881 2821 6043 2854
rect 6115 2821 7169 2854
rect 5881 2787 5939 2821
rect 5973 2787 6029 2821
rect 6115 2787 6119 2821
rect 6153 2787 6209 2821
rect 6243 2787 6299 2821
rect 6333 2787 6389 2821
rect 6423 2787 6479 2821
rect 6513 2787 6569 2821
rect 6603 2787 6659 2821
rect 6693 2787 6749 2821
rect 6783 2787 6839 2821
rect 6873 2787 6929 2821
rect 6963 2787 7019 2821
rect 7053 2787 7169 2821
rect 5881 2755 6043 2787
rect 6115 2755 7169 2787
rect 5881 2720 5980 2755
rect 5881 2691 5916 2720
rect 5950 2691 5980 2720
rect 7070 2720 7169 2755
rect 4493 2596 4528 2619
rect 4562 2596 4592 2619
rect 4493 2540 4592 2596
rect 4493 2506 4528 2540
rect 4562 2506 4592 2540
rect 4493 2450 4592 2506
rect 4493 2416 4528 2450
rect 4562 2416 4592 2450
rect 4493 2360 4592 2416
rect 4493 2326 4528 2360
rect 4562 2326 4592 2360
rect 4493 2270 4592 2326
rect 4493 2236 4528 2270
rect 4562 2236 4592 2270
rect 4493 2180 4592 2236
rect 4493 2146 4528 2180
rect 4562 2146 4592 2180
rect 4493 2090 4592 2146
rect 4493 2056 4528 2090
rect 4562 2056 4592 2090
rect 4493 2000 4592 2056
rect 4493 1966 4528 2000
rect 4562 1966 4592 2000
rect 4493 1910 4592 1966
rect 4493 1876 4528 1910
rect 4562 1876 4592 1910
rect 4493 1820 4592 1876
rect 4493 1786 4528 1820
rect 4562 1786 4592 1820
rect 4493 1730 4592 1786
rect 4493 1696 4528 1730
rect 4562 1696 4592 1730
rect 4728 2672 5546 2691
rect 4728 2638 4751 2672
rect 4785 2638 4841 2672
rect 4875 2638 4931 2672
rect 4965 2638 5021 2672
rect 5055 2638 5111 2672
rect 5145 2638 5201 2672
rect 5235 2638 5291 2672
rect 5325 2638 5381 2672
rect 5415 2638 5471 2672
rect 5505 2638 5546 2672
rect 4728 2619 5546 2638
rect 4656 2614 4728 2619
rect 4656 2580 4675 2614
rect 4709 2580 4728 2614
rect 4656 2524 4728 2580
rect 5546 2580 5618 2619
rect 4656 2490 4675 2524
rect 4709 2490 4728 2524
rect 4656 2434 4728 2490
rect 4656 2400 4675 2434
rect 4709 2400 4728 2434
rect 4656 2344 4728 2400
rect 4656 2310 4675 2344
rect 4709 2310 4728 2344
rect 4656 2254 4728 2310
rect 4656 2220 4675 2254
rect 4709 2220 4728 2254
rect 4656 2164 4728 2220
rect 4656 2130 4675 2164
rect 4709 2130 4728 2164
rect 4656 2074 4728 2130
rect 4656 2040 4675 2074
rect 4709 2040 4728 2074
rect 4656 1984 4728 2040
rect 4656 1950 4675 1984
rect 4709 1950 4728 1984
rect 4656 1894 4728 1950
rect 4656 1860 4675 1894
rect 4709 1860 4728 1894
rect 4790 2498 5484 2557
rect 4790 2464 4849 2498
rect 4883 2470 4939 2498
rect 4911 2464 4939 2470
rect 4973 2470 5029 2498
rect 4973 2464 4977 2470
rect 4790 2436 4877 2464
rect 4911 2436 4977 2464
rect 5011 2464 5029 2470
rect 5063 2470 5119 2498
rect 5063 2464 5077 2470
rect 5011 2436 5077 2464
rect 5111 2464 5119 2470
rect 5153 2470 5209 2498
rect 5243 2470 5299 2498
rect 5333 2470 5389 2498
rect 5153 2464 5177 2470
rect 5243 2464 5277 2470
rect 5333 2464 5377 2470
rect 5423 2464 5484 2498
rect 5111 2436 5177 2464
rect 5211 2436 5277 2464
rect 5311 2436 5377 2464
rect 5411 2436 5484 2464
rect 4790 2408 5484 2436
rect 4790 2374 4849 2408
rect 4883 2374 4939 2408
rect 4973 2374 5029 2408
rect 5063 2374 5119 2408
rect 5153 2374 5209 2408
rect 5243 2374 5299 2408
rect 5333 2374 5389 2408
rect 5423 2374 5484 2408
rect 4790 2370 5484 2374
rect 4790 2336 4877 2370
rect 4911 2336 4977 2370
rect 5011 2336 5077 2370
rect 5111 2336 5177 2370
rect 5211 2336 5277 2370
rect 5311 2336 5377 2370
rect 5411 2336 5484 2370
rect 4790 2318 5484 2336
rect 4790 2284 4849 2318
rect 4883 2284 4939 2318
rect 4973 2284 5029 2318
rect 5063 2284 5119 2318
rect 5153 2284 5209 2318
rect 5243 2284 5299 2318
rect 5333 2284 5389 2318
rect 5423 2284 5484 2318
rect 4790 2270 5484 2284
rect 4790 2236 4877 2270
rect 4911 2236 4977 2270
rect 5011 2236 5077 2270
rect 5111 2236 5177 2270
rect 5211 2236 5277 2270
rect 5311 2236 5377 2270
rect 5411 2236 5484 2270
rect 4790 2228 5484 2236
rect 4790 2194 4849 2228
rect 4883 2194 4939 2228
rect 4973 2194 5029 2228
rect 5063 2194 5119 2228
rect 5153 2194 5209 2228
rect 5243 2194 5299 2228
rect 5333 2194 5389 2228
rect 5423 2194 5484 2228
rect 4790 2170 5484 2194
rect 4790 2138 4877 2170
rect 4911 2138 4977 2170
rect 4790 2104 4849 2138
rect 4911 2136 4939 2138
rect 4883 2104 4939 2136
rect 4973 2136 4977 2138
rect 5011 2138 5077 2170
rect 5011 2136 5029 2138
rect 4973 2104 5029 2136
rect 5063 2136 5077 2138
rect 5111 2138 5177 2170
rect 5211 2138 5277 2170
rect 5311 2138 5377 2170
rect 5411 2138 5484 2170
rect 5111 2136 5119 2138
rect 5063 2104 5119 2136
rect 5153 2136 5177 2138
rect 5243 2136 5277 2138
rect 5333 2136 5377 2138
rect 5153 2104 5209 2136
rect 5243 2104 5299 2136
rect 5333 2104 5389 2136
rect 5423 2104 5484 2138
rect 4790 2070 5484 2104
rect 4790 2048 4877 2070
rect 4911 2048 4977 2070
rect 4790 2014 4849 2048
rect 4911 2036 4939 2048
rect 4883 2014 4939 2036
rect 4973 2036 4977 2048
rect 5011 2048 5077 2070
rect 5011 2036 5029 2048
rect 4973 2014 5029 2036
rect 5063 2036 5077 2048
rect 5111 2048 5177 2070
rect 5211 2048 5277 2070
rect 5311 2048 5377 2070
rect 5411 2048 5484 2070
rect 5111 2036 5119 2048
rect 5063 2014 5119 2036
rect 5153 2036 5177 2048
rect 5243 2036 5277 2048
rect 5333 2036 5377 2048
rect 5153 2014 5209 2036
rect 5243 2014 5299 2036
rect 5333 2014 5389 2036
rect 5423 2014 5484 2048
rect 4790 1970 5484 2014
rect 4790 1958 4877 1970
rect 4911 1958 4977 1970
rect 4790 1924 4849 1958
rect 4911 1936 4939 1958
rect 4883 1924 4939 1936
rect 4973 1936 4977 1958
rect 5011 1958 5077 1970
rect 5011 1936 5029 1958
rect 4973 1924 5029 1936
rect 5063 1936 5077 1958
rect 5111 1958 5177 1970
rect 5211 1958 5277 1970
rect 5311 1958 5377 1970
rect 5411 1958 5484 1970
rect 5111 1936 5119 1958
rect 5063 1924 5119 1936
rect 5153 1936 5177 1958
rect 5243 1936 5277 1958
rect 5333 1936 5377 1958
rect 5153 1924 5209 1936
rect 5243 1924 5299 1936
rect 5333 1924 5389 1936
rect 5423 1924 5484 1958
rect 4790 1863 5484 1924
rect 5546 2546 5565 2580
rect 5599 2546 5618 2580
rect 5546 2490 5618 2546
rect 5546 2456 5565 2490
rect 5599 2456 5618 2490
rect 5546 2400 5618 2456
rect 5546 2366 5565 2400
rect 5599 2366 5618 2400
rect 5546 2310 5618 2366
rect 5546 2276 5565 2310
rect 5599 2276 5618 2310
rect 5546 2220 5618 2276
rect 5546 2186 5565 2220
rect 5599 2186 5618 2220
rect 5546 2130 5618 2186
rect 5546 2096 5565 2130
rect 5599 2096 5618 2130
rect 5546 2040 5618 2096
rect 5546 2006 5565 2040
rect 5599 2006 5618 2040
rect 5546 1950 5618 2006
rect 5546 1916 5565 1950
rect 5599 1916 5618 1950
rect 4656 1801 4728 1860
rect 5546 1860 5618 1916
rect 5546 1826 5565 1860
rect 5599 1826 5618 1860
rect 5546 1801 5618 1826
rect 4656 1782 5618 1801
rect 4656 1748 4732 1782
rect 4766 1748 4822 1782
rect 4856 1748 4912 1782
rect 4946 1748 5002 1782
rect 5036 1748 5092 1782
rect 5126 1748 5182 1782
rect 5216 1748 5272 1782
rect 5306 1748 5362 1782
rect 5396 1748 5452 1782
rect 5486 1748 5618 1782
rect 4656 1729 5618 1748
rect 5979 2619 5980 2691
rect 6115 2672 7006 2691
rect 6115 2638 6139 2672
rect 6173 2638 6229 2672
rect 6263 2638 6319 2672
rect 6353 2638 6409 2672
rect 6443 2638 6499 2672
rect 6533 2638 6589 2672
rect 6623 2638 6679 2672
rect 6713 2638 6769 2672
rect 6803 2638 6859 2672
rect 6893 2638 7006 2672
rect 6115 2619 7006 2638
rect 5682 2596 5715 2619
rect 5749 2596 5781 2619
rect 5682 2540 5781 2596
rect 5682 2506 5715 2540
rect 5749 2506 5781 2540
rect 5682 2450 5781 2506
rect 5682 2416 5715 2450
rect 5749 2416 5781 2450
rect 5682 2360 5781 2416
rect 5682 2326 5715 2360
rect 5749 2326 5781 2360
rect 5682 2270 5781 2326
rect 5682 2236 5715 2270
rect 5749 2236 5781 2270
rect 5682 2180 5781 2236
rect 5682 2146 5715 2180
rect 5749 2146 5781 2180
rect 5682 2090 5781 2146
rect 5682 2056 5715 2090
rect 5749 2056 5781 2090
rect 5682 2000 5781 2056
rect 5682 1966 5715 2000
rect 5749 1966 5781 2000
rect 5682 1910 5781 1966
rect 5682 1876 5715 1910
rect 5749 1876 5781 1910
rect 5682 1820 5781 1876
rect 5682 1786 5715 1820
rect 5749 1786 5781 1820
rect 5682 1730 5781 1786
rect 4493 1665 4592 1696
rect 5682 1696 5715 1730
rect 5749 1696 5781 1730
rect 5682 1665 5781 1696
rect 4493 1634 5781 1665
rect 4493 1600 4551 1634
rect 4585 1600 4641 1634
rect 4675 1600 4731 1634
rect 4765 1600 4821 1634
rect 4855 1600 4911 1634
rect 4945 1600 5001 1634
rect 5035 1600 5091 1634
rect 5125 1600 5181 1634
rect 5215 1600 5271 1634
rect 5305 1600 5361 1634
rect 5395 1600 5451 1634
rect 5485 1600 5541 1634
rect 5575 1600 5631 1634
rect 5665 1600 5781 1634
rect 4493 1566 5781 1600
rect 5881 2596 5916 2619
rect 5950 2596 5980 2619
rect 5881 2540 5980 2596
rect 5881 2506 5916 2540
rect 5950 2506 5980 2540
rect 5881 2450 5980 2506
rect 5881 2416 5916 2450
rect 5950 2416 5980 2450
rect 5881 2360 5980 2416
rect 5881 2326 5916 2360
rect 5950 2326 5980 2360
rect 5881 2270 5980 2326
rect 5881 2236 5916 2270
rect 5950 2236 5980 2270
rect 5881 2180 5980 2236
rect 5881 2146 5916 2180
rect 5950 2146 5980 2180
rect 5881 2090 5980 2146
rect 5881 2056 5916 2090
rect 5950 2056 5980 2090
rect 5881 2000 5980 2056
rect 5881 1966 5916 2000
rect 5950 1966 5980 2000
rect 5881 1910 5980 1966
rect 5881 1876 5916 1910
rect 5950 1876 5980 1910
rect 5881 1820 5980 1876
rect 5881 1786 5916 1820
rect 5950 1786 5980 1820
rect 5881 1730 5980 1786
rect 5881 1696 5916 1730
rect 5950 1696 5980 1730
rect 6044 2614 6116 2619
rect 6044 2580 6063 2614
rect 6097 2580 6116 2614
rect 6044 2524 6116 2580
rect 6934 2580 7006 2619
rect 6044 2490 6063 2524
rect 6097 2490 6116 2524
rect 6044 2434 6116 2490
rect 6044 2400 6063 2434
rect 6097 2400 6116 2434
rect 6044 2344 6116 2400
rect 6044 2310 6063 2344
rect 6097 2310 6116 2344
rect 6044 2254 6116 2310
rect 6044 2220 6063 2254
rect 6097 2220 6116 2254
rect 6044 2164 6116 2220
rect 6044 2130 6063 2164
rect 6097 2130 6116 2164
rect 6044 2074 6116 2130
rect 6044 2040 6063 2074
rect 6097 2040 6116 2074
rect 6044 1984 6116 2040
rect 6044 1950 6063 1984
rect 6097 1950 6116 1984
rect 6044 1894 6116 1950
rect 6044 1860 6063 1894
rect 6097 1860 6116 1894
rect 6178 2498 6872 2557
rect 6178 2464 6237 2498
rect 6271 2470 6327 2498
rect 6299 2464 6327 2470
rect 6361 2470 6417 2498
rect 6361 2464 6365 2470
rect 6178 2436 6265 2464
rect 6299 2436 6365 2464
rect 6399 2464 6417 2470
rect 6451 2470 6507 2498
rect 6451 2464 6465 2470
rect 6399 2436 6465 2464
rect 6499 2464 6507 2470
rect 6541 2470 6597 2498
rect 6631 2470 6687 2498
rect 6721 2470 6777 2498
rect 6541 2464 6565 2470
rect 6631 2464 6665 2470
rect 6721 2464 6765 2470
rect 6811 2464 6872 2498
rect 6499 2436 6565 2464
rect 6599 2436 6665 2464
rect 6699 2436 6765 2464
rect 6799 2436 6872 2464
rect 6178 2408 6872 2436
rect 6178 2374 6237 2408
rect 6271 2374 6327 2408
rect 6361 2374 6417 2408
rect 6451 2374 6507 2408
rect 6541 2374 6597 2408
rect 6631 2374 6687 2408
rect 6721 2374 6777 2408
rect 6811 2374 6872 2408
rect 6178 2370 6872 2374
rect 6178 2336 6265 2370
rect 6299 2336 6365 2370
rect 6399 2336 6465 2370
rect 6499 2336 6565 2370
rect 6599 2336 6665 2370
rect 6699 2336 6765 2370
rect 6799 2336 6872 2370
rect 6178 2318 6872 2336
rect 6178 2284 6237 2318
rect 6271 2284 6327 2318
rect 6361 2284 6417 2318
rect 6451 2284 6507 2318
rect 6541 2284 6597 2318
rect 6631 2284 6687 2318
rect 6721 2284 6777 2318
rect 6811 2284 6872 2318
rect 6178 2270 6872 2284
rect 6178 2236 6265 2270
rect 6299 2236 6365 2270
rect 6399 2236 6465 2270
rect 6499 2236 6565 2270
rect 6599 2236 6665 2270
rect 6699 2236 6765 2270
rect 6799 2236 6872 2270
rect 6178 2228 6872 2236
rect 6178 2194 6237 2228
rect 6271 2194 6327 2228
rect 6361 2194 6417 2228
rect 6451 2194 6507 2228
rect 6541 2194 6597 2228
rect 6631 2194 6687 2228
rect 6721 2194 6777 2228
rect 6811 2194 6872 2228
rect 6178 2170 6872 2194
rect 6178 2138 6265 2170
rect 6299 2138 6365 2170
rect 6178 2104 6237 2138
rect 6299 2136 6327 2138
rect 6271 2104 6327 2136
rect 6361 2136 6365 2138
rect 6399 2138 6465 2170
rect 6399 2136 6417 2138
rect 6361 2104 6417 2136
rect 6451 2136 6465 2138
rect 6499 2138 6565 2170
rect 6599 2138 6665 2170
rect 6699 2138 6765 2170
rect 6799 2138 6872 2170
rect 6499 2136 6507 2138
rect 6451 2104 6507 2136
rect 6541 2136 6565 2138
rect 6631 2136 6665 2138
rect 6721 2136 6765 2138
rect 6541 2104 6597 2136
rect 6631 2104 6687 2136
rect 6721 2104 6777 2136
rect 6811 2104 6872 2138
rect 6178 2070 6872 2104
rect 6178 2048 6265 2070
rect 6299 2048 6365 2070
rect 6178 2014 6237 2048
rect 6299 2036 6327 2048
rect 6271 2014 6327 2036
rect 6361 2036 6365 2048
rect 6399 2048 6465 2070
rect 6399 2036 6417 2048
rect 6361 2014 6417 2036
rect 6451 2036 6465 2048
rect 6499 2048 6565 2070
rect 6599 2048 6665 2070
rect 6699 2048 6765 2070
rect 6799 2048 6872 2070
rect 6499 2036 6507 2048
rect 6451 2014 6507 2036
rect 6541 2036 6565 2048
rect 6631 2036 6665 2048
rect 6721 2036 6765 2048
rect 6541 2014 6597 2036
rect 6631 2014 6687 2036
rect 6721 2014 6777 2036
rect 6811 2014 6872 2048
rect 6178 1970 6872 2014
rect 6178 1958 6265 1970
rect 6299 1958 6365 1970
rect 6178 1924 6237 1958
rect 6299 1936 6327 1958
rect 6271 1924 6327 1936
rect 6361 1936 6365 1958
rect 6399 1958 6465 1970
rect 6399 1936 6417 1958
rect 6361 1924 6417 1936
rect 6451 1936 6465 1958
rect 6499 1958 6565 1970
rect 6599 1958 6665 1970
rect 6699 1958 6765 1970
rect 6799 1958 6872 1970
rect 6499 1936 6507 1958
rect 6451 1924 6507 1936
rect 6541 1936 6565 1958
rect 6631 1936 6665 1958
rect 6721 1936 6765 1958
rect 6541 1924 6597 1936
rect 6631 1924 6687 1936
rect 6721 1924 6777 1936
rect 6811 1924 6872 1958
rect 6178 1863 6872 1924
rect 6934 2546 6953 2580
rect 6987 2546 7006 2580
rect 6934 2490 7006 2546
rect 6934 2456 6953 2490
rect 6987 2456 7006 2490
rect 6934 2400 7006 2456
rect 6934 2366 6953 2400
rect 6987 2366 7006 2400
rect 6934 2310 7006 2366
rect 6934 2276 6953 2310
rect 6987 2276 7006 2310
rect 6934 2220 7006 2276
rect 6934 2186 6953 2220
rect 6987 2186 7006 2220
rect 6934 2130 7006 2186
rect 6934 2096 6953 2130
rect 6987 2096 7006 2130
rect 6934 2040 7006 2096
rect 6934 2006 6953 2040
rect 6987 2006 7006 2040
rect 6934 1950 7006 2006
rect 6934 1916 6953 1950
rect 6987 1916 7006 1950
rect 6044 1801 6116 1860
rect 6934 1860 7006 1916
rect 6934 1826 6953 1860
rect 6987 1826 7006 1860
rect 6934 1801 7006 1826
rect 6044 1782 7006 1801
rect 6044 1748 6120 1782
rect 6154 1748 6210 1782
rect 6244 1748 6300 1782
rect 6334 1748 6390 1782
rect 6424 1748 6480 1782
rect 6514 1748 6570 1782
rect 6604 1748 6660 1782
rect 6694 1748 6750 1782
rect 6784 1748 6840 1782
rect 6874 1748 7006 1782
rect 6044 1729 7006 1748
rect 7070 2686 7103 2720
rect 7137 2686 7169 2720
rect 7070 2630 7169 2686
rect 7070 2596 7103 2630
rect 7137 2596 7169 2630
rect 7070 2540 7169 2596
rect 7070 2506 7103 2540
rect 7137 2506 7169 2540
rect 7070 2450 7169 2506
rect 7070 2416 7103 2450
rect 7137 2416 7169 2450
rect 7070 2360 7169 2416
rect 7070 2326 7103 2360
rect 7137 2326 7169 2360
rect 7070 2270 7169 2326
rect 7070 2236 7103 2270
rect 7137 2236 7169 2270
rect 7070 2180 7169 2236
rect 7070 2146 7103 2180
rect 7137 2146 7169 2180
rect 7070 2090 7169 2146
rect 7070 2056 7103 2090
rect 7137 2056 7169 2090
rect 7070 2000 7169 2056
rect 7070 1966 7103 2000
rect 7137 1966 7169 2000
rect 7070 1910 7169 1966
rect 7070 1876 7103 1910
rect 7137 1876 7169 1910
rect 7070 1820 7169 1876
rect 7070 1786 7103 1820
rect 7137 1786 7169 1820
rect 7070 1730 7169 1786
rect 5881 1665 5980 1696
rect 7070 1696 7103 1730
rect 7137 1696 7169 1730
rect 7070 1665 7169 1696
rect 5881 1634 7169 1665
rect 5881 1600 5939 1634
rect 5973 1600 6029 1634
rect 6063 1600 6119 1634
rect 6153 1600 6209 1634
rect 6243 1600 6299 1634
rect 6333 1600 6389 1634
rect 6423 1600 6479 1634
rect 6513 1600 6569 1634
rect 6603 1600 6659 1634
rect 6693 1600 6749 1634
rect 6783 1600 6839 1634
rect 6873 1600 6929 1634
rect 6963 1600 7019 1634
rect 7053 1600 7169 1634
rect 5881 1566 7169 1600
rect -17937 -401 -17903 -375
rect 9167 -401 9201 -375
rect -17937 -435 -17877 -401
rect 9141 -435 9201 -401
<< viali >>
rect -17500 22657 -17440 22691
rect -17440 22657 8642 22691
rect 8642 22657 8702 22691
rect -17500 22631 -17466 22657
rect -17500 20912 -17466 22631
rect 8668 22631 8702 22657
rect -17337 22507 -16940 22545
rect -13538 22507 -13141 22545
rect -13001 22507 -12604 22545
rect -9202 22507 -8805 22545
rect -8665 22507 -8268 22545
rect -4866 22507 -4469 22545
rect -4329 22507 -3932 22545
rect -530 22507 -133 22545
rect 7 22507 404 22545
rect 3806 22507 4203 22545
rect 4343 22507 4740 22545
rect 8142 22507 8539 22545
rect -17337 22341 -16940 22379
rect -13538 22341 -13141 22379
rect -13001 22341 -12604 22379
rect -9202 22341 -8805 22379
rect -8665 22341 -8268 22379
rect -4866 22341 -4469 22379
rect -4329 22341 -3932 22379
rect -530 22341 -133 22379
rect 7 22341 404 22379
rect 3806 22341 4203 22379
rect 4343 22341 4740 22379
rect 8142 22341 8539 22379
rect -17337 22175 -16940 22213
rect -13538 22175 -13141 22213
rect -13001 22175 -12604 22213
rect -9202 22175 -8805 22213
rect -8665 22175 -8268 22213
rect -4866 22175 -4469 22213
rect -4329 22175 -3932 22213
rect -530 22175 -133 22213
rect 7 22175 404 22213
rect 3806 22175 4203 22213
rect 4343 22175 4740 22213
rect 8142 22175 8539 22213
rect -17337 22009 -16940 22047
rect -13538 22009 -13141 22047
rect -13001 22009 -12604 22047
rect -9202 22009 -8805 22047
rect -8665 22009 -8268 22047
rect -4866 22009 -4469 22047
rect -4329 22009 -3932 22047
rect -530 22009 -133 22047
rect 7 22009 404 22047
rect 3806 22009 4203 22047
rect 4343 22009 4740 22047
rect 8142 22009 8539 22047
rect -17337 21843 -16940 21881
rect -13538 21843 -13141 21881
rect -13001 21843 -12604 21881
rect -9202 21843 -8805 21881
rect -8665 21843 -8268 21881
rect -4866 21843 -4469 21881
rect -4329 21843 -3932 21881
rect -530 21843 -133 21881
rect 7 21843 404 21881
rect 3806 21843 4203 21881
rect 4343 21843 4740 21881
rect 8142 21843 8539 21881
rect -17337 21677 -16940 21715
rect -13538 21677 -13141 21715
rect -13001 21677 -12604 21715
rect -9202 21677 -8805 21715
rect -8665 21677 -8268 21715
rect -4866 21677 -4469 21715
rect -4329 21677 -3932 21715
rect -530 21677 -133 21715
rect 7 21677 404 21715
rect 3806 21677 4203 21715
rect 4343 21677 4740 21715
rect 8142 21677 8539 21715
rect -17337 21511 -16940 21549
rect -13538 21511 -13141 21549
rect -13001 21511 -12604 21549
rect -9202 21511 -8805 21549
rect -8665 21511 -8268 21549
rect -4866 21511 -4469 21549
rect -4329 21511 -3932 21549
rect -530 21511 -133 21549
rect 7 21511 404 21549
rect 3806 21511 4203 21549
rect 4343 21511 4740 21549
rect 8142 21511 8539 21549
rect -17337 21345 -16940 21383
rect -13538 21345 -13141 21383
rect -13001 21345 -12604 21383
rect -9202 21345 -8805 21383
rect -8665 21345 -8268 21383
rect -4866 21345 -4469 21383
rect -4329 21345 -3932 21383
rect -530 21345 -133 21383
rect 7 21345 404 21383
rect 3806 21345 4203 21383
rect 4343 21345 4740 21383
rect 8142 21345 8539 21383
rect -17337 21179 -16940 21217
rect -13538 21179 -13141 21217
rect -13001 21179 -12604 21217
rect -9202 21179 -8805 21217
rect -8665 21179 -8268 21217
rect -4866 21179 -4469 21217
rect -4329 21179 -3932 21217
rect -530 21179 -133 21217
rect 7 21179 404 21217
rect 3806 21179 4203 21217
rect 4343 21179 4740 21217
rect 8142 21179 8539 21217
rect -17337 21013 -16940 21051
rect -13538 21013 -13141 21051
rect -13001 21013 -12604 21051
rect -9202 21013 -8805 21051
rect -8665 21013 -8268 21051
rect -4866 21013 -4469 21051
rect -4329 21013 -3932 21051
rect -530 21013 -133 21051
rect 7 21013 404 21051
rect 3806 21013 4203 21051
rect 4343 21013 4740 21051
rect 8142 21013 8539 21051
rect -17500 20886 -17466 20912
rect 8668 20912 8702 22631
rect 8668 20886 8702 20912
rect -17500 20852 -17440 20886
rect -17440 20852 8642 20886
rect 8642 20852 8702 20886
rect -13149 20761 -13053 20795
rect -13053 20761 8591 20795
rect 8591 20761 8687 20795
rect -13149 20699 -13115 20761
rect -13149 19399 -13115 20699
rect 8653 20699 8687 20761
rect -13001 20611 -12604 20649
rect -9202 20611 -8805 20649
rect -8665 20611 -8268 20649
rect -4866 20611 -4469 20649
rect -4329 20611 -3932 20649
rect -530 20611 -133 20649
rect 7 20611 404 20649
rect 3806 20611 4203 20649
rect 4343 20611 4740 20649
rect 8142 20611 8539 20649
rect -13001 20445 -12604 20483
rect -9202 20445 -8805 20483
rect -8665 20445 -8268 20483
rect -4866 20445 -4469 20483
rect -4329 20445 -3932 20483
rect -530 20445 -133 20483
rect 7 20445 404 20483
rect 3806 20445 4203 20483
rect 4343 20445 4740 20483
rect 8142 20445 8539 20483
rect -13001 20279 -12604 20317
rect -9202 20279 -8805 20317
rect -8665 20279 -8268 20317
rect -4866 20279 -4469 20317
rect -4329 20279 -3932 20317
rect -530 20279 -133 20317
rect 7 20279 404 20317
rect 3806 20279 4203 20317
rect 4343 20279 4740 20317
rect 8142 20279 8539 20317
rect -13001 20113 -12604 20151
rect -9202 20113 -8805 20151
rect -8665 20113 -8268 20151
rect -4866 20113 -4469 20151
rect -4329 20113 -3932 20151
rect -530 20113 -133 20151
rect 7 20113 404 20151
rect 3806 20113 4203 20151
rect 4343 20113 4740 20151
rect 8142 20113 8539 20151
rect -13001 19947 -12604 19985
rect -9202 19947 -8805 19985
rect -8665 19947 -8268 19985
rect -4866 19947 -4469 19985
rect -4329 19947 -3932 19985
rect -530 19947 -133 19985
rect 7 19947 404 19985
rect 3806 19947 4203 19985
rect 4343 19947 4740 19985
rect 8142 19947 8539 19985
rect -13001 19781 -12604 19819
rect -9202 19781 -8805 19819
rect -8665 19781 -8268 19819
rect -4866 19781 -4469 19819
rect -4329 19781 -3932 19819
rect -530 19781 -133 19819
rect 7 19781 404 19819
rect 3806 19781 4203 19819
rect 4343 19781 4740 19819
rect 8142 19781 8539 19819
rect -13001 19615 -12604 19653
rect -9202 19615 -8805 19653
rect -8665 19615 -8268 19653
rect -4866 19615 -4469 19653
rect -4329 19615 -3932 19653
rect -530 19615 -133 19653
rect 7 19615 404 19653
rect 3806 19615 4203 19653
rect 4343 19615 4740 19653
rect 8142 19615 8539 19653
rect -13001 19449 -12604 19487
rect -9202 19449 -8805 19487
rect -8665 19449 -8268 19487
rect -4866 19449 -4469 19487
rect -4329 19449 -3932 19487
rect -530 19449 -133 19487
rect 7 19449 404 19487
rect 3806 19449 4203 19487
rect 4343 19449 4740 19487
rect 8142 19449 8539 19487
rect -13149 19337 -13115 19399
rect 8653 19399 8687 20699
rect 8653 19337 8687 19399
rect -13149 19303 -13053 19337
rect -13053 19303 8591 19337
rect 8591 19303 8687 19337
rect -7017 19047 -6620 19085
rect -4938 19047 -4541 19085
rect -4401 19047 -4004 19085
rect -2322 19047 -1925 19085
rect -1785 19047 -1388 19085
rect 294 19047 691 19085
rect 831 19047 1228 19085
rect 2910 19047 3307 19085
rect 3447 19047 3844 19085
rect 5526 19047 5923 19085
rect 6063 19047 6460 19085
rect 8142 19047 8539 19085
rect -7017 18881 -6620 18919
rect -4938 18881 -4541 18919
rect -4401 18881 -4004 18919
rect -2322 18881 -1925 18919
rect -1785 18881 -1388 18919
rect 294 18881 691 18919
rect 831 18881 1228 18919
rect 2910 18881 3307 18919
rect 3447 18881 3844 18919
rect 5526 18881 5923 18919
rect 6063 18881 6460 18919
rect 8142 18881 8539 18919
rect -7017 18715 -6620 18753
rect -4938 18715 -4541 18753
rect -4401 18715 -4004 18753
rect -2322 18715 -1925 18753
rect -1785 18715 -1388 18753
rect 294 18715 691 18753
rect 831 18715 1228 18753
rect 2910 18715 3307 18753
rect 3447 18715 3844 18753
rect 5526 18715 5923 18753
rect 6063 18715 6460 18753
rect 8142 18715 8539 18753
rect -7017 18549 -6620 18587
rect -4938 18549 -4541 18587
rect -4401 18549 -4004 18587
rect -2322 18549 -1925 18587
rect -1785 18549 -1388 18587
rect 294 18549 691 18587
rect 831 18549 1228 18587
rect 2910 18549 3307 18587
rect 3447 18549 3844 18587
rect 5526 18549 5923 18587
rect 6063 18549 6460 18587
rect 8142 18549 8539 18587
rect -7017 18383 -6620 18421
rect -4938 18383 -4541 18421
rect -4401 18383 -4004 18421
rect -2322 18383 -1925 18421
rect -1785 18383 -1388 18421
rect 294 18383 691 18421
rect 831 18383 1228 18421
rect 2910 18383 3307 18421
rect 3447 18383 3844 18421
rect 5526 18383 5923 18421
rect 6063 18383 6460 18421
rect 8142 18383 8539 18421
rect -7017 18217 -6620 18255
rect -4938 18217 -4541 18255
rect -4401 18217 -4004 18255
rect -2322 18217 -1925 18255
rect -1785 18217 -1388 18255
rect 294 18217 691 18255
rect 831 18217 1228 18255
rect 2910 18217 3307 18255
rect 3447 18217 3844 18255
rect 5526 18217 5923 18255
rect 6063 18217 6460 18255
rect 8142 18217 8539 18255
rect -7017 18051 -6620 18089
rect -4938 18051 -4541 18089
rect -4401 18051 -4004 18089
rect -2322 18051 -1925 18089
rect -1785 18051 -1388 18089
rect 294 18051 691 18089
rect 831 18051 1228 18089
rect 2910 18051 3307 18089
rect 3447 18051 3844 18089
rect 5526 18051 5923 18089
rect 6063 18051 6460 18089
rect 8142 18051 8539 18089
rect -7017 17885 -6620 17923
rect -4938 17885 -4541 17923
rect -4401 17885 -4004 17923
rect -2322 17885 -1925 17923
rect -1785 17885 -1388 17923
rect 294 17885 691 17923
rect 831 17885 1228 17923
rect 2910 17885 3307 17923
rect 3447 17885 3844 17923
rect 5526 17885 5923 17923
rect 6063 17885 6460 17923
rect 8142 17885 8539 17923
rect -16699 17607 -16606 17641
rect -16606 17607 -7986 17641
rect -7986 17607 -7901 17641
rect -16699 17581 -16665 17607
rect -16699 15724 -16665 17581
rect -7935 17581 -7901 17607
rect -16517 17513 -16483 17547
rect -8109 17513 -8075 17547
rect -16517 17278 -16483 17454
rect -16429 17278 -16395 17454
rect -14371 17278 -14337 17454
rect -12313 17278 -12279 17454
rect -10255 17278 -10221 17454
rect -8197 17278 -8163 17454
rect -8109 17278 -8075 17454
rect -15875 17185 -14891 17219
rect -13817 17185 -12833 17219
rect -11759 17185 -10775 17219
rect -9701 17185 -8717 17219
rect -15875 17034 -14891 17068
rect -13817 17034 -12833 17068
rect -11759 17034 -10775 17068
rect -9701 17034 -8717 17068
rect -16517 16799 -16483 16975
rect -16429 16799 -16395 16975
rect -14371 16799 -14337 16975
rect -12313 16799 -12279 16975
rect -10255 16799 -10221 16975
rect -8197 16799 -8163 16975
rect -8109 16799 -8075 16975
rect -15875 16706 -14891 16740
rect -13817 16706 -12833 16740
rect -11759 16706 -10775 16740
rect -9701 16706 -8717 16740
rect -16517 16635 -16483 16669
rect -8109 16635 -8075 16669
rect -15875 16564 -14891 16598
rect -13817 16564 -12833 16598
rect -11759 16564 -10775 16598
rect -9701 16564 -8717 16598
rect -16517 16329 -16483 16505
rect -16429 16329 -16395 16505
rect -14371 16329 -14337 16505
rect -12313 16329 -12279 16505
rect -10255 16329 -10221 16505
rect -8197 16329 -8163 16505
rect -8109 16329 -8075 16505
rect -15875 16236 -14891 16270
rect -13817 16236 -12833 16270
rect -11759 16236 -10775 16270
rect -9701 16236 -8717 16270
rect -15875 16085 -14891 16119
rect -13817 16085 -12833 16119
rect -11759 16085 -10775 16119
rect -9701 16085 -8717 16119
rect -16517 15850 -16483 16026
rect -16429 15850 -16395 16026
rect -14371 15850 -14337 16026
rect -12313 15850 -12279 16026
rect -10255 15850 -10221 16026
rect -8197 15850 -8163 16026
rect -8109 15850 -8075 16026
rect -16517 15757 -16483 15791
rect -8109 15757 -8075 15791
rect -16699 15698 -16665 15724
rect -7935 15724 -7901 17581
rect -1270 17574 -1210 17608
rect -1210 17574 -404 17608
rect -404 17574 -344 17608
rect -7935 15698 -7901 15724
rect -16699 15664 -16606 15698
rect -16606 15664 -7986 15698
rect -7986 15664 -7901 15698
rect -7670 17518 -7585 17552
rect -7585 17518 -3081 17552
rect -3081 17518 -2996 17552
rect -7670 17492 -7636 17518
rect -7670 15718 -7636 17492
rect -3030 17492 -2996 17518
rect -7496 17419 -7462 17453
rect -3204 17419 -3170 17453
rect -7496 17184 -7462 17360
rect -7408 17184 -7374 17360
rect -5350 17184 -5316 17360
rect -3292 17184 -3258 17360
rect -3204 17184 -3170 17360
rect -6854 17091 -5870 17125
rect -4796 17091 -3812 17125
rect -7496 16987 -7462 17021
rect -3204 16987 -3170 17021
rect -7496 16752 -7462 16928
rect -7408 16752 -7374 16928
rect -5350 16752 -5316 16928
rect -3292 16752 -3258 16928
rect -3204 16752 -3170 16928
rect -6854 16659 -5870 16693
rect -4796 16659 -3812 16693
rect -6854 16517 -5870 16551
rect -4796 16517 -3812 16551
rect -7496 16282 -7462 16458
rect -7408 16282 -7374 16458
rect -5350 16282 -5316 16458
rect -3292 16282 -3258 16458
rect -3204 16282 -3170 16458
rect -7496 16189 -7462 16223
rect -3204 16189 -3170 16223
rect -6854 16085 -5870 16119
rect -4796 16085 -3812 16119
rect -7496 15850 -7462 16026
rect -7408 15850 -7374 16026
rect -5350 15850 -5316 16026
rect -3292 15850 -3258 16026
rect -3204 15850 -3170 16026
rect -7496 15757 -7462 15791
rect -3204 15757 -3170 15791
rect -7670 15692 -7636 15718
rect -3030 15718 -2996 17492
rect -1270 17541 -1236 17574
rect -1270 16854 -1236 17541
rect -378 17541 -344 17574
rect -1170 17490 -1136 17524
rect -978 17490 -894 17524
rect -720 17490 -636 17524
rect -478 17490 -444 17524
rect -1170 17264 -1136 17440
rect -1082 17264 -1048 17440
rect -824 17264 -790 17440
rect -566 17264 -532 17440
rect -478 17264 -444 17440
rect -978 17180 -894 17214
rect -720 17180 -636 17214
rect -1170 16954 -1136 17130
rect -1082 16954 -1048 17130
rect -824 16954 -790 17130
rect -566 16954 -532 17130
rect -478 16954 -444 17130
rect -1170 16870 -1136 16904
rect -978 16870 -894 16904
rect -720 16870 -636 16904
rect -478 16870 -444 16904
rect -1270 16820 -1236 16854
rect -378 16843 -344 17541
rect -378 16820 -344 16843
rect -1270 16786 -1210 16820
rect -1210 16786 -404 16820
rect -404 16786 -344 16820
rect -209 17587 -149 17621
rect -149 17587 8627 17621
rect 8627 17587 8687 17621
rect -209 17539 -175 17587
rect -209 15985 -175 17539
rect -92 17502 -58 17536
rect 5332 17502 7316 17536
rect 8536 17502 8570 17536
rect -92 17276 -58 17452
rect -4 17276 30 17452
rect 108 17276 142 17452
rect 4166 17276 4200 17452
rect 4278 17276 4312 17452
rect 8336 17276 8370 17452
rect 8448 17276 8482 17452
rect 8536 17276 8570 17452
rect 8653 17539 8687 17587
rect -92 17108 -58 17142
rect 8536 17108 8570 17142
rect -92 16882 -58 17058
rect -4 16882 30 17058
rect 108 16882 142 17058
rect 4166 16882 4200 17058
rect 4278 16882 4312 17058
rect 8336 16882 8370 17058
rect 8448 16882 8482 17058
rect 8536 16882 8570 17058
rect -92 16488 -58 16664
rect -4 16488 30 16664
rect 108 16488 142 16664
rect 4166 16488 4200 16664
rect 4278 16488 4312 16664
rect 8336 16488 8370 16664
rect 8448 16488 8482 16664
rect 8536 16488 8570 16664
rect -92 16404 -58 16438
rect 8536 16404 8570 16438
rect -92 16094 -58 16270
rect -4 16094 30 16270
rect 108 16094 142 16270
rect 4166 16094 4200 16270
rect 4278 16094 4312 16270
rect 8336 16094 8370 16270
rect 8448 16094 8482 16270
rect 8536 16094 8570 16270
rect -92 16010 -58 16044
rect 1162 16010 3146 16044
rect 8536 16010 8570 16044
rect -209 15959 -175 15985
rect 8653 15985 8687 17539
rect 8653 15959 8687 15985
rect -209 15925 -149 15959
rect -149 15925 8627 15959
rect 8627 15925 8687 15959
rect -3030 15692 -2996 15718
rect -7670 15658 -7585 15692
rect -7585 15658 -3081 15692
rect -3081 15658 -2996 15692
rect -1220 15829 -1160 15863
rect -1160 15829 2568 15863
rect 2568 15829 2628 15863
rect -1220 15803 -1186 15829
rect -12483 15558 -12423 15592
rect -12423 15558 -7986 15592
rect -7986 15558 -7926 15592
rect -12483 15532 -12449 15558
rect -12483 14722 -12449 15532
rect -7960 15532 -7926 15558
rect -11726 15471 -10742 15505
rect -9668 15471 -8684 15505
rect -12368 15236 -12334 15412
rect -12280 15236 -12246 15412
rect -10222 15236 -10188 15412
rect -8164 15236 -8130 15412
rect -8076 15236 -8042 15412
rect -12368 15110 -12334 15144
rect -8076 15110 -8042 15144
rect -12368 14842 -12334 15018
rect -12280 14842 -12246 15018
rect -10222 14842 -10188 15018
rect -8164 14842 -8130 15018
rect -8076 14842 -8042 15018
rect -11726 14749 -10742 14783
rect -9668 14749 -8684 14783
rect -12483 14696 -12449 14722
rect -7960 14722 -7926 15532
rect -7562 15543 -7502 15577
rect -7502 15543 -3096 15577
rect -3096 15543 -3036 15577
rect -7562 15517 -7528 15543
rect -7562 14785 -7528 15517
rect -3070 15517 -3036 15543
rect -7462 15301 -7428 15477
rect -7374 15301 -7340 15477
rect -5316 15301 -5282 15477
rect -3258 15301 -3224 15477
rect -3170 15301 -3136 15477
rect -7462 15207 -7428 15241
rect -6820 15208 -5836 15242
rect -4762 15208 -3778 15242
rect -3170 15208 -3136 15242
rect -7462 15060 -7428 15094
rect -6820 15060 -5836 15094
rect -4762 15060 -3778 15094
rect -3170 15060 -3136 15094
rect -7462 14825 -7428 15001
rect -7374 14825 -7340 15001
rect -5316 14825 -5282 15001
rect -3258 14825 -3224 15001
rect -3170 14825 -3136 15001
rect -7562 14759 -7528 14785
rect -3070 14785 -3036 15517
rect -3070 14759 -3036 14785
rect -7562 14725 -7502 14759
rect -7502 14725 -3096 14759
rect -3096 14725 -3036 14759
rect -1220 14763 -1186 15803
rect 2594 15803 2628 15829
rect -1062 15679 -665 15717
rect 237 15679 634 15717
rect 774 15679 1171 15717
rect 2073 15679 2470 15717
rect -1062 15513 -665 15551
rect 237 15513 634 15551
rect 774 15513 1171 15551
rect 2073 15513 2470 15551
rect -1062 15347 -665 15385
rect 237 15347 634 15385
rect 774 15347 1171 15385
rect 2073 15347 2470 15385
rect -1062 15181 -665 15219
rect 237 15181 634 15219
rect 774 15181 1171 15219
rect 2073 15181 2470 15219
rect -1062 15015 -665 15053
rect 237 15015 634 15053
rect 774 15015 1171 15053
rect 2073 15015 2470 15053
rect -1062 14849 -665 14887
rect 237 14849 634 14887
rect 774 14849 1171 14887
rect 2073 14849 2470 14887
rect -1220 14737 -1186 14763
rect 2594 14763 2628 15803
rect 2865 15744 2927 15778
rect 2927 15744 8625 15778
rect 8625 15744 8687 15778
rect 2865 15703 2899 15744
rect 2865 14861 2899 15703
rect 8653 15703 8687 15744
rect 3805 15584 5089 15618
rect 6463 15584 7747 15618
rect 3013 15378 3047 15534
rect 3101 15378 3135 15534
rect 5759 15378 5793 15534
rect 8417 15378 8451 15534
rect 8505 15378 8539 15534
rect 3013 15294 3047 15328
rect 3805 15294 5089 15328
rect 6463 15294 7747 15328
rect 8505 15294 8539 15328
rect 3013 15152 3047 15186
rect 3805 15152 5089 15186
rect 6463 15152 7747 15186
rect 8505 15152 8539 15186
rect 3013 14946 3047 15102
rect 3101 14946 3135 15102
rect 5759 14946 5793 15102
rect 8417 14946 8451 15102
rect 8505 14946 8539 15102
rect 2865 14820 2899 14861
rect 8653 14861 8687 15703
rect 8653 14820 8687 14861
rect 2865 14786 2927 14820
rect 2927 14786 8625 14820
rect 8625 14786 8687 14820
rect 2594 14737 2628 14763
rect -7960 14696 -7926 14722
rect -1220 14703 -1160 14737
rect -1160 14703 2568 14737
rect 2568 14703 2628 14737
rect -12483 14662 -12423 14696
rect -12423 14662 -7986 14696
rect -7986 14662 -7926 14696
rect 854 12216 1022 12250
rect 1112 12216 1280 12250
rect 704 11390 738 12166
rect 792 11390 826 12166
rect 1050 11390 1084 12166
rect 1308 11390 1342 12166
rect 1396 11390 1430 12166
rect 704 11264 738 11298
rect 1396 11264 1430 11298
rect 604 10291 638 10471
rect 704 10396 738 11172
rect 792 10396 826 11172
rect 1050 10396 1084 11172
rect 1308 10396 1342 11172
rect 1396 10396 1430 11172
rect 854 10312 1022 10346
rect 1112 10312 1280 10346
rect 1746 12216 1914 12250
rect 2004 12216 2172 12250
rect 1596 11390 1630 12166
rect 1684 11390 1718 12166
rect 1942 11390 1976 12166
rect 2200 11390 2234 12166
rect 2288 11390 2322 12166
rect 1596 11264 1630 11298
rect 2288 11264 2322 11298
rect 1596 10396 1630 11172
rect 1684 10396 1718 11172
rect 1942 10396 1976 11172
rect 2200 10396 2234 11172
rect 2288 10396 2322 11172
rect 1746 10312 1914 10346
rect 2004 10312 2172 10346
rect 2638 12216 2806 12250
rect 2896 12216 3064 12250
rect 2488 11390 2522 12166
rect 2576 11390 2610 12166
rect 2834 11390 2868 12166
rect 3092 11390 3126 12166
rect 3180 11390 3214 12166
rect 2488 11264 2522 11298
rect 3180 11264 3214 11298
rect 2488 10396 2522 11172
rect 2576 10396 2610 11172
rect 2834 10396 2868 11172
rect 3092 10396 3126 11172
rect 3180 10396 3214 11172
rect 2638 10312 2806 10346
rect 2896 10312 3064 10346
rect 3530 12216 3698 12250
rect 3788 12216 3956 12250
rect 3380 11390 3414 12166
rect 3468 11390 3502 12166
rect 3726 11390 3760 12166
rect 3984 11390 4018 12166
rect 4072 11390 4106 12166
rect 3380 11264 3414 11298
rect 4072 11264 4106 11298
rect 3380 10396 3414 11172
rect 3468 10396 3502 11172
rect 3726 10396 3760 11172
rect 3984 10396 4018 11172
rect 4072 10396 4106 11172
rect 3530 10312 3698 10346
rect 3788 10312 3956 10346
rect 4344 12167 4378 12201
rect 4428 12167 4604 12201
rect 4428 12079 4604 12113
rect 4654 11883 4688 12051
rect 4428 11821 4604 11855
rect 4654 11625 4688 11793
rect 4428 11563 4604 11597
rect 4344 11475 4378 11509
rect 4428 11475 4604 11509
rect 4344 11053 4378 11087
rect 4428 11053 4604 11087
rect 4428 10965 4604 10999
rect 4654 10769 4688 10937
rect 4428 10707 4604 10741
rect 4654 10511 4688 10679
rect 4428 10449 4604 10483
rect 4344 10361 4378 10395
rect 4428 10361 4604 10395
rect 5001 11778 5377 11812
rect 5469 11778 5503 11812
rect 5595 11778 5971 11812
rect 5001 11690 5377 11724
rect 5595 11690 5971 11724
rect 4908 11386 4942 11570
rect 6030 11386 6064 11570
rect 5001 11232 5377 11266
rect 5595 11232 5971 11266
rect 4908 10928 4942 11112
rect 6030 10928 6064 11112
rect 5001 10774 5377 10808
rect 5595 10774 5971 10808
rect 5001 10686 5377 10720
rect 5469 10686 5503 10720
rect 5595 10686 5971 10720
rect 757 9973 937 10007
rect 713 8016 719 8022
rect 719 8016 747 8022
rect 713 7988 747 8016
rect 813 7988 847 8022
rect 913 7988 947 8022
rect 1013 8016 1045 8022
rect 1045 8016 1047 8022
rect 1113 8016 1135 8022
rect 1135 8016 1147 8022
rect 1213 8016 1225 8022
rect 1225 8016 1247 8022
rect 1013 7988 1047 8016
rect 1113 7988 1147 8016
rect 1213 7988 1247 8016
rect 713 7888 747 7922
rect 813 7888 847 7922
rect 913 7888 947 7922
rect 1013 7888 1047 7922
rect 1113 7888 1147 7922
rect 1213 7888 1247 7922
rect 713 7788 747 7822
rect 813 7788 847 7822
rect 913 7788 947 7822
rect 1013 7788 1047 7822
rect 1113 7788 1147 7822
rect 1213 7788 1247 7822
rect 713 7690 747 7722
rect 713 7688 719 7690
rect 719 7688 747 7690
rect 813 7688 847 7722
rect 913 7688 947 7722
rect 1013 7690 1047 7722
rect 1113 7690 1147 7722
rect 1213 7690 1247 7722
rect 1013 7688 1045 7690
rect 1045 7688 1047 7690
rect 1113 7688 1135 7690
rect 1135 7688 1147 7690
rect 1213 7688 1225 7690
rect 1225 7688 1247 7690
rect 713 7600 747 7622
rect 713 7588 719 7600
rect 719 7588 747 7600
rect 813 7588 847 7622
rect 913 7588 947 7622
rect 1013 7600 1047 7622
rect 1113 7600 1147 7622
rect 1213 7600 1247 7622
rect 1013 7588 1045 7600
rect 1045 7588 1047 7600
rect 1113 7588 1135 7600
rect 1135 7588 1147 7600
rect 1213 7588 1225 7600
rect 1225 7588 1247 7600
rect 713 7510 747 7522
rect 713 7488 719 7510
rect 719 7488 747 7510
rect 813 7488 847 7522
rect 913 7488 947 7522
rect 1013 7510 1047 7522
rect 1113 7510 1147 7522
rect 1213 7510 1247 7522
rect 1013 7488 1045 7510
rect 1045 7488 1047 7510
rect 1113 7488 1135 7510
rect 1135 7488 1147 7510
rect 1213 7488 1225 7510
rect 1225 7488 1247 7510
rect 1382 7281 1454 7353
rect 1518 7338 1551 7353
rect 1551 7338 1585 7353
rect 1585 7338 1617 7353
rect 1518 7282 1617 7338
rect 1518 7281 1551 7282
rect 1551 7281 1585 7282
rect 1585 7281 1617 7282
rect 1382 7186 1454 7217
rect 1382 7152 1411 7186
rect 1411 7152 1454 7186
rect 1382 7118 1454 7152
rect 2101 8016 2107 8022
rect 2107 8016 2135 8022
rect 2101 7988 2135 8016
rect 2201 7988 2235 8022
rect 2301 7988 2335 8022
rect 2401 8016 2433 8022
rect 2433 8016 2435 8022
rect 2501 8016 2523 8022
rect 2523 8016 2535 8022
rect 2601 8016 2613 8022
rect 2613 8016 2635 8022
rect 2401 7988 2435 8016
rect 2501 7988 2535 8016
rect 2601 7988 2635 8016
rect 2101 7888 2135 7922
rect 2201 7888 2235 7922
rect 2301 7888 2335 7922
rect 2401 7888 2435 7922
rect 2501 7888 2535 7922
rect 2601 7888 2635 7922
rect 2101 7788 2135 7822
rect 2201 7788 2235 7822
rect 2301 7788 2335 7822
rect 2401 7788 2435 7822
rect 2501 7788 2535 7822
rect 2601 7788 2635 7822
rect 2101 7690 2135 7722
rect 2101 7688 2107 7690
rect 2107 7688 2135 7690
rect 2201 7688 2235 7722
rect 2301 7688 2335 7722
rect 2401 7690 2435 7722
rect 2501 7690 2535 7722
rect 2601 7690 2635 7722
rect 2401 7688 2433 7690
rect 2433 7688 2435 7690
rect 2501 7688 2523 7690
rect 2523 7688 2535 7690
rect 2601 7688 2613 7690
rect 2613 7688 2635 7690
rect 2101 7600 2135 7622
rect 2101 7588 2107 7600
rect 2107 7588 2135 7600
rect 2201 7588 2235 7622
rect 2301 7588 2335 7622
rect 2401 7600 2435 7622
rect 2501 7600 2535 7622
rect 2601 7600 2635 7622
rect 2401 7588 2433 7600
rect 2433 7588 2435 7600
rect 2501 7588 2523 7600
rect 2523 7588 2535 7600
rect 2601 7588 2613 7600
rect 2613 7588 2635 7600
rect 2101 7510 2135 7522
rect 2101 7488 2107 7510
rect 2107 7488 2135 7510
rect 2201 7488 2235 7522
rect 2301 7488 2335 7522
rect 2401 7510 2435 7522
rect 2501 7510 2535 7522
rect 2601 7510 2635 7522
rect 2401 7488 2433 7510
rect 2433 7488 2435 7510
rect 2501 7488 2523 7510
rect 2523 7488 2535 7510
rect 2601 7488 2613 7510
rect 2613 7488 2635 7510
rect 2770 7281 2842 7353
rect 2906 7338 2939 7353
rect 2939 7338 2973 7353
rect 2973 7338 3005 7353
rect 2906 7282 3005 7338
rect 2906 7281 2939 7282
rect 2939 7281 2973 7282
rect 2973 7281 3005 7282
rect 3105 7338 3140 7353
rect 3140 7338 3174 7353
rect 3174 7338 3204 7353
rect 3105 7282 3204 7338
rect 3105 7281 3140 7282
rect 3140 7281 3174 7282
rect 3174 7281 3204 7282
rect 3489 8016 3495 8022
rect 3495 8016 3523 8022
rect 3489 7988 3523 8016
rect 3589 7988 3623 8022
rect 3689 7988 3723 8022
rect 3789 8016 3821 8022
rect 3821 8016 3823 8022
rect 3889 8016 3911 8022
rect 3911 8016 3923 8022
rect 3989 8016 4001 8022
rect 4001 8016 4023 8022
rect 3789 7988 3823 8016
rect 3889 7988 3923 8016
rect 3989 7988 4023 8016
rect 3489 7888 3523 7922
rect 3589 7888 3623 7922
rect 3689 7888 3723 7922
rect 3789 7888 3823 7922
rect 3889 7888 3923 7922
rect 3989 7888 4023 7922
rect 3489 7788 3523 7822
rect 3589 7788 3623 7822
rect 3689 7788 3723 7822
rect 3789 7788 3823 7822
rect 3889 7788 3923 7822
rect 3989 7788 4023 7822
rect 3489 7690 3523 7722
rect 3489 7688 3495 7690
rect 3495 7688 3523 7690
rect 3589 7688 3623 7722
rect 3689 7688 3723 7722
rect 3789 7690 3823 7722
rect 3889 7690 3923 7722
rect 3989 7690 4023 7722
rect 3789 7688 3821 7690
rect 3821 7688 3823 7690
rect 3889 7688 3911 7690
rect 3911 7688 3923 7690
rect 3989 7688 4001 7690
rect 4001 7688 4023 7690
rect 3489 7600 3523 7622
rect 3489 7588 3495 7600
rect 3495 7588 3523 7600
rect 3589 7588 3623 7622
rect 3689 7588 3723 7622
rect 3789 7600 3823 7622
rect 3889 7600 3923 7622
rect 3989 7600 4023 7622
rect 3789 7588 3821 7600
rect 3821 7588 3823 7600
rect 3889 7588 3911 7600
rect 3911 7588 3923 7600
rect 3989 7588 4001 7600
rect 4001 7588 4023 7600
rect 3489 7510 3523 7522
rect 3489 7488 3495 7510
rect 3495 7488 3523 7510
rect 3589 7488 3623 7522
rect 3689 7488 3723 7522
rect 3789 7510 3823 7522
rect 3889 7510 3923 7522
rect 3989 7510 4023 7522
rect 3789 7488 3821 7510
rect 3821 7488 3823 7510
rect 3889 7488 3911 7510
rect 3911 7488 3923 7510
rect 3989 7488 4001 7510
rect 4001 7488 4023 7510
rect 3268 7281 3340 7353
rect 4158 7281 4230 7353
rect 4294 7338 4327 7353
rect 4327 7338 4361 7353
rect 4361 7338 4393 7353
rect 4294 7282 4393 7338
rect 4294 7281 4327 7282
rect 4327 7281 4361 7282
rect 4361 7281 4393 7282
rect 4493 7338 4528 7353
rect 4528 7338 4562 7353
rect 4562 7338 4592 7353
rect 4493 7282 4592 7338
rect 4493 7281 4528 7282
rect 4528 7281 4562 7282
rect 4562 7281 4592 7282
rect 4877 8016 4883 8022
rect 4883 8016 4911 8022
rect 4877 7988 4911 8016
rect 4977 7988 5011 8022
rect 5077 7988 5111 8022
rect 5177 8016 5209 8022
rect 5209 8016 5211 8022
rect 5277 8016 5299 8022
rect 5299 8016 5311 8022
rect 5377 8016 5389 8022
rect 5389 8016 5411 8022
rect 5177 7988 5211 8016
rect 5277 7988 5311 8016
rect 5377 7988 5411 8016
rect 4877 7888 4911 7922
rect 4977 7888 5011 7922
rect 5077 7888 5111 7922
rect 5177 7888 5211 7922
rect 5277 7888 5311 7922
rect 5377 7888 5411 7922
rect 4877 7788 4911 7822
rect 4977 7788 5011 7822
rect 5077 7788 5111 7822
rect 5177 7788 5211 7822
rect 5277 7788 5311 7822
rect 5377 7788 5411 7822
rect 4877 7690 4911 7722
rect 4877 7688 4883 7690
rect 4883 7688 4911 7690
rect 4977 7688 5011 7722
rect 5077 7688 5111 7722
rect 5177 7690 5211 7722
rect 5277 7690 5311 7722
rect 5377 7690 5411 7722
rect 5177 7688 5209 7690
rect 5209 7688 5211 7690
rect 5277 7688 5299 7690
rect 5299 7688 5311 7690
rect 5377 7688 5389 7690
rect 5389 7688 5411 7690
rect 4877 7600 4911 7622
rect 4877 7588 4883 7600
rect 4883 7588 4911 7600
rect 4977 7588 5011 7622
rect 5077 7588 5111 7622
rect 5177 7600 5211 7622
rect 5277 7600 5311 7622
rect 5377 7600 5411 7622
rect 5177 7588 5209 7600
rect 5209 7588 5211 7600
rect 5277 7588 5299 7600
rect 5299 7588 5311 7600
rect 5377 7588 5389 7600
rect 5389 7588 5411 7600
rect 4877 7510 4911 7522
rect 4877 7488 4883 7510
rect 4883 7488 4911 7510
rect 4977 7488 5011 7522
rect 5077 7488 5111 7522
rect 5177 7510 5211 7522
rect 5277 7510 5311 7522
rect 5377 7510 5411 7522
rect 5177 7488 5209 7510
rect 5209 7488 5211 7510
rect 5277 7488 5299 7510
rect 5299 7488 5311 7510
rect 5377 7488 5389 7510
rect 5389 7488 5411 7510
rect 4656 7281 4728 7353
rect 5546 7281 5618 7353
rect 5682 7338 5715 7353
rect 5715 7338 5749 7353
rect 5749 7338 5781 7353
rect 5682 7282 5781 7338
rect 5682 7281 5715 7282
rect 5715 7281 5749 7282
rect 5749 7281 5781 7282
rect 5881 7338 5916 7353
rect 5916 7338 5950 7353
rect 5950 7338 5980 7353
rect 5881 7282 5980 7338
rect 5881 7281 5916 7282
rect 5916 7281 5950 7282
rect 5950 7281 5980 7282
rect 6265 8016 6271 8022
rect 6271 8016 6299 8022
rect 6265 7988 6299 8016
rect 6365 7988 6399 8022
rect 6465 7988 6499 8022
rect 6565 8016 6597 8022
rect 6597 8016 6599 8022
rect 6665 8016 6687 8022
rect 6687 8016 6699 8022
rect 6765 8016 6777 8022
rect 6777 8016 6799 8022
rect 6565 7988 6599 8016
rect 6665 7988 6699 8016
rect 6765 7988 6799 8016
rect 6265 7888 6299 7922
rect 6365 7888 6399 7922
rect 6465 7888 6499 7922
rect 6565 7888 6599 7922
rect 6665 7888 6699 7922
rect 6765 7888 6799 7922
rect 6265 7788 6299 7822
rect 6365 7788 6399 7822
rect 6465 7788 6499 7822
rect 6565 7788 6599 7822
rect 6665 7788 6699 7822
rect 6765 7788 6799 7822
rect 6265 7690 6299 7722
rect 6265 7688 6271 7690
rect 6271 7688 6299 7690
rect 6365 7688 6399 7722
rect 6465 7688 6499 7722
rect 6565 7690 6599 7722
rect 6665 7690 6699 7722
rect 6765 7690 6799 7722
rect 6565 7688 6597 7690
rect 6597 7688 6599 7690
rect 6665 7688 6687 7690
rect 6687 7688 6699 7690
rect 6765 7688 6777 7690
rect 6777 7688 6799 7690
rect 6265 7600 6299 7622
rect 6265 7588 6271 7600
rect 6271 7588 6299 7600
rect 6365 7588 6399 7622
rect 6465 7588 6499 7622
rect 6565 7600 6599 7622
rect 6665 7600 6699 7622
rect 6765 7600 6799 7622
rect 6565 7588 6597 7600
rect 6597 7588 6599 7600
rect 6665 7588 6687 7600
rect 6687 7588 6699 7600
rect 6765 7588 6777 7600
rect 6777 7588 6799 7600
rect 6265 7510 6299 7522
rect 6265 7488 6271 7510
rect 6271 7488 6299 7510
rect 6365 7488 6399 7522
rect 6465 7488 6499 7522
rect 6565 7510 6599 7522
rect 6665 7510 6699 7522
rect 6765 7510 6799 7522
rect 6565 7488 6597 7510
rect 6597 7488 6599 7510
rect 6665 7488 6687 7510
rect 6687 7488 6699 7510
rect 6765 7488 6777 7510
rect 6777 7488 6799 7510
rect 6044 7281 6116 7353
rect 6044 7186 6116 7217
rect 6044 7152 6063 7186
rect 6063 7152 6116 7186
rect 6044 7118 6116 7152
rect 1382 6985 1454 7018
rect 1382 6951 1411 6985
rect 1411 6951 1454 6985
rect 1382 6919 1454 6951
rect 1382 6783 1454 6855
rect 713 6628 719 6634
rect 719 6628 747 6634
rect 713 6600 747 6628
rect 813 6600 847 6634
rect 913 6600 947 6634
rect 1013 6628 1045 6634
rect 1045 6628 1047 6634
rect 1113 6628 1135 6634
rect 1135 6628 1147 6634
rect 1213 6628 1225 6634
rect 1225 6628 1247 6634
rect 1013 6600 1047 6628
rect 1113 6600 1147 6628
rect 1213 6600 1247 6628
rect 713 6500 747 6534
rect 813 6500 847 6534
rect 913 6500 947 6534
rect 1013 6500 1047 6534
rect 1113 6500 1147 6534
rect 1213 6500 1247 6534
rect 713 6400 747 6434
rect 813 6400 847 6434
rect 913 6400 947 6434
rect 1013 6400 1047 6434
rect 1113 6400 1147 6434
rect 1213 6400 1247 6434
rect 713 6302 747 6334
rect 713 6300 719 6302
rect 719 6300 747 6302
rect 813 6300 847 6334
rect 913 6300 947 6334
rect 1013 6302 1047 6334
rect 1113 6302 1147 6334
rect 1213 6302 1247 6334
rect 1013 6300 1045 6302
rect 1045 6300 1047 6302
rect 1113 6300 1135 6302
rect 1135 6300 1147 6302
rect 1213 6300 1225 6302
rect 1225 6300 1247 6302
rect 713 6212 747 6234
rect 713 6200 719 6212
rect 719 6200 747 6212
rect 813 6200 847 6234
rect 913 6200 947 6234
rect 1013 6212 1047 6234
rect 1113 6212 1147 6234
rect 1213 6212 1247 6234
rect 1013 6200 1045 6212
rect 1045 6200 1047 6212
rect 1113 6200 1135 6212
rect 1135 6200 1147 6212
rect 1213 6200 1225 6212
rect 1225 6200 1247 6212
rect 713 6122 747 6134
rect 713 6100 719 6122
rect 719 6100 747 6122
rect 813 6100 847 6134
rect 913 6100 947 6134
rect 1013 6122 1047 6134
rect 1113 6122 1147 6134
rect 1213 6122 1247 6134
rect 1013 6100 1045 6122
rect 1045 6100 1047 6122
rect 1113 6100 1135 6122
rect 1135 6100 1147 6122
rect 1213 6100 1225 6122
rect 1225 6100 1247 6122
rect 1382 5893 1454 5965
rect 1382 5798 1454 5829
rect 1382 5764 1411 5798
rect 1411 5764 1454 5798
rect 1382 5730 1454 5764
rect 2101 6628 2107 6634
rect 2107 6628 2135 6634
rect 2101 6600 2135 6628
rect 2201 6600 2235 6634
rect 2301 6600 2335 6634
rect 2401 6628 2433 6634
rect 2433 6628 2435 6634
rect 2501 6628 2523 6634
rect 2523 6628 2535 6634
rect 2601 6628 2613 6634
rect 2613 6628 2635 6634
rect 2401 6600 2435 6628
rect 2501 6600 2535 6628
rect 2601 6600 2635 6628
rect 2101 6500 2135 6534
rect 2201 6500 2235 6534
rect 2301 6500 2335 6534
rect 2401 6500 2435 6534
rect 2501 6500 2535 6534
rect 2601 6500 2635 6534
rect 2101 6400 2135 6434
rect 2201 6400 2235 6434
rect 2301 6400 2335 6434
rect 2401 6400 2435 6434
rect 2501 6400 2535 6434
rect 2601 6400 2635 6434
rect 2101 6302 2135 6334
rect 2101 6300 2107 6302
rect 2107 6300 2135 6302
rect 2201 6300 2235 6334
rect 2301 6300 2335 6334
rect 2401 6302 2435 6334
rect 2501 6302 2535 6334
rect 2601 6302 2635 6334
rect 2401 6300 2433 6302
rect 2433 6300 2435 6302
rect 2501 6300 2523 6302
rect 2523 6300 2535 6302
rect 2601 6300 2613 6302
rect 2613 6300 2635 6302
rect 2101 6212 2135 6234
rect 2101 6200 2107 6212
rect 2107 6200 2135 6212
rect 2201 6200 2235 6234
rect 2301 6200 2335 6234
rect 2401 6212 2435 6234
rect 2501 6212 2535 6234
rect 2601 6212 2635 6234
rect 2401 6200 2433 6212
rect 2433 6200 2435 6212
rect 2501 6200 2523 6212
rect 2523 6200 2535 6212
rect 2601 6200 2613 6212
rect 2613 6200 2635 6212
rect 2101 6122 2135 6134
rect 2101 6100 2107 6122
rect 2107 6100 2135 6122
rect 2201 6100 2235 6134
rect 2301 6100 2335 6134
rect 2401 6122 2435 6134
rect 2501 6122 2535 6134
rect 2601 6122 2635 6134
rect 2401 6100 2433 6122
rect 2433 6100 2435 6122
rect 2501 6100 2523 6122
rect 2523 6100 2535 6122
rect 2601 6100 2613 6122
rect 2613 6100 2635 6122
rect 2770 5893 2842 5965
rect 2906 5950 2939 5965
rect 2939 5950 2973 5965
rect 2973 5950 3005 5965
rect 2906 5894 3005 5950
rect 2906 5893 2939 5894
rect 2939 5893 2973 5894
rect 2973 5893 3005 5894
rect 2770 5798 2842 5829
rect 2770 5764 2799 5798
rect 2799 5764 2842 5798
rect 2770 5730 2842 5764
rect 3105 5950 3140 5965
rect 3140 5950 3174 5965
rect 3174 5950 3204 5965
rect 3105 5894 3204 5950
rect 3105 5893 3140 5894
rect 3140 5893 3174 5894
rect 3174 5893 3204 5894
rect 3489 6628 3495 6634
rect 3495 6628 3523 6634
rect 3489 6600 3523 6628
rect 3589 6600 3623 6634
rect 3689 6600 3723 6634
rect 3789 6628 3821 6634
rect 3821 6628 3823 6634
rect 3889 6628 3911 6634
rect 3911 6628 3923 6634
rect 3989 6628 4001 6634
rect 4001 6628 4023 6634
rect 3789 6600 3823 6628
rect 3889 6600 3923 6628
rect 3989 6600 4023 6628
rect 3489 6500 3523 6534
rect 3589 6500 3623 6534
rect 3689 6500 3723 6534
rect 3789 6500 3823 6534
rect 3889 6500 3923 6534
rect 3989 6500 4023 6534
rect 3489 6400 3523 6434
rect 3589 6400 3623 6434
rect 3689 6400 3723 6434
rect 3789 6400 3823 6434
rect 3889 6400 3923 6434
rect 3989 6400 4023 6434
rect 3489 6302 3523 6334
rect 3489 6300 3495 6302
rect 3495 6300 3523 6302
rect 3589 6300 3623 6334
rect 3689 6300 3723 6334
rect 3789 6302 3823 6334
rect 3889 6302 3923 6334
rect 3989 6302 4023 6334
rect 3789 6300 3821 6302
rect 3821 6300 3823 6302
rect 3889 6300 3911 6302
rect 3911 6300 3923 6302
rect 3989 6300 4001 6302
rect 4001 6300 4023 6302
rect 3489 6212 3523 6234
rect 3489 6200 3495 6212
rect 3495 6200 3523 6212
rect 3589 6200 3623 6234
rect 3689 6200 3723 6234
rect 3789 6212 3823 6234
rect 3889 6212 3923 6234
rect 3989 6212 4023 6234
rect 3789 6200 3821 6212
rect 3821 6200 3823 6212
rect 3889 6200 3911 6212
rect 3911 6200 3923 6212
rect 3989 6200 4001 6212
rect 4001 6200 4023 6212
rect 3489 6122 3523 6134
rect 3489 6100 3495 6122
rect 3495 6100 3523 6122
rect 3589 6100 3623 6134
rect 3689 6100 3723 6134
rect 3789 6122 3823 6134
rect 3889 6122 3923 6134
rect 3989 6122 4023 6134
rect 3789 6100 3821 6122
rect 3821 6100 3823 6122
rect 3889 6100 3911 6122
rect 3911 6100 3923 6122
rect 3989 6100 4001 6122
rect 4001 6100 4023 6122
rect 3268 5893 3340 5965
rect 4158 5893 4230 5965
rect 4294 5950 4327 5965
rect 4327 5950 4361 5965
rect 4361 5950 4393 5965
rect 4294 5894 4393 5950
rect 4294 5893 4327 5894
rect 4327 5893 4361 5894
rect 4361 5893 4393 5894
rect 4493 5950 4528 5965
rect 4528 5950 4562 5965
rect 4562 5950 4592 5965
rect 4493 5894 4592 5950
rect 4493 5893 4528 5894
rect 4528 5893 4562 5894
rect 4562 5893 4592 5894
rect 4877 6628 4883 6634
rect 4883 6628 4911 6634
rect 4877 6600 4911 6628
rect 4977 6600 5011 6634
rect 5077 6600 5111 6634
rect 5177 6628 5209 6634
rect 5209 6628 5211 6634
rect 5277 6628 5299 6634
rect 5299 6628 5311 6634
rect 5377 6628 5389 6634
rect 5389 6628 5411 6634
rect 5177 6600 5211 6628
rect 5277 6600 5311 6628
rect 5377 6600 5411 6628
rect 4877 6500 4911 6534
rect 4977 6500 5011 6534
rect 5077 6500 5111 6534
rect 5177 6500 5211 6534
rect 5277 6500 5311 6534
rect 5377 6500 5411 6534
rect 4877 6400 4911 6434
rect 4977 6400 5011 6434
rect 5077 6400 5111 6434
rect 5177 6400 5211 6434
rect 5277 6400 5311 6434
rect 5377 6400 5411 6434
rect 4877 6302 4911 6334
rect 4877 6300 4883 6302
rect 4883 6300 4911 6302
rect 4977 6300 5011 6334
rect 5077 6300 5111 6334
rect 5177 6302 5211 6334
rect 5277 6302 5311 6334
rect 5377 6302 5411 6334
rect 5177 6300 5209 6302
rect 5209 6300 5211 6302
rect 5277 6300 5299 6302
rect 5299 6300 5311 6302
rect 5377 6300 5389 6302
rect 5389 6300 5411 6302
rect 4877 6212 4911 6234
rect 4877 6200 4883 6212
rect 4883 6200 4911 6212
rect 4977 6200 5011 6234
rect 5077 6200 5111 6234
rect 5177 6212 5211 6234
rect 5277 6212 5311 6234
rect 5377 6212 5411 6234
rect 5177 6200 5209 6212
rect 5209 6200 5211 6212
rect 5277 6200 5299 6212
rect 5299 6200 5311 6212
rect 5377 6200 5389 6212
rect 5389 6200 5411 6212
rect 4877 6122 4911 6134
rect 4877 6100 4883 6122
rect 4883 6100 4911 6122
rect 4977 6100 5011 6134
rect 5077 6100 5111 6134
rect 5177 6122 5211 6134
rect 5277 6122 5311 6134
rect 5377 6122 5411 6134
rect 5177 6100 5209 6122
rect 5209 6100 5211 6122
rect 5277 6100 5299 6122
rect 5299 6100 5311 6122
rect 5377 6100 5389 6122
rect 5389 6100 5411 6122
rect 4656 5893 4728 5965
rect 4656 5798 4728 5829
rect 4656 5764 4675 5798
rect 4675 5764 4728 5798
rect 4656 5730 4728 5764
rect 6044 6985 6116 7018
rect 6044 6951 6063 6985
rect 6063 6951 6116 6985
rect 6044 6919 6116 6951
rect 6044 6783 6116 6855
rect 6265 6628 6271 6634
rect 6271 6628 6299 6634
rect 6265 6600 6299 6628
rect 6365 6600 6399 6634
rect 6465 6600 6499 6634
rect 6565 6628 6597 6634
rect 6597 6628 6599 6634
rect 6665 6628 6687 6634
rect 6687 6628 6699 6634
rect 6765 6628 6777 6634
rect 6777 6628 6799 6634
rect 6565 6600 6599 6628
rect 6665 6600 6699 6628
rect 6765 6600 6799 6628
rect 6265 6500 6299 6534
rect 6365 6500 6399 6534
rect 6465 6500 6499 6534
rect 6565 6500 6599 6534
rect 6665 6500 6699 6534
rect 6765 6500 6799 6534
rect 6265 6400 6299 6434
rect 6365 6400 6399 6434
rect 6465 6400 6499 6434
rect 6565 6400 6599 6434
rect 6665 6400 6699 6434
rect 6765 6400 6799 6434
rect 6265 6302 6299 6334
rect 6265 6300 6271 6302
rect 6271 6300 6299 6302
rect 6365 6300 6399 6334
rect 6465 6300 6499 6334
rect 6565 6302 6599 6334
rect 6665 6302 6699 6334
rect 6765 6302 6799 6334
rect 6565 6300 6597 6302
rect 6597 6300 6599 6302
rect 6665 6300 6687 6302
rect 6687 6300 6699 6302
rect 6765 6300 6777 6302
rect 6777 6300 6799 6302
rect 6265 6212 6299 6234
rect 6265 6200 6271 6212
rect 6271 6200 6299 6212
rect 6365 6200 6399 6234
rect 6465 6200 6499 6234
rect 6565 6212 6599 6234
rect 6665 6212 6699 6234
rect 6765 6212 6799 6234
rect 6565 6200 6597 6212
rect 6597 6200 6599 6212
rect 6665 6200 6687 6212
rect 6687 6200 6699 6212
rect 6765 6200 6777 6212
rect 6777 6200 6799 6212
rect 6265 6122 6299 6134
rect 6265 6100 6271 6122
rect 6271 6100 6299 6122
rect 6365 6100 6399 6134
rect 6465 6100 6499 6134
rect 6565 6122 6599 6134
rect 6665 6122 6699 6134
rect 6765 6122 6799 6134
rect 6565 6100 6597 6122
rect 6597 6100 6599 6122
rect 6665 6100 6687 6122
rect 6687 6100 6699 6122
rect 6765 6100 6777 6122
rect 6777 6100 6799 6122
rect 6044 5893 6116 5965
rect 6044 5798 6116 5829
rect 6044 5764 6063 5798
rect 6063 5764 6116 5798
rect 6044 5730 6116 5764
rect 1382 5597 1454 5630
rect 1382 5563 1411 5597
rect 1411 5563 1454 5597
rect 1382 5531 1454 5563
rect 1382 5395 1454 5467
rect 713 5240 719 5246
rect 719 5240 747 5246
rect 713 5212 747 5240
rect 813 5212 847 5246
rect 913 5212 947 5246
rect 1013 5240 1045 5246
rect 1045 5240 1047 5246
rect 1113 5240 1135 5246
rect 1135 5240 1147 5246
rect 1213 5240 1225 5246
rect 1225 5240 1247 5246
rect 1013 5212 1047 5240
rect 1113 5212 1147 5240
rect 1213 5212 1247 5240
rect 713 5112 747 5146
rect 813 5112 847 5146
rect 913 5112 947 5146
rect 1013 5112 1047 5146
rect 1113 5112 1147 5146
rect 1213 5112 1247 5146
rect 713 5012 747 5046
rect 813 5012 847 5046
rect 913 5012 947 5046
rect 1013 5012 1047 5046
rect 1113 5012 1147 5046
rect 1213 5012 1247 5046
rect 713 4914 747 4946
rect 713 4912 719 4914
rect 719 4912 747 4914
rect 813 4912 847 4946
rect 913 4912 947 4946
rect 1013 4914 1047 4946
rect 1113 4914 1147 4946
rect 1213 4914 1247 4946
rect 1013 4912 1045 4914
rect 1045 4912 1047 4914
rect 1113 4912 1135 4914
rect 1135 4912 1147 4914
rect 1213 4912 1225 4914
rect 1225 4912 1247 4914
rect 713 4824 747 4846
rect 713 4812 719 4824
rect 719 4812 747 4824
rect 813 4812 847 4846
rect 913 4812 947 4846
rect 1013 4824 1047 4846
rect 1113 4824 1147 4846
rect 1213 4824 1247 4846
rect 1013 4812 1045 4824
rect 1045 4812 1047 4824
rect 1113 4812 1135 4824
rect 1135 4812 1147 4824
rect 1213 4812 1225 4824
rect 1225 4812 1247 4824
rect 713 4734 747 4746
rect 713 4712 719 4734
rect 719 4712 747 4734
rect 813 4712 847 4746
rect 913 4712 947 4746
rect 1013 4734 1047 4746
rect 1113 4734 1147 4746
rect 1213 4734 1247 4746
rect 1013 4712 1045 4734
rect 1045 4712 1047 4734
rect 1113 4712 1135 4734
rect 1135 4712 1147 4734
rect 1213 4712 1225 4734
rect 1225 4712 1247 4734
rect 1382 4505 1454 4577
rect 1382 4410 1454 4441
rect 1382 4376 1411 4410
rect 1411 4376 1454 4410
rect 1382 4342 1454 4376
rect 2770 5597 2842 5630
rect 2770 5563 2799 5597
rect 2799 5563 2842 5597
rect 2770 5531 2842 5563
rect 2770 5395 2842 5467
rect 2101 5240 2107 5246
rect 2107 5240 2135 5246
rect 2101 5212 2135 5240
rect 2201 5212 2235 5246
rect 2301 5212 2335 5246
rect 2401 5240 2433 5246
rect 2433 5240 2435 5246
rect 2501 5240 2523 5246
rect 2523 5240 2535 5246
rect 2601 5240 2613 5246
rect 2613 5240 2635 5246
rect 2401 5212 2435 5240
rect 2501 5212 2535 5240
rect 2601 5212 2635 5240
rect 2101 5112 2135 5146
rect 2201 5112 2235 5146
rect 2301 5112 2335 5146
rect 2401 5112 2435 5146
rect 2501 5112 2535 5146
rect 2601 5112 2635 5146
rect 2101 5012 2135 5046
rect 2201 5012 2235 5046
rect 2301 5012 2335 5046
rect 2401 5012 2435 5046
rect 2501 5012 2535 5046
rect 2601 5012 2635 5046
rect 2101 4914 2135 4946
rect 2101 4912 2107 4914
rect 2107 4912 2135 4914
rect 2201 4912 2235 4946
rect 2301 4912 2335 4946
rect 2401 4914 2435 4946
rect 2501 4914 2535 4946
rect 2601 4914 2635 4946
rect 2401 4912 2433 4914
rect 2433 4912 2435 4914
rect 2501 4912 2523 4914
rect 2523 4912 2535 4914
rect 2601 4912 2613 4914
rect 2613 4912 2635 4914
rect 2101 4824 2135 4846
rect 2101 4812 2107 4824
rect 2107 4812 2135 4824
rect 2201 4812 2235 4846
rect 2301 4812 2335 4846
rect 2401 4824 2435 4846
rect 2501 4824 2535 4846
rect 2601 4824 2635 4846
rect 2401 4812 2433 4824
rect 2433 4812 2435 4824
rect 2501 4812 2523 4824
rect 2523 4812 2535 4824
rect 2601 4812 2613 4824
rect 2613 4812 2635 4824
rect 2101 4734 2135 4746
rect 2101 4712 2107 4734
rect 2107 4712 2135 4734
rect 2201 4712 2235 4746
rect 2301 4712 2335 4746
rect 2401 4734 2435 4746
rect 2501 4734 2535 4746
rect 2601 4734 2635 4746
rect 2401 4712 2433 4734
rect 2433 4712 2435 4734
rect 2501 4712 2523 4734
rect 2523 4712 2535 4734
rect 2601 4712 2613 4734
rect 2613 4712 2635 4734
rect 2770 4505 2842 4577
rect 2770 4410 2842 4441
rect 2770 4376 2799 4410
rect 2799 4376 2842 4410
rect 2770 4342 2842 4376
rect 3268 5597 3340 5630
rect 4158 5597 4230 5630
rect 3268 5563 3287 5597
rect 3287 5563 3340 5597
rect 4158 5563 4187 5597
rect 4187 5563 4230 5597
rect 3268 5531 3340 5563
rect 4158 5531 4230 5563
rect 3105 5462 3140 5467
rect 3140 5462 3174 5467
rect 3174 5462 3204 5467
rect 3105 5406 3204 5462
rect 3105 5395 3140 5406
rect 3140 5395 3174 5406
rect 3174 5395 3204 5406
rect 3105 4562 3140 4577
rect 3140 4562 3174 4577
rect 3174 4562 3204 4577
rect 3105 4506 3204 4562
rect 3105 4505 3140 4506
rect 3140 4505 3174 4506
rect 3174 4505 3204 4506
rect 3268 5395 3340 5467
rect 4158 5395 4230 5467
rect 3489 5240 3495 5246
rect 3495 5240 3523 5246
rect 3489 5212 3523 5240
rect 3589 5212 3623 5246
rect 3689 5212 3723 5246
rect 3789 5240 3821 5246
rect 3821 5240 3823 5246
rect 3889 5240 3911 5246
rect 3911 5240 3923 5246
rect 3989 5240 4001 5246
rect 4001 5240 4023 5246
rect 3789 5212 3823 5240
rect 3889 5212 3923 5240
rect 3989 5212 4023 5240
rect 3489 5112 3523 5146
rect 3589 5112 3623 5146
rect 3689 5112 3723 5146
rect 3789 5112 3823 5146
rect 3889 5112 3923 5146
rect 3989 5112 4023 5146
rect 3489 5012 3523 5046
rect 3589 5012 3623 5046
rect 3689 5012 3723 5046
rect 3789 5012 3823 5046
rect 3889 5012 3923 5046
rect 3989 5012 4023 5046
rect 3489 4914 3523 4946
rect 3489 4912 3495 4914
rect 3495 4912 3523 4914
rect 3589 4912 3623 4946
rect 3689 4912 3723 4946
rect 3789 4914 3823 4946
rect 3889 4914 3923 4946
rect 3989 4914 4023 4946
rect 3789 4912 3821 4914
rect 3821 4912 3823 4914
rect 3889 4912 3911 4914
rect 3911 4912 3923 4914
rect 3989 4912 4001 4914
rect 4001 4912 4023 4914
rect 3489 4824 3523 4846
rect 3489 4812 3495 4824
rect 3495 4812 3523 4824
rect 3589 4812 3623 4846
rect 3689 4812 3723 4846
rect 3789 4824 3823 4846
rect 3889 4824 3923 4846
rect 3989 4824 4023 4846
rect 3789 4812 3821 4824
rect 3821 4812 3823 4824
rect 3889 4812 3911 4824
rect 3911 4812 3923 4824
rect 3989 4812 4001 4824
rect 4001 4812 4023 4824
rect 3489 4734 3523 4746
rect 3489 4712 3495 4734
rect 3495 4712 3523 4734
rect 3589 4712 3623 4746
rect 3689 4712 3723 4746
rect 3789 4734 3823 4746
rect 3889 4734 3923 4746
rect 3989 4734 4023 4746
rect 3789 4712 3821 4734
rect 3821 4712 3823 4734
rect 3889 4712 3911 4734
rect 3911 4712 3923 4734
rect 3989 4712 4001 4734
rect 4001 4712 4023 4734
rect 3268 4505 3340 4577
rect 4158 4505 4230 4577
rect 4294 5462 4327 5467
rect 4327 5462 4361 5467
rect 4361 5462 4393 5467
rect 4294 5406 4393 5462
rect 4294 5395 4327 5406
rect 4327 5395 4361 5406
rect 4361 5395 4393 5406
rect 4294 4562 4327 4577
rect 4327 4562 4361 4577
rect 4361 4562 4393 4577
rect 4294 4506 4393 4562
rect 4294 4505 4327 4506
rect 4327 4505 4361 4506
rect 4361 4505 4393 4506
rect 3268 4410 3340 4441
rect 4158 4410 4230 4441
rect 3268 4376 3287 4410
rect 3287 4376 3340 4410
rect 4158 4376 4187 4410
rect 4187 4376 4230 4410
rect 3268 4342 3340 4376
rect 4158 4342 4230 4376
rect 4656 5597 4728 5630
rect 4656 5563 4675 5597
rect 4675 5563 4728 5597
rect 4656 5531 4728 5563
rect 4656 5395 4728 5467
rect 4877 5240 4883 5246
rect 4883 5240 4911 5246
rect 4877 5212 4911 5240
rect 4977 5212 5011 5246
rect 5077 5212 5111 5246
rect 5177 5240 5209 5246
rect 5209 5240 5211 5246
rect 5277 5240 5299 5246
rect 5299 5240 5311 5246
rect 5377 5240 5389 5246
rect 5389 5240 5411 5246
rect 5177 5212 5211 5240
rect 5277 5212 5311 5240
rect 5377 5212 5411 5240
rect 4877 5112 4911 5146
rect 4977 5112 5011 5146
rect 5077 5112 5111 5146
rect 5177 5112 5211 5146
rect 5277 5112 5311 5146
rect 5377 5112 5411 5146
rect 4877 5012 4911 5046
rect 4977 5012 5011 5046
rect 5077 5012 5111 5046
rect 5177 5012 5211 5046
rect 5277 5012 5311 5046
rect 5377 5012 5411 5046
rect 4877 4914 4911 4946
rect 4877 4912 4883 4914
rect 4883 4912 4911 4914
rect 4977 4912 5011 4946
rect 5077 4912 5111 4946
rect 5177 4914 5211 4946
rect 5277 4914 5311 4946
rect 5377 4914 5411 4946
rect 5177 4912 5209 4914
rect 5209 4912 5211 4914
rect 5277 4912 5299 4914
rect 5299 4912 5311 4914
rect 5377 4912 5389 4914
rect 5389 4912 5411 4914
rect 4877 4824 4911 4846
rect 4877 4812 4883 4824
rect 4883 4812 4911 4824
rect 4977 4812 5011 4846
rect 5077 4812 5111 4846
rect 5177 4824 5211 4846
rect 5277 4824 5311 4846
rect 5377 4824 5411 4846
rect 5177 4812 5209 4824
rect 5209 4812 5211 4824
rect 5277 4812 5299 4824
rect 5299 4812 5311 4824
rect 5377 4812 5389 4824
rect 5389 4812 5411 4824
rect 4877 4734 4911 4746
rect 4877 4712 4883 4734
rect 4883 4712 4911 4734
rect 4977 4712 5011 4746
rect 5077 4712 5111 4746
rect 5177 4734 5211 4746
rect 5277 4734 5311 4746
rect 5377 4734 5411 4746
rect 5177 4712 5209 4734
rect 5209 4712 5211 4734
rect 5277 4712 5299 4734
rect 5299 4712 5311 4734
rect 5377 4712 5389 4734
rect 5389 4712 5411 4734
rect 4656 4505 4728 4577
rect 4656 4410 4728 4441
rect 4656 4376 4675 4410
rect 4675 4376 4728 4410
rect 4656 4342 4728 4376
rect 6044 5597 6116 5630
rect 6044 5563 6063 5597
rect 6063 5563 6116 5597
rect 6044 5531 6116 5563
rect 6044 5395 6116 5467
rect 6265 5240 6271 5246
rect 6271 5240 6299 5246
rect 6265 5212 6299 5240
rect 6365 5212 6399 5246
rect 6465 5212 6499 5246
rect 6565 5240 6597 5246
rect 6597 5240 6599 5246
rect 6665 5240 6687 5246
rect 6687 5240 6699 5246
rect 6765 5240 6777 5246
rect 6777 5240 6799 5246
rect 6565 5212 6599 5240
rect 6665 5212 6699 5240
rect 6765 5212 6799 5240
rect 6265 5112 6299 5146
rect 6365 5112 6399 5146
rect 6465 5112 6499 5146
rect 6565 5112 6599 5146
rect 6665 5112 6699 5146
rect 6765 5112 6799 5146
rect 6265 5012 6299 5046
rect 6365 5012 6399 5046
rect 6465 5012 6499 5046
rect 6565 5012 6599 5046
rect 6665 5012 6699 5046
rect 6765 5012 6799 5046
rect 6265 4914 6299 4946
rect 6265 4912 6271 4914
rect 6271 4912 6299 4914
rect 6365 4912 6399 4946
rect 6465 4912 6499 4946
rect 6565 4914 6599 4946
rect 6665 4914 6699 4946
rect 6765 4914 6799 4946
rect 6565 4912 6597 4914
rect 6597 4912 6599 4914
rect 6665 4912 6687 4914
rect 6687 4912 6699 4914
rect 6765 4912 6777 4914
rect 6777 4912 6799 4914
rect 6265 4824 6299 4846
rect 6265 4812 6271 4824
rect 6271 4812 6299 4824
rect 6365 4812 6399 4846
rect 6465 4812 6499 4846
rect 6565 4824 6599 4846
rect 6665 4824 6699 4846
rect 6765 4824 6799 4846
rect 6565 4812 6597 4824
rect 6597 4812 6599 4824
rect 6665 4812 6687 4824
rect 6687 4812 6699 4824
rect 6765 4812 6777 4824
rect 6777 4812 6799 4824
rect 6265 4734 6299 4746
rect 6265 4712 6271 4734
rect 6271 4712 6299 4734
rect 6365 4712 6399 4746
rect 6465 4712 6499 4746
rect 6565 4734 6599 4746
rect 6665 4734 6699 4746
rect 6765 4734 6799 4746
rect 6565 4712 6597 4734
rect 6597 4712 6599 4734
rect 6665 4712 6687 4734
rect 6687 4712 6699 4734
rect 6765 4712 6777 4734
rect 6777 4712 6799 4734
rect 6044 4505 6116 4577
rect 6044 4410 6116 4441
rect 6044 4376 6063 4410
rect 6063 4376 6116 4410
rect 6044 4342 6116 4376
rect 1382 4209 1454 4242
rect 1382 4175 1411 4209
rect 1411 4175 1454 4209
rect 1382 4143 1454 4175
rect 1382 4007 1454 4079
rect 713 3852 719 3858
rect 719 3852 747 3858
rect 713 3824 747 3852
rect 813 3824 847 3858
rect 913 3824 947 3858
rect 1013 3852 1045 3858
rect 1045 3852 1047 3858
rect 1113 3852 1135 3858
rect 1135 3852 1147 3858
rect 1213 3852 1225 3858
rect 1225 3852 1247 3858
rect 1013 3824 1047 3852
rect 1113 3824 1147 3852
rect 1213 3824 1247 3852
rect 713 3724 747 3758
rect 813 3724 847 3758
rect 913 3724 947 3758
rect 1013 3724 1047 3758
rect 1113 3724 1147 3758
rect 1213 3724 1247 3758
rect 713 3624 747 3658
rect 813 3624 847 3658
rect 913 3624 947 3658
rect 1013 3624 1047 3658
rect 1113 3624 1147 3658
rect 1213 3624 1247 3658
rect 713 3526 747 3558
rect 713 3524 719 3526
rect 719 3524 747 3526
rect 813 3524 847 3558
rect 913 3524 947 3558
rect 1013 3526 1047 3558
rect 1113 3526 1147 3558
rect 1213 3526 1247 3558
rect 1013 3524 1045 3526
rect 1045 3524 1047 3526
rect 1113 3524 1135 3526
rect 1135 3524 1147 3526
rect 1213 3524 1225 3526
rect 1225 3524 1247 3526
rect 713 3436 747 3458
rect 713 3424 719 3436
rect 719 3424 747 3436
rect 813 3424 847 3458
rect 913 3424 947 3458
rect 1013 3436 1047 3458
rect 1113 3436 1147 3458
rect 1213 3436 1247 3458
rect 1013 3424 1045 3436
rect 1045 3424 1047 3436
rect 1113 3424 1135 3436
rect 1135 3424 1147 3436
rect 1213 3424 1225 3436
rect 1225 3424 1247 3436
rect 713 3346 747 3358
rect 713 3324 719 3346
rect 719 3324 747 3346
rect 813 3324 847 3358
rect 913 3324 947 3358
rect 1013 3346 1047 3358
rect 1113 3346 1147 3358
rect 1213 3346 1247 3358
rect 1013 3324 1045 3346
rect 1045 3324 1047 3346
rect 1113 3324 1135 3346
rect 1135 3324 1147 3346
rect 1213 3324 1225 3346
rect 1225 3324 1247 3346
rect 1382 3117 1454 3189
rect 1382 3022 1454 3053
rect 1382 2988 1411 3022
rect 1411 2988 1454 3022
rect 1382 2954 1454 2988
rect 2770 4209 2842 4242
rect 2770 4175 2799 4209
rect 2799 4175 2842 4209
rect 2770 4143 2842 4175
rect 2770 4007 2842 4079
rect 2101 3852 2107 3858
rect 2107 3852 2135 3858
rect 2101 3824 2135 3852
rect 2201 3824 2235 3858
rect 2301 3824 2335 3858
rect 2401 3852 2433 3858
rect 2433 3852 2435 3858
rect 2501 3852 2523 3858
rect 2523 3852 2535 3858
rect 2601 3852 2613 3858
rect 2613 3852 2635 3858
rect 2401 3824 2435 3852
rect 2501 3824 2535 3852
rect 2601 3824 2635 3852
rect 2101 3724 2135 3758
rect 2201 3724 2235 3758
rect 2301 3724 2335 3758
rect 2401 3724 2435 3758
rect 2501 3724 2535 3758
rect 2601 3724 2635 3758
rect 2101 3624 2135 3658
rect 2201 3624 2235 3658
rect 2301 3624 2335 3658
rect 2401 3624 2435 3658
rect 2501 3624 2535 3658
rect 2601 3624 2635 3658
rect 2101 3526 2135 3558
rect 2101 3524 2107 3526
rect 2107 3524 2135 3526
rect 2201 3524 2235 3558
rect 2301 3524 2335 3558
rect 2401 3526 2435 3558
rect 2501 3526 2535 3558
rect 2601 3526 2635 3558
rect 2401 3524 2433 3526
rect 2433 3524 2435 3526
rect 2501 3524 2523 3526
rect 2523 3524 2535 3526
rect 2601 3524 2613 3526
rect 2613 3524 2635 3526
rect 2101 3436 2135 3458
rect 2101 3424 2107 3436
rect 2107 3424 2135 3436
rect 2201 3424 2235 3458
rect 2301 3424 2335 3458
rect 2401 3436 2435 3458
rect 2501 3436 2535 3458
rect 2601 3436 2635 3458
rect 2401 3424 2433 3436
rect 2433 3424 2435 3436
rect 2501 3424 2523 3436
rect 2523 3424 2535 3436
rect 2601 3424 2613 3436
rect 2613 3424 2635 3436
rect 2101 3346 2135 3358
rect 2101 3324 2107 3346
rect 2107 3324 2135 3346
rect 2201 3324 2235 3358
rect 2301 3324 2335 3358
rect 2401 3346 2435 3358
rect 2501 3346 2535 3358
rect 2601 3346 2635 3358
rect 2401 3324 2433 3346
rect 2433 3324 2435 3346
rect 2501 3324 2523 3346
rect 2523 3324 2535 3346
rect 2601 3324 2613 3346
rect 2613 3324 2635 3346
rect 2906 4074 2939 4079
rect 2939 4074 2973 4079
rect 2973 4074 3005 4079
rect 2906 4018 3005 4074
rect 2906 4007 2939 4018
rect 2939 4007 2973 4018
rect 2973 4007 3005 4018
rect 3105 4074 3140 4079
rect 3140 4074 3174 4079
rect 3174 4074 3204 4079
rect 3105 4018 3204 4074
rect 3105 4007 3140 4018
rect 3140 4007 3174 4018
rect 3174 4007 3204 4018
rect 3268 4007 3340 4079
rect 4158 4007 4230 4079
rect 3489 3852 3495 3858
rect 3495 3852 3523 3858
rect 3489 3824 3523 3852
rect 3589 3824 3623 3858
rect 3689 3824 3723 3858
rect 3789 3852 3821 3858
rect 3821 3852 3823 3858
rect 3889 3852 3911 3858
rect 3911 3852 3923 3858
rect 3989 3852 4001 3858
rect 4001 3852 4023 3858
rect 3789 3824 3823 3852
rect 3889 3824 3923 3852
rect 3989 3824 4023 3852
rect 3489 3724 3523 3758
rect 3589 3724 3623 3758
rect 3689 3724 3723 3758
rect 3789 3724 3823 3758
rect 3889 3724 3923 3758
rect 3989 3724 4023 3758
rect 3489 3624 3523 3658
rect 3589 3624 3623 3658
rect 3689 3624 3723 3658
rect 3789 3624 3823 3658
rect 3889 3624 3923 3658
rect 3989 3624 4023 3658
rect 3489 3526 3523 3558
rect 3489 3524 3495 3526
rect 3495 3524 3523 3526
rect 3589 3524 3623 3558
rect 3689 3524 3723 3558
rect 3789 3526 3823 3558
rect 3889 3526 3923 3558
rect 3989 3526 4023 3558
rect 3789 3524 3821 3526
rect 3821 3524 3823 3526
rect 3889 3524 3911 3526
rect 3911 3524 3923 3526
rect 3989 3524 4001 3526
rect 4001 3524 4023 3526
rect 3489 3436 3523 3458
rect 3489 3424 3495 3436
rect 3495 3424 3523 3436
rect 3589 3424 3623 3458
rect 3689 3424 3723 3458
rect 3789 3436 3823 3458
rect 3889 3436 3923 3458
rect 3989 3436 4023 3458
rect 3789 3424 3821 3436
rect 3821 3424 3823 3436
rect 3889 3424 3911 3436
rect 3911 3424 3923 3436
rect 3989 3424 4001 3436
rect 4001 3424 4023 3436
rect 3489 3346 3523 3358
rect 3489 3324 3495 3346
rect 3495 3324 3523 3346
rect 3589 3324 3623 3358
rect 3689 3324 3723 3358
rect 3789 3346 3823 3358
rect 3889 3346 3923 3358
rect 3989 3346 4023 3358
rect 3789 3324 3821 3346
rect 3821 3324 3823 3346
rect 3889 3324 3911 3346
rect 3911 3324 3923 3346
rect 3989 3324 4001 3346
rect 4001 3324 4023 3346
rect 4294 4074 4327 4079
rect 4327 4074 4361 4079
rect 4361 4074 4393 4079
rect 4294 4018 4393 4074
rect 4294 4007 4327 4018
rect 4327 4007 4361 4018
rect 4361 4007 4393 4018
rect 4656 4209 4728 4242
rect 4656 4175 4675 4209
rect 4675 4175 4728 4209
rect 4656 4143 4728 4175
rect 4493 4074 4528 4079
rect 4528 4074 4562 4079
rect 4562 4074 4592 4079
rect 4493 4018 4592 4074
rect 4493 4007 4528 4018
rect 4528 4007 4562 4018
rect 4562 4007 4592 4018
rect 4656 4007 4728 4079
rect 4877 3852 4883 3858
rect 4883 3852 4911 3858
rect 4877 3824 4911 3852
rect 4977 3824 5011 3858
rect 5077 3824 5111 3858
rect 5177 3852 5209 3858
rect 5209 3852 5211 3858
rect 5277 3852 5299 3858
rect 5299 3852 5311 3858
rect 5377 3852 5389 3858
rect 5389 3852 5411 3858
rect 5177 3824 5211 3852
rect 5277 3824 5311 3852
rect 5377 3824 5411 3852
rect 4877 3724 4911 3758
rect 4977 3724 5011 3758
rect 5077 3724 5111 3758
rect 5177 3724 5211 3758
rect 5277 3724 5311 3758
rect 5377 3724 5411 3758
rect 4877 3624 4911 3658
rect 4977 3624 5011 3658
rect 5077 3624 5111 3658
rect 5177 3624 5211 3658
rect 5277 3624 5311 3658
rect 5377 3624 5411 3658
rect 4877 3526 4911 3558
rect 4877 3524 4883 3526
rect 4883 3524 4911 3526
rect 4977 3524 5011 3558
rect 5077 3524 5111 3558
rect 5177 3526 5211 3558
rect 5277 3526 5311 3558
rect 5377 3526 5411 3558
rect 5177 3524 5209 3526
rect 5209 3524 5211 3526
rect 5277 3524 5299 3526
rect 5299 3524 5311 3526
rect 5377 3524 5389 3526
rect 5389 3524 5411 3526
rect 4877 3436 4911 3458
rect 4877 3424 4883 3436
rect 4883 3424 4911 3436
rect 4977 3424 5011 3458
rect 5077 3424 5111 3458
rect 5177 3436 5211 3458
rect 5277 3436 5311 3458
rect 5377 3436 5411 3458
rect 5177 3424 5209 3436
rect 5209 3424 5211 3436
rect 5277 3424 5299 3436
rect 5299 3424 5311 3436
rect 5377 3424 5389 3436
rect 5389 3424 5411 3436
rect 4877 3346 4911 3358
rect 4877 3324 4883 3346
rect 4883 3324 4911 3346
rect 4977 3324 5011 3358
rect 5077 3324 5111 3358
rect 5177 3346 5211 3358
rect 5277 3346 5311 3358
rect 5377 3346 5411 3358
rect 5177 3324 5209 3346
rect 5209 3324 5211 3346
rect 5277 3324 5299 3346
rect 5299 3324 5311 3346
rect 5377 3324 5389 3346
rect 5389 3324 5411 3346
rect 6044 4209 6116 4242
rect 6044 4175 6063 4209
rect 6063 4175 6116 4209
rect 6044 4143 6116 4175
rect 6044 4007 6116 4079
rect 6265 3852 6271 3858
rect 6271 3852 6299 3858
rect 6265 3824 6299 3852
rect 6365 3824 6399 3858
rect 6465 3824 6499 3858
rect 6565 3852 6597 3858
rect 6597 3852 6599 3858
rect 6665 3852 6687 3858
rect 6687 3852 6699 3858
rect 6765 3852 6777 3858
rect 6777 3852 6799 3858
rect 6565 3824 6599 3852
rect 6665 3824 6699 3852
rect 6765 3824 6799 3852
rect 6265 3724 6299 3758
rect 6365 3724 6399 3758
rect 6465 3724 6499 3758
rect 6565 3724 6599 3758
rect 6665 3724 6699 3758
rect 6765 3724 6799 3758
rect 6265 3624 6299 3658
rect 6365 3624 6399 3658
rect 6465 3624 6499 3658
rect 6565 3624 6599 3658
rect 6665 3624 6699 3658
rect 6765 3624 6799 3658
rect 6265 3526 6299 3558
rect 6265 3524 6271 3526
rect 6271 3524 6299 3526
rect 6365 3524 6399 3558
rect 6465 3524 6499 3558
rect 6565 3526 6599 3558
rect 6665 3526 6699 3558
rect 6765 3526 6799 3558
rect 6565 3524 6597 3526
rect 6597 3524 6599 3526
rect 6665 3524 6687 3526
rect 6687 3524 6699 3526
rect 6765 3524 6777 3526
rect 6777 3524 6799 3526
rect 6265 3436 6299 3458
rect 6265 3424 6271 3436
rect 6271 3424 6299 3436
rect 6365 3424 6399 3458
rect 6465 3424 6499 3458
rect 6565 3436 6599 3458
rect 6665 3436 6699 3458
rect 6765 3436 6799 3458
rect 6565 3424 6597 3436
rect 6597 3424 6599 3436
rect 6665 3424 6687 3436
rect 6687 3424 6699 3436
rect 6765 3424 6777 3436
rect 6777 3424 6799 3436
rect 6265 3346 6299 3358
rect 6265 3324 6271 3346
rect 6271 3324 6299 3346
rect 6365 3324 6399 3358
rect 6465 3324 6499 3358
rect 6565 3346 6599 3358
rect 6665 3346 6699 3358
rect 6765 3346 6799 3358
rect 6565 3324 6597 3346
rect 6597 3324 6599 3346
rect 6665 3324 6687 3346
rect 6687 3324 6699 3346
rect 6765 3324 6777 3346
rect 6777 3324 6799 3346
rect 6044 3117 6116 3189
rect 6044 3022 6116 3053
rect 6044 2988 6063 3022
rect 6063 2988 6116 3022
rect 6044 2954 6116 2988
rect 1382 2821 1454 2854
rect 1382 2787 1411 2821
rect 1411 2787 1454 2821
rect 1382 2755 1454 2787
rect 1382 2619 1454 2691
rect 713 2464 719 2470
rect 719 2464 747 2470
rect 713 2436 747 2464
rect 813 2436 847 2470
rect 913 2436 947 2470
rect 1013 2464 1045 2470
rect 1045 2464 1047 2470
rect 1113 2464 1135 2470
rect 1135 2464 1147 2470
rect 1213 2464 1225 2470
rect 1225 2464 1247 2470
rect 1013 2436 1047 2464
rect 1113 2436 1147 2464
rect 1213 2436 1247 2464
rect 713 2336 747 2370
rect 813 2336 847 2370
rect 913 2336 947 2370
rect 1013 2336 1047 2370
rect 1113 2336 1147 2370
rect 1213 2336 1247 2370
rect 713 2236 747 2270
rect 813 2236 847 2270
rect 913 2236 947 2270
rect 1013 2236 1047 2270
rect 1113 2236 1147 2270
rect 1213 2236 1247 2270
rect 713 2138 747 2170
rect 713 2136 719 2138
rect 719 2136 747 2138
rect 813 2136 847 2170
rect 913 2136 947 2170
rect 1013 2138 1047 2170
rect 1113 2138 1147 2170
rect 1213 2138 1247 2170
rect 1013 2136 1045 2138
rect 1045 2136 1047 2138
rect 1113 2136 1135 2138
rect 1135 2136 1147 2138
rect 1213 2136 1225 2138
rect 1225 2136 1247 2138
rect 713 2048 747 2070
rect 713 2036 719 2048
rect 719 2036 747 2048
rect 813 2036 847 2070
rect 913 2036 947 2070
rect 1013 2048 1047 2070
rect 1113 2048 1147 2070
rect 1213 2048 1247 2070
rect 1013 2036 1045 2048
rect 1045 2036 1047 2048
rect 1113 2036 1135 2048
rect 1135 2036 1147 2048
rect 1213 2036 1225 2048
rect 1225 2036 1247 2048
rect 713 1958 747 1970
rect 713 1936 719 1958
rect 719 1936 747 1958
rect 813 1936 847 1970
rect 913 1936 947 1970
rect 1013 1958 1047 1970
rect 1113 1958 1147 1970
rect 1213 1958 1247 1970
rect 1013 1936 1045 1958
rect 1045 1936 1047 1958
rect 1113 1936 1135 1958
rect 1135 1936 1147 1958
rect 1213 1936 1225 1958
rect 1225 1936 1247 1958
rect 1518 2686 1551 2691
rect 1551 2686 1585 2691
rect 1585 2686 1617 2691
rect 1518 2630 1617 2686
rect 1518 2619 1551 2630
rect 1551 2619 1585 2630
rect 1585 2619 1617 2630
rect 1717 2686 1752 2691
rect 1752 2686 1786 2691
rect 1786 2686 1816 2691
rect 1717 2630 1816 2686
rect 1717 2619 1752 2630
rect 1752 2619 1786 2630
rect 1786 2619 1816 2630
rect 1880 2619 1952 2691
rect 2770 2619 2842 2691
rect 2101 2464 2107 2470
rect 2107 2464 2135 2470
rect 2101 2436 2135 2464
rect 2201 2436 2235 2470
rect 2301 2436 2335 2470
rect 2401 2464 2433 2470
rect 2433 2464 2435 2470
rect 2501 2464 2523 2470
rect 2523 2464 2535 2470
rect 2601 2464 2613 2470
rect 2613 2464 2635 2470
rect 2401 2436 2435 2464
rect 2501 2436 2535 2464
rect 2601 2436 2635 2464
rect 2101 2336 2135 2370
rect 2201 2336 2235 2370
rect 2301 2336 2335 2370
rect 2401 2336 2435 2370
rect 2501 2336 2535 2370
rect 2601 2336 2635 2370
rect 2101 2236 2135 2270
rect 2201 2236 2235 2270
rect 2301 2236 2335 2270
rect 2401 2236 2435 2270
rect 2501 2236 2535 2270
rect 2601 2236 2635 2270
rect 2101 2138 2135 2170
rect 2101 2136 2107 2138
rect 2107 2136 2135 2138
rect 2201 2136 2235 2170
rect 2301 2136 2335 2170
rect 2401 2138 2435 2170
rect 2501 2138 2535 2170
rect 2601 2138 2635 2170
rect 2401 2136 2433 2138
rect 2433 2136 2435 2138
rect 2501 2136 2523 2138
rect 2523 2136 2535 2138
rect 2601 2136 2613 2138
rect 2613 2136 2635 2138
rect 2101 2048 2135 2070
rect 2101 2036 2107 2048
rect 2107 2036 2135 2048
rect 2201 2036 2235 2070
rect 2301 2036 2335 2070
rect 2401 2048 2435 2070
rect 2501 2048 2535 2070
rect 2601 2048 2635 2070
rect 2401 2036 2433 2048
rect 2433 2036 2435 2048
rect 2501 2036 2523 2048
rect 2523 2036 2535 2048
rect 2601 2036 2613 2048
rect 2613 2036 2635 2048
rect 2101 1958 2135 1970
rect 2101 1936 2107 1958
rect 2107 1936 2135 1958
rect 2201 1936 2235 1970
rect 2301 1936 2335 1970
rect 2401 1958 2435 1970
rect 2501 1958 2535 1970
rect 2601 1958 2635 1970
rect 2401 1936 2433 1958
rect 2433 1936 2435 1958
rect 2501 1936 2523 1958
rect 2523 1936 2535 1958
rect 2601 1936 2613 1958
rect 2613 1936 2635 1958
rect 2906 2686 2939 2691
rect 2939 2686 2973 2691
rect 2973 2686 3005 2691
rect 2906 2630 3005 2686
rect 2906 2619 2939 2630
rect 2939 2619 2973 2630
rect 2973 2619 3005 2630
rect 3105 2686 3140 2691
rect 3140 2686 3174 2691
rect 3174 2686 3204 2691
rect 3105 2630 3204 2686
rect 3105 2619 3140 2630
rect 3140 2619 3174 2630
rect 3174 2619 3204 2630
rect 3268 2619 3340 2691
rect 4158 2619 4230 2691
rect 3489 2464 3495 2470
rect 3495 2464 3523 2470
rect 3489 2436 3523 2464
rect 3589 2436 3623 2470
rect 3689 2436 3723 2470
rect 3789 2464 3821 2470
rect 3821 2464 3823 2470
rect 3889 2464 3911 2470
rect 3911 2464 3923 2470
rect 3989 2464 4001 2470
rect 4001 2464 4023 2470
rect 3789 2436 3823 2464
rect 3889 2436 3923 2464
rect 3989 2436 4023 2464
rect 3489 2336 3523 2370
rect 3589 2336 3623 2370
rect 3689 2336 3723 2370
rect 3789 2336 3823 2370
rect 3889 2336 3923 2370
rect 3989 2336 4023 2370
rect 3489 2236 3523 2270
rect 3589 2236 3623 2270
rect 3689 2236 3723 2270
rect 3789 2236 3823 2270
rect 3889 2236 3923 2270
rect 3989 2236 4023 2270
rect 3489 2138 3523 2170
rect 3489 2136 3495 2138
rect 3495 2136 3523 2138
rect 3589 2136 3623 2170
rect 3689 2136 3723 2170
rect 3789 2138 3823 2170
rect 3889 2138 3923 2170
rect 3989 2138 4023 2170
rect 3789 2136 3821 2138
rect 3821 2136 3823 2138
rect 3889 2136 3911 2138
rect 3911 2136 3923 2138
rect 3989 2136 4001 2138
rect 4001 2136 4023 2138
rect 3489 2048 3523 2070
rect 3489 2036 3495 2048
rect 3495 2036 3523 2048
rect 3589 2036 3623 2070
rect 3689 2036 3723 2070
rect 3789 2048 3823 2070
rect 3889 2048 3923 2070
rect 3989 2048 4023 2070
rect 3789 2036 3821 2048
rect 3821 2036 3823 2048
rect 3889 2036 3911 2048
rect 3911 2036 3923 2048
rect 3989 2036 4001 2048
rect 4001 2036 4023 2048
rect 3489 1958 3523 1970
rect 3489 1936 3495 1958
rect 3495 1936 3523 1958
rect 3589 1936 3623 1970
rect 3689 1936 3723 1970
rect 3789 1958 3823 1970
rect 3889 1958 3923 1970
rect 3989 1958 4023 1970
rect 3789 1936 3821 1958
rect 3821 1936 3823 1958
rect 3889 1936 3911 1958
rect 3911 1936 3923 1958
rect 3989 1936 4001 1958
rect 4001 1936 4023 1958
rect 4294 2686 4327 2691
rect 4327 2686 4361 2691
rect 4361 2686 4393 2691
rect 4294 2630 4393 2686
rect 4294 2619 4327 2630
rect 4327 2619 4361 2630
rect 4361 2619 4393 2630
rect 6043 2821 6115 2854
rect 6043 2787 6063 2821
rect 6063 2787 6115 2821
rect 6043 2755 6115 2787
rect 4493 2686 4528 2691
rect 4528 2686 4562 2691
rect 4562 2686 4592 2691
rect 4493 2630 4592 2686
rect 4493 2619 4528 2630
rect 4528 2619 4562 2630
rect 4562 2619 4592 2630
rect 4656 2619 4728 2691
rect 5546 2619 5618 2691
rect 4877 2464 4883 2470
rect 4883 2464 4911 2470
rect 4877 2436 4911 2464
rect 4977 2436 5011 2470
rect 5077 2436 5111 2470
rect 5177 2464 5209 2470
rect 5209 2464 5211 2470
rect 5277 2464 5299 2470
rect 5299 2464 5311 2470
rect 5377 2464 5389 2470
rect 5389 2464 5411 2470
rect 5177 2436 5211 2464
rect 5277 2436 5311 2464
rect 5377 2436 5411 2464
rect 4877 2336 4911 2370
rect 4977 2336 5011 2370
rect 5077 2336 5111 2370
rect 5177 2336 5211 2370
rect 5277 2336 5311 2370
rect 5377 2336 5411 2370
rect 4877 2236 4911 2270
rect 4977 2236 5011 2270
rect 5077 2236 5111 2270
rect 5177 2236 5211 2270
rect 5277 2236 5311 2270
rect 5377 2236 5411 2270
rect 4877 2138 4911 2170
rect 4877 2136 4883 2138
rect 4883 2136 4911 2138
rect 4977 2136 5011 2170
rect 5077 2136 5111 2170
rect 5177 2138 5211 2170
rect 5277 2138 5311 2170
rect 5377 2138 5411 2170
rect 5177 2136 5209 2138
rect 5209 2136 5211 2138
rect 5277 2136 5299 2138
rect 5299 2136 5311 2138
rect 5377 2136 5389 2138
rect 5389 2136 5411 2138
rect 4877 2048 4911 2070
rect 4877 2036 4883 2048
rect 4883 2036 4911 2048
rect 4977 2036 5011 2070
rect 5077 2036 5111 2070
rect 5177 2048 5211 2070
rect 5277 2048 5311 2070
rect 5377 2048 5411 2070
rect 5177 2036 5209 2048
rect 5209 2036 5211 2048
rect 5277 2036 5299 2048
rect 5299 2036 5311 2048
rect 5377 2036 5389 2048
rect 5389 2036 5411 2048
rect 4877 1958 4911 1970
rect 4877 1936 4883 1958
rect 4883 1936 4911 1958
rect 4977 1936 5011 1970
rect 5077 1936 5111 1970
rect 5177 1958 5211 1970
rect 5277 1958 5311 1970
rect 5377 1958 5411 1970
rect 5177 1936 5209 1958
rect 5209 1936 5211 1958
rect 5277 1936 5299 1958
rect 5299 1936 5311 1958
rect 5377 1936 5389 1958
rect 5389 1936 5411 1958
rect 5682 2686 5715 2691
rect 5715 2686 5749 2691
rect 5749 2686 5781 2691
rect 5682 2630 5781 2686
rect 5682 2619 5715 2630
rect 5715 2619 5749 2630
rect 5749 2619 5781 2630
rect 5880 2686 5916 2691
rect 5916 2686 5950 2691
rect 5950 2686 5979 2691
rect 5880 2630 5979 2686
rect 5880 2619 5916 2630
rect 5916 2619 5950 2630
rect 5950 2619 5979 2630
rect 6043 2619 6115 2691
rect 6265 2464 6271 2470
rect 6271 2464 6299 2470
rect 6265 2436 6299 2464
rect 6365 2436 6399 2470
rect 6465 2436 6499 2470
rect 6565 2464 6597 2470
rect 6597 2464 6599 2470
rect 6665 2464 6687 2470
rect 6687 2464 6699 2470
rect 6765 2464 6777 2470
rect 6777 2464 6799 2470
rect 6565 2436 6599 2464
rect 6665 2436 6699 2464
rect 6765 2436 6799 2464
rect 6265 2336 6299 2370
rect 6365 2336 6399 2370
rect 6465 2336 6499 2370
rect 6565 2336 6599 2370
rect 6665 2336 6699 2370
rect 6765 2336 6799 2370
rect 6265 2236 6299 2270
rect 6365 2236 6399 2270
rect 6465 2236 6499 2270
rect 6565 2236 6599 2270
rect 6665 2236 6699 2270
rect 6765 2236 6799 2270
rect 6265 2138 6299 2170
rect 6265 2136 6271 2138
rect 6271 2136 6299 2138
rect 6365 2136 6399 2170
rect 6465 2136 6499 2170
rect 6565 2138 6599 2170
rect 6665 2138 6699 2170
rect 6765 2138 6799 2170
rect 6565 2136 6597 2138
rect 6597 2136 6599 2138
rect 6665 2136 6687 2138
rect 6687 2136 6699 2138
rect 6765 2136 6777 2138
rect 6777 2136 6799 2138
rect 6265 2048 6299 2070
rect 6265 2036 6271 2048
rect 6271 2036 6299 2048
rect 6365 2036 6399 2070
rect 6465 2036 6499 2070
rect 6565 2048 6599 2070
rect 6665 2048 6699 2070
rect 6765 2048 6799 2070
rect 6565 2036 6597 2048
rect 6597 2036 6599 2048
rect 6665 2036 6687 2048
rect 6687 2036 6699 2048
rect 6765 2036 6777 2048
rect 6777 2036 6799 2048
rect 6265 1958 6299 1970
rect 6265 1936 6271 1958
rect 6271 1936 6299 1958
rect 6365 1936 6399 1970
rect 6465 1936 6499 1970
rect 6565 1958 6599 1970
rect 6665 1958 6699 1970
rect 6765 1958 6799 1970
rect 6565 1936 6597 1958
rect 6597 1936 6599 1958
rect 6665 1936 6687 1958
rect 6687 1936 6699 1958
rect 6765 1936 6777 1958
rect 6777 1936 6799 1958
<< metal1 >>
rect -17506 22697 -17460 22701
rect 8662 22697 8708 22701
rect -17512 22691 8714 22697
rect -17512 22651 -17500 22691
rect -17506 20892 -17500 22651
rect -17512 20852 -17500 20892
rect -17466 22651 8668 22657
rect -17466 22551 -17460 22651
rect 8662 22551 8668 22651
rect -17466 22545 -16928 22551
rect -17466 22507 -17337 22545
rect -16940 22507 -16928 22545
rect -17466 22501 -16928 22507
rect -13550 22545 -12592 22551
rect -13550 22507 -13538 22545
rect -13141 22507 -13001 22545
rect -12604 22507 -12592 22545
rect -13550 22501 -12592 22507
rect -9214 22545 -8256 22551
rect -9214 22507 -9202 22545
rect -8805 22507 -8665 22545
rect -8268 22507 -8256 22545
rect -9214 22501 -8256 22507
rect -4878 22545 -3920 22551
rect -4878 22507 -4866 22545
rect -4469 22507 -4329 22545
rect -3932 22507 -3920 22545
rect -4878 22501 -3920 22507
rect -542 22545 416 22551
rect -542 22507 -530 22545
rect -133 22507 7 22545
rect 404 22507 416 22545
rect -542 22501 416 22507
rect 3794 22545 4752 22551
rect 3794 22507 3806 22545
rect 4203 22507 4343 22545
rect 4740 22507 4752 22545
rect 3794 22501 4752 22507
rect 8130 22545 8668 22551
rect 8130 22507 8142 22545
rect 8539 22507 8668 22545
rect 8130 22501 8668 22507
rect -17466 21057 -17460 22501
rect -17365 22325 -17355 22395
rect -16923 22325 -16913 22395
rect -13001 22386 -12949 22396
rect -13550 22379 -13046 22385
rect -13550 22341 -13538 22379
rect -13141 22341 -13046 22379
rect -13550 22335 -13046 22341
rect -13013 22335 -13001 22385
rect -8857 22386 -8805 22396
rect -12949 22379 -12592 22385
rect -12604 22341 -12592 22379
rect -17365 22159 -17355 22229
rect -16923 22159 -16913 22229
rect -13193 22220 -13141 22230
rect -13550 22213 -13193 22219
rect -13096 22219 -13046 22335
rect -12949 22335 -12592 22341
rect -9214 22379 -8857 22385
rect -4329 22386 -4277 22396
rect -9214 22341 -9202 22379
rect -9214 22335 -8857 22341
rect -13001 22324 -12949 22334
rect -8805 22335 -8793 22385
rect -8760 22379 -8256 22385
rect -8760 22341 -8665 22379
rect -8268 22341 -8256 22379
rect -8760 22335 -8256 22341
rect -4878 22379 -4374 22385
rect -4878 22341 -4866 22379
rect -4469 22341 -4374 22379
rect -4878 22335 -4374 22341
rect -4341 22335 -4329 22385
rect -185 22386 -133 22396
rect -4277 22379 -3920 22385
rect -3932 22341 -3920 22379
rect -8857 22324 -8805 22334
rect -8760 22219 -8710 22335
rect -8665 22220 -8613 22230
rect -13550 22175 -13538 22213
rect -13550 22169 -13193 22175
rect -13141 22169 -13129 22219
rect -13096 22213 -12592 22219
rect -13096 22175 -13001 22213
rect -12604 22175 -12592 22213
rect -13096 22169 -12592 22175
rect -9214 22213 -8710 22219
rect -9214 22175 -9202 22213
rect -8805 22175 -8710 22213
rect -9214 22169 -8710 22175
rect -8677 22169 -8665 22219
rect -4521 22220 -4469 22230
rect -8613 22213 -8256 22219
rect -8268 22175 -8256 22213
rect -13193 22158 -13141 22168
rect -8613 22169 -8256 22175
rect -4878 22213 -4521 22219
rect -4424 22219 -4374 22335
rect -4277 22335 -3920 22341
rect -542 22379 -185 22385
rect 4343 22386 4395 22396
rect -542 22341 -530 22379
rect -542 22335 -185 22341
rect -4329 22324 -4277 22334
rect -133 22335 -121 22385
rect -88 22379 416 22385
rect -88 22341 7 22379
rect 404 22341 416 22379
rect -88 22335 416 22341
rect 3794 22379 4298 22385
rect 3794 22341 3806 22379
rect 4203 22341 4298 22379
rect 3794 22335 4298 22341
rect 4331 22335 4343 22385
rect 8487 22386 8539 22396
rect 4395 22379 4752 22385
rect 4740 22341 4752 22379
rect -185 22324 -133 22334
rect -88 22219 -38 22335
rect 7 22220 59 22230
rect -4878 22175 -4866 22213
rect -4878 22169 -4521 22175
rect -8665 22158 -8613 22168
rect -4469 22169 -4457 22219
rect -4424 22213 -3920 22219
rect -4424 22175 -4329 22213
rect -3932 22175 -3920 22213
rect -4424 22169 -3920 22175
rect -542 22213 -38 22219
rect -542 22175 -530 22213
rect -133 22175 -38 22213
rect -542 22169 -38 22175
rect -5 22169 7 22219
rect 4151 22220 4203 22230
rect 59 22213 416 22219
rect 404 22175 416 22213
rect -4521 22158 -4469 22168
rect 59 22169 416 22175
rect 3794 22213 4151 22219
rect 4248 22219 4298 22335
rect 4395 22335 4752 22341
rect 8130 22379 8487 22385
rect 8130 22341 8142 22379
rect 8130 22335 8487 22341
rect 4343 22324 4395 22334
rect 8539 22335 8551 22385
rect 8487 22324 8539 22334
rect 3794 22175 3806 22213
rect 3794 22169 4151 22175
rect 7 22158 59 22168
rect 4203 22169 4215 22219
rect 4248 22213 4752 22219
rect 4248 22175 4343 22213
rect 4740 22175 4752 22213
rect 4248 22169 4752 22175
rect 8130 22213 8634 22219
rect 8130 22175 8142 22213
rect 8539 22175 8634 22213
rect 8130 22169 8634 22175
rect 4151 22158 4203 22168
rect -13001 22054 -12949 22064
rect -17432 22047 -16928 22053
rect -17432 22009 -17337 22047
rect -16940 22009 -16928 22047
rect -17432 22003 -16928 22009
rect -13550 22047 -13046 22053
rect -13550 22009 -13538 22047
rect -13141 22009 -13046 22047
rect -13550 22003 -13046 22009
rect -13013 22003 -13001 22053
rect -8857 22054 -8805 22064
rect -12949 22047 -12592 22053
rect -12604 22009 -12592 22047
rect -17432 21555 -17382 22003
rect -13193 21888 -13141 21898
rect -17349 21881 -16928 21887
rect -17349 21843 -17337 21881
rect -16940 21843 -16928 21881
rect -17349 21837 -16928 21843
rect -13550 21881 -13193 21887
rect -13096 21887 -13046 22003
rect -12949 22003 -12592 22009
rect -9214 22047 -8857 22053
rect -4329 22054 -4277 22064
rect -9214 22009 -9202 22047
rect -9214 22003 -8857 22009
rect -13001 21992 -12949 22002
rect -8805 22003 -8793 22053
rect -8760 22047 -8256 22053
rect -8760 22009 -8665 22047
rect -8268 22009 -8256 22047
rect -8760 22003 -8256 22009
rect -4878 22047 -4374 22053
rect -4878 22009 -4866 22047
rect -4469 22009 -4374 22047
rect -4878 22003 -4374 22009
rect -4341 22003 -4329 22053
rect -185 22054 -133 22064
rect 4343 22054 4395 22064
rect -4277 22047 -3920 22053
rect -3932 22009 -3920 22047
rect -8857 21992 -8805 22002
rect -8760 21887 -8710 22003
rect -4424 21964 -4374 22003
rect -4277 22003 -3920 22009
rect -542 22047 -185 22053
rect 342 22053 352 22054
rect -542 22009 -530 22047
rect -542 22003 -185 22009
rect -4329 21992 -4277 22002
rect -133 22003 -121 22053
rect -88 22047 352 22053
rect 404 22053 414 22054
rect -88 22009 7 22047
rect -88 22003 352 22009
rect -185 21992 -133 22002
rect -88 21964 -38 22003
rect 342 22002 352 22003
rect 404 22003 416 22053
rect 3794 22047 4298 22053
rect 3794 22009 3806 22047
rect 4203 22009 4298 22047
rect 3794 22003 4298 22009
rect 4331 22003 4343 22053
rect 8487 22054 8539 22064
rect 4395 22047 4752 22053
rect 4740 22009 4752 22047
rect 404 22002 414 22003
rect -4424 21926 -38 21964
rect -8665 21888 -8613 21898
rect -13550 21843 -13538 21881
rect -13550 21837 -13193 21843
rect -17349 21721 -17299 21837
rect -13141 21837 -13129 21887
rect -13096 21881 -12592 21887
rect -13096 21843 -13001 21881
rect -12604 21843 -12592 21881
rect -13096 21837 -12592 21843
rect -9214 21881 -8710 21887
rect -9214 21843 -9202 21881
rect -8805 21843 -8710 21881
rect -9214 21837 -8710 21843
rect -8677 21837 -8665 21887
rect -4521 21888 -4469 21898
rect 7 21888 59 21898
rect -8613 21881 -8256 21887
rect -8268 21843 -8256 21881
rect -13193 21826 -13141 21836
rect -8613 21837 -8256 21843
rect -4878 21881 -4521 21887
rect -540 21887 -530 21888
rect -4878 21843 -4866 21881
rect -4878 21837 -4521 21843
rect -8665 21826 -8613 21836
rect -4469 21837 -4457 21887
rect -4341 21881 -3920 21887
rect -4341 21843 -4329 21881
rect -3932 21843 -3920 21881
rect -4341 21837 -3920 21843
rect -542 21837 -530 21887
rect -133 21887 -123 21888
rect -4521 21826 -4469 21836
rect -4341 21798 -4294 21837
rect -540 21836 -530 21837
rect -133 21837 -121 21887
rect -5 21837 7 21887
rect 4151 21888 4203 21898
rect 59 21881 416 21887
rect 404 21843 416 21881
rect -133 21836 -123 21837
rect 59 21837 416 21843
rect 3794 21881 4151 21887
rect 4248 21887 4298 22003
rect 4395 22003 4752 22009
rect 8130 22047 8487 22053
rect 8130 22009 8142 22047
rect 8130 22003 8487 22009
rect 4343 21992 4395 22002
rect 8539 22003 8551 22053
rect 8487 21992 8539 22002
rect 4678 21887 4688 21888
rect 3794 21843 3806 21881
rect 3794 21837 4151 21843
rect 7 21826 59 21836
rect 4203 21837 4215 21887
rect 4248 21881 4688 21887
rect 4740 21887 4750 21888
rect 8584 21887 8634 22169
rect 4248 21843 4343 21881
rect 4248 21837 4688 21843
rect 4678 21836 4688 21837
rect 4740 21837 4752 21887
rect 8130 21881 8634 21887
rect 8130 21843 8142 21881
rect 8539 21843 8634 21881
rect 8130 21837 8634 21843
rect 4740 21836 4750 21837
rect 4151 21826 4203 21836
rect -4504 21751 -4294 21798
rect -13193 21722 -13141 21732
rect -17349 21715 -16928 21721
rect -17349 21677 -17337 21715
rect -16940 21677 -16928 21715
rect -17349 21671 -16928 21677
rect -13550 21715 -13193 21721
rect -8665 21722 -8613 21732
rect -13550 21677 -13538 21715
rect -13550 21671 -13193 21677
rect -13141 21671 -13129 21721
rect -13096 21715 -12592 21721
rect -13096 21677 -13001 21715
rect -12604 21677 -12592 21715
rect -13096 21671 -12592 21677
rect -9214 21715 -8710 21721
rect -9214 21677 -9202 21715
rect -8805 21677 -8710 21715
rect -9214 21671 -8710 21677
rect -8677 21671 -8665 21721
rect -4504 21721 -4457 21751
rect 7 21722 59 21732
rect -8613 21715 -8256 21721
rect -8268 21677 -8256 21715
rect -13193 21660 -13141 21670
rect -13096 21555 -13046 21671
rect -13001 21556 -12949 21566
rect -17432 21549 -16928 21555
rect -17432 21511 -17337 21549
rect -16940 21511 -16928 21549
rect -17432 21505 -16928 21511
rect -13550 21549 -13046 21555
rect -13550 21511 -13538 21549
rect -13141 21511 -13046 21549
rect -13550 21505 -13046 21511
rect -13013 21505 -13001 21555
rect -8857 21556 -8805 21566
rect -12949 21549 -12592 21555
rect -12604 21511 -12592 21549
rect -12949 21505 -12592 21511
rect -9214 21549 -8857 21555
rect -8760 21555 -8710 21671
rect -8613 21671 -8256 21677
rect -4878 21715 -4457 21721
rect -4878 21677 -4866 21715
rect -4469 21677 -4457 21715
rect -4878 21671 -4457 21677
rect -4424 21715 -3920 21721
rect -4424 21677 -4329 21715
rect -3932 21677 -3920 21715
rect -4424 21671 -3920 21677
rect -542 21715 -38 21721
rect -542 21677 -530 21715
rect -133 21677 -38 21715
rect -542 21671 -38 21677
rect -5 21671 7 21721
rect 4151 21722 4203 21732
rect 59 21715 416 21721
rect 404 21677 416 21715
rect -8665 21660 -8613 21670
rect -4424 21643 -4374 21671
rect -88 21643 -38 21671
rect 59 21671 416 21677
rect 3794 21715 4151 21721
rect 3794 21677 3806 21715
rect 3794 21671 4151 21677
rect 7 21660 59 21670
rect 4203 21671 4215 21721
rect 4248 21715 4752 21721
rect 4248 21677 4343 21715
rect 4740 21677 4752 21715
rect 4248 21671 4752 21677
rect 8130 21715 8634 21721
rect 8130 21677 8142 21715
rect 8539 21677 8634 21715
rect 8130 21671 8634 21677
rect 4151 21660 4203 21670
rect -4424 21594 -38 21643
rect -4424 21555 -4374 21594
rect -4329 21556 -4277 21566
rect -9214 21511 -9202 21549
rect -9214 21505 -8857 21511
rect -13001 21494 -12949 21504
rect -8805 21505 -8793 21555
rect -8760 21549 -8256 21555
rect -8760 21511 -8665 21549
rect -8268 21511 -8256 21549
rect -8760 21505 -8256 21511
rect -4878 21549 -4374 21555
rect -4878 21511 -4866 21549
rect -4469 21511 -4374 21549
rect -4878 21505 -4374 21511
rect -4341 21505 -4329 21555
rect -185 21556 -133 21566
rect -4277 21549 -3920 21555
rect -3932 21511 -3920 21549
rect -8857 21494 -8805 21504
rect -4277 21505 -3920 21511
rect -542 21549 -185 21555
rect -88 21555 -38 21594
rect 4248 21555 4298 21671
rect 4343 21556 4395 21566
rect -542 21511 -530 21549
rect -542 21505 -185 21511
rect -4329 21494 -4277 21504
rect -133 21505 -121 21555
rect -88 21549 416 21555
rect -88 21511 7 21549
rect 404 21511 416 21549
rect -88 21505 416 21511
rect 3794 21549 4298 21555
rect 3794 21511 3806 21549
rect 4203 21511 4298 21549
rect 3794 21505 4298 21511
rect 4331 21505 4343 21555
rect 8487 21556 8539 21566
rect 4395 21549 4752 21555
rect 4740 21511 4752 21549
rect -185 21494 -133 21504
rect 4395 21505 4752 21511
rect 8130 21549 8487 21555
rect 8130 21511 8142 21549
rect 8130 21505 8487 21511
rect 4343 21494 4395 21504
rect 8539 21505 8551 21555
rect 8487 21494 8539 21504
rect -13193 21390 -13141 21400
rect -17074 21389 -17064 21390
rect -17349 21383 -17064 21389
rect -16940 21389 -16930 21390
rect -17349 21345 -17337 21383
rect -17349 21339 -17064 21345
rect -17074 21338 -17064 21339
rect -16940 21339 -16928 21389
rect -13550 21383 -13193 21389
rect -8665 21390 -8613 21400
rect -13550 21345 -13538 21383
rect -13550 21339 -13193 21345
rect -16940 21338 -16930 21339
rect -13141 21339 -13129 21389
rect -13096 21383 -12592 21389
rect -13096 21345 -13001 21383
rect -12604 21345 -12592 21383
rect -13096 21339 -12592 21345
rect -9214 21383 -8710 21389
rect -9214 21345 -9202 21383
rect -8805 21345 -8710 21383
rect -9214 21339 -8710 21345
rect -8677 21339 -8665 21389
rect -4521 21390 -4469 21400
rect -8613 21383 -8256 21389
rect -8268 21345 -8256 21383
rect -13193 21328 -13141 21338
rect -17336 21223 -17326 21234
rect -17349 21217 -17326 21223
rect -17254 21223 -17244 21234
rect -13096 21223 -13046 21339
rect -13001 21224 -12949 21234
rect -17254 21217 -16928 21223
rect -17349 21179 -17337 21217
rect -16940 21179 -16928 21217
rect -17349 21173 -17326 21179
rect -17336 21162 -17326 21173
rect -17254 21173 -16928 21179
rect -13550 21217 -13046 21223
rect -13550 21179 -13538 21217
rect -13141 21179 -13046 21217
rect -13550 21173 -13046 21179
rect -13013 21173 -13001 21223
rect -8857 21224 -8805 21234
rect -12949 21217 -12592 21223
rect -12604 21179 -12592 21217
rect -17254 21162 -17244 21173
rect -12949 21173 -12592 21179
rect -9214 21217 -8857 21223
rect -8760 21223 -8710 21339
rect -8613 21339 -8256 21345
rect -4878 21383 -4521 21389
rect 7 21390 59 21400
rect -4878 21345 -4866 21383
rect -4878 21339 -4521 21345
rect -8665 21328 -8613 21338
rect -4469 21339 -4457 21389
rect -4424 21383 -3920 21389
rect -4424 21345 -4329 21383
rect -3932 21345 -3920 21383
rect -4424 21339 -3920 21345
rect -542 21383 -38 21389
rect -542 21345 -530 21383
rect -133 21345 -38 21383
rect -542 21339 -38 21345
rect -5 21339 7 21389
rect 4151 21390 4203 21400
rect 59 21383 416 21389
rect 404 21345 416 21383
rect -4521 21328 -4469 21338
rect -4424 21223 -4374 21339
rect -4329 21224 -4277 21234
rect -9214 21179 -9202 21217
rect -9214 21173 -8857 21179
rect -13001 21162 -12949 21172
rect -8805 21173 -8793 21223
rect -8760 21217 -8256 21223
rect -8760 21179 -8665 21217
rect -8268 21179 -8256 21217
rect -8760 21173 -8256 21179
rect -4878 21217 -4374 21223
rect -4878 21179 -4866 21217
rect -4469 21179 -4374 21217
rect -4878 21173 -4374 21179
rect -4341 21173 -4329 21223
rect -185 21224 -133 21234
rect -4277 21217 -3920 21223
rect -3932 21179 -3920 21217
rect -8857 21162 -8805 21172
rect -4277 21173 -3920 21179
rect -542 21217 -185 21223
rect -88 21223 -38 21339
rect 59 21339 416 21345
rect 3794 21383 4151 21389
rect 8584 21389 8634 21671
rect 3794 21345 3806 21383
rect 3794 21339 4151 21345
rect 7 21328 59 21338
rect 4203 21339 4215 21389
rect 4248 21383 4752 21389
rect 4248 21345 4343 21383
rect 4740 21345 4752 21383
rect 4248 21339 4752 21345
rect 8130 21383 8634 21389
rect 8130 21345 8142 21383
rect 8539 21345 8634 21383
rect 8130 21339 8634 21345
rect 4151 21328 4203 21338
rect 4248 21223 4298 21339
rect 4343 21224 4395 21234
rect -542 21179 -530 21217
rect -542 21173 -185 21179
rect -4329 21162 -4277 21172
rect -133 21173 -121 21223
rect -88 21217 416 21223
rect -88 21179 7 21217
rect 404 21179 416 21217
rect -88 21173 416 21179
rect 3794 21217 4298 21223
rect 3794 21179 3806 21217
rect 4203 21179 4298 21217
rect 3794 21173 4298 21179
rect 4331 21173 4343 21223
rect 8487 21224 8539 21234
rect 4395 21217 4752 21223
rect 4740 21179 4752 21217
rect -185 21162 -133 21172
rect 4395 21173 4752 21179
rect 8130 21217 8487 21223
rect 8130 21179 8142 21217
rect 8130 21173 8487 21179
rect 4343 21162 4395 21172
rect 8539 21173 8551 21223
rect 8487 21162 8539 21172
rect 8662 21057 8668 22501
rect -17466 21051 -16928 21057
rect -17466 21013 -17337 21051
rect -16940 21013 -16928 21051
rect -17466 21007 -16928 21013
rect -13550 21051 -12592 21057
rect -13550 21013 -13538 21051
rect -13141 21013 -13001 21051
rect -12604 21013 -12592 21051
rect -13550 21007 -12592 21013
rect -9214 21051 -8256 21057
rect -9214 21013 -9202 21051
rect -8805 21013 -8665 21051
rect -8268 21013 -8256 21051
rect -9214 21007 -8256 21013
rect -4878 21051 -3920 21057
rect -4878 21013 -4866 21051
rect -4469 21013 -4329 21051
rect -3932 21013 -3920 21051
rect -4878 21007 -3920 21013
rect -542 21051 416 21057
rect -542 21013 -530 21051
rect -133 21013 7 21051
rect 404 21013 416 21051
rect -542 21007 416 21013
rect 3794 21051 4752 21057
rect 3794 21013 3806 21051
rect 4203 21013 4343 21051
rect 4740 21013 4752 21051
rect 3794 21007 4752 21013
rect 8130 21051 8668 21057
rect 8130 21013 8142 21051
rect 8539 21013 8668 21051
rect 8130 21007 8668 21013
rect -17466 20892 -17460 21007
rect 8662 20892 8668 21007
rect -17466 20886 8668 20892
rect 8702 22651 8714 22691
rect 8702 20892 8708 22651
rect 8702 20852 8714 20892
rect -17512 20846 8714 20852
rect -17506 20840 -17460 20846
rect -17402 20218 -16759 20846
rect -13155 20801 -13109 20807
rect -13038 20801 -12065 20846
rect 8662 20840 8708 20846
rect 8647 20801 8693 20807
rect -13161 20795 8699 20801
rect -13161 20755 -13149 20795
rect -17412 20077 -17402 20218
rect -16759 20077 -16749 20218
rect -13155 19343 -13149 20755
rect -13161 19303 -13149 19343
rect -13115 20755 8653 20761
rect -13115 19343 -13109 20755
rect -13013 20655 -12955 20755
rect 8493 20655 8552 20755
rect -13013 20649 -12592 20655
rect -13013 20611 -13001 20649
rect -12604 20611 -12592 20649
rect -13013 20605 -12592 20611
rect -9214 20649 -8256 20655
rect -9214 20611 -9202 20649
rect -8805 20611 -8665 20649
rect -8268 20611 -8256 20649
rect -9214 20605 -8256 20611
rect -4878 20649 -3920 20655
rect -4878 20611 -4866 20649
rect -4469 20611 -4329 20649
rect -3932 20611 -3920 20649
rect -4878 20605 -3920 20611
rect -542 20649 416 20655
rect -542 20611 -530 20649
rect -133 20611 7 20649
rect 404 20611 416 20649
rect -542 20605 416 20611
rect 3794 20649 4752 20655
rect 3794 20611 3806 20649
rect 4203 20611 4343 20649
rect 4740 20611 4752 20649
rect 3794 20605 4752 20611
rect 8130 20650 8552 20655
rect 8130 20649 8551 20650
rect 8130 20611 8142 20649
rect 8539 20611 8551 20649
rect 8130 20605 8551 20611
rect -13013 20489 -12955 20605
rect -13013 20483 -12592 20489
rect -13013 20445 -13001 20483
rect -12604 20445 -12592 20483
rect -13013 20439 -12592 20445
rect -9214 20483 -8256 20489
rect -9214 20445 -9202 20483
rect -8805 20445 -8665 20483
rect -8268 20445 -8256 20483
rect -9214 20439 -8256 20445
rect -4878 20483 -3920 20489
rect -4878 20445 -4866 20483
rect -4469 20445 -4329 20483
rect -3932 20445 -3920 20483
rect -4878 20439 -3920 20445
rect -542 20483 416 20489
rect -542 20445 -530 20483
rect -133 20445 7 20483
rect 404 20445 416 20483
rect -542 20439 416 20445
rect 3794 20483 4752 20489
rect 3794 20445 3806 20483
rect 4203 20445 4343 20483
rect 4740 20445 4752 20483
rect 3794 20439 4752 20445
rect 8130 20483 8551 20489
rect 8130 20445 8142 20483
rect 8539 20445 8551 20483
rect 8130 20439 8551 20445
rect 8501 20323 8551 20439
rect -13013 20317 -12592 20323
rect -13013 20279 -13001 20317
rect -12604 20279 -12592 20317
rect -13013 20273 -12592 20279
rect -9214 20317 -8256 20323
rect -9214 20279 -9202 20317
rect -8805 20279 -8665 20317
rect -8268 20279 -8256 20317
rect -9214 20273 -8256 20279
rect -4878 20317 -3920 20323
rect -4878 20279 -4866 20317
rect -4469 20279 -4329 20317
rect -3932 20279 -3920 20317
rect -4878 20273 -3920 20279
rect -542 20317 416 20323
rect -542 20279 -530 20317
rect -133 20279 7 20317
rect 404 20279 416 20317
rect -542 20273 416 20279
rect 3794 20317 4752 20323
rect 3794 20279 3806 20317
rect 4203 20279 4343 20317
rect 4740 20279 4752 20317
rect 3794 20273 4752 20279
rect 8130 20317 8551 20323
rect 8130 20279 8142 20317
rect 8539 20279 8551 20317
rect 8130 20273 8551 20279
rect -13013 20157 -12963 20273
rect -13013 20151 -12592 20157
rect -13013 20113 -13001 20151
rect -12604 20113 -12592 20151
rect -13013 20107 -12592 20113
rect -9214 20151 -8256 20157
rect -9214 20113 -9202 20151
rect -8805 20113 -8665 20151
rect -8268 20113 -8256 20151
rect -9214 20107 -8256 20113
rect -4878 20151 -3920 20157
rect -4878 20113 -4866 20151
rect -4469 20113 -4329 20151
rect -3932 20113 -3920 20151
rect -4878 20107 -3920 20113
rect -542 20151 416 20157
rect -542 20113 -530 20151
rect -133 20113 7 20151
rect 404 20113 416 20151
rect -542 20107 416 20113
rect 3794 20151 4752 20157
rect 3794 20113 3806 20151
rect 4203 20113 4343 20151
rect 4740 20113 4752 20151
rect 3794 20107 4752 20113
rect 8130 20151 8551 20157
rect 8130 20113 8142 20151
rect 8539 20113 8551 20151
rect 8130 20107 8551 20113
rect -13013 20106 -12963 20107
rect 8501 19991 8551 20107
rect -13013 19985 -12592 19991
rect -13013 19947 -13001 19985
rect -12604 19947 -12592 19985
rect -13013 19941 -12592 19947
rect -9214 19985 -8256 19991
rect -9214 19947 -9202 19985
rect -8805 19947 -8665 19985
rect -8268 19947 -8256 19985
rect -9214 19941 -8256 19947
rect -4878 19985 -3920 19991
rect -4878 19947 -4866 19985
rect -4469 19947 -4329 19985
rect -3932 19947 -3920 19985
rect -4878 19941 -3920 19947
rect -542 19985 416 19991
rect -542 19947 -530 19985
rect -133 19947 7 19985
rect 404 19947 416 19985
rect -542 19941 416 19947
rect 3794 19985 4752 19991
rect 3794 19947 3806 19985
rect 4203 19947 4343 19985
rect 4740 19947 4752 19985
rect 3794 19941 4752 19947
rect 8130 19985 8551 19991
rect 8130 19947 8142 19985
rect 8539 19947 8551 19985
rect 8130 19941 8551 19947
rect -13013 19825 -12963 19941
rect -13013 19819 -12592 19825
rect -13013 19781 -13001 19819
rect -12604 19781 -12592 19819
rect -13013 19775 -12592 19781
rect -9214 19819 -8256 19825
rect -9214 19781 -9202 19819
rect -8805 19781 -8665 19819
rect -8268 19781 -8256 19819
rect -9214 19775 -8256 19781
rect -4878 19819 -3920 19825
rect -4878 19781 -4866 19819
rect -4469 19781 -4329 19819
rect -3932 19781 -3920 19819
rect -4878 19775 -3920 19781
rect -542 19819 416 19825
rect -542 19781 -530 19819
rect -133 19781 7 19819
rect 404 19781 416 19819
rect -542 19775 416 19781
rect 3794 19819 4752 19825
rect 3794 19781 3806 19819
rect 4203 19781 4343 19819
rect 4740 19781 4752 19819
rect 3794 19775 4752 19781
rect 8130 19819 8551 19825
rect 8130 19781 8142 19819
rect 8539 19781 8551 19819
rect 8130 19775 8551 19781
rect -13013 19774 -12963 19775
rect -13011 19659 -13001 19660
rect -13013 19609 -13001 19659
rect -12604 19659 -12594 19660
rect 8501 19659 8551 19775
rect -13011 19608 -13001 19609
rect -12604 19609 -12592 19659
rect -9214 19653 -8256 19659
rect -9214 19615 -9202 19653
rect -8805 19615 -8665 19653
rect -8268 19615 -8256 19653
rect -9214 19609 -8256 19615
rect -4878 19653 -3920 19659
rect -4878 19615 -4866 19653
rect -4469 19615 -4329 19653
rect -3932 19615 -3920 19653
rect -4878 19609 -3920 19615
rect -542 19653 416 19659
rect -542 19615 -530 19653
rect -133 19615 7 19653
rect 404 19615 416 19653
rect -542 19609 416 19615
rect 3794 19653 4752 19659
rect 3794 19615 3806 19653
rect 4203 19615 4343 19653
rect 4740 19615 4752 19653
rect 3794 19609 4752 19615
rect 8130 19653 8551 19659
rect 8130 19615 8142 19653
rect 8539 19615 8551 19653
rect 8130 19609 8551 19615
rect -12604 19608 -12594 19609
rect -13013 19487 -12592 19493
rect -13013 19449 -13001 19487
rect -12604 19449 -12592 19487
rect -13013 19443 -12592 19449
rect -9214 19487 -8256 19493
rect -9214 19449 -9202 19487
rect -8805 19449 -8665 19487
rect -8268 19449 -8256 19487
rect -9214 19443 -8256 19449
rect -4878 19487 -3920 19493
rect -4878 19449 -4866 19487
rect -4469 19449 -4329 19487
rect -3932 19449 -3920 19487
rect -4878 19443 -3920 19449
rect -542 19487 416 19493
rect -542 19449 -530 19487
rect -133 19449 7 19487
rect 404 19449 416 19487
rect -542 19443 416 19449
rect 3794 19487 4752 19493
rect 3794 19449 3806 19487
rect 4203 19449 4343 19487
rect 4740 19449 4752 19487
rect 3794 19443 4752 19449
rect 8130 19487 8551 19493
rect 8130 19449 8142 19487
rect 8539 19449 8551 19487
rect 8130 19443 8551 19449
rect -13013 19343 -12955 19443
rect 8493 19343 8551 19443
rect 8647 19343 8653 20755
rect -13115 19337 8653 19343
rect 8687 20755 8699 20795
rect 8687 19343 8693 20755
rect 8687 19303 8699 19343
rect -13161 19297 8699 19303
rect -13155 19291 -13109 19297
rect 8647 19291 8693 19297
rect -1351 19175 257 19185
rect -7112 19124 -1351 19174
rect -7112 18435 -7062 19124
rect -7029 19091 -6979 19124
rect -4579 19091 -4529 19124
rect -7029 19085 -6608 19091
rect -7029 19047 -7017 19085
rect -6620 19047 -6608 19085
rect -7029 19041 -6608 19047
rect -4950 19085 -4529 19091
rect -4950 19047 -4938 19085
rect -4541 19047 -4529 19085
rect -4950 19041 -4529 19047
rect -4413 19091 -4363 19124
rect -1963 19091 -1913 19124
rect -4413 19085 -3992 19091
rect -4413 19047 -4401 19085
rect -4004 19047 -3992 19085
rect -4413 19041 -3992 19047
rect -2334 19085 -1913 19091
rect -2334 19047 -2322 19085
rect -1925 19047 -1913 19085
rect -2334 19041 -1913 19047
rect -7029 18925 -6979 19041
rect -4579 18925 -4529 19041
rect -1880 18925 -1830 19124
rect -7029 18919 -6608 18925
rect -7029 18881 -7017 18919
rect -6620 18881 -6608 18919
rect -7029 18875 -6608 18881
rect -4950 18919 -4529 18925
rect -4950 18881 -4938 18919
rect -4541 18881 -4529 18919
rect -4950 18875 -4529 18881
rect -4496 18919 -3992 18925
rect -4496 18881 -4401 18919
rect -4004 18881 -3992 18919
rect -4496 18875 -3992 18881
rect -2334 18919 -1830 18925
rect -2334 18881 -2322 18919
rect -1925 18881 -1830 18919
rect -2334 18875 -1830 18881
rect -1797 19091 -1747 19124
rect 1265 19175 2873 19185
rect 257 19124 1265 19174
rect -1351 19113 257 19123
rect 653 19091 703 19124
rect -1797 19085 -1376 19091
rect -1797 19047 -1785 19085
rect -1388 19047 -1376 19085
rect -1797 19041 -1376 19047
rect 282 19085 703 19091
rect 282 19047 294 19085
rect 691 19047 703 19085
rect 282 19041 703 19047
rect 819 19091 869 19124
rect 2873 19124 8634 19174
rect 1265 19113 2873 19123
rect 3269 19091 3319 19124
rect 819 19085 1240 19091
rect 819 19047 831 19085
rect 1228 19047 1240 19085
rect 819 19041 1240 19047
rect 2898 19085 3319 19091
rect 2898 19047 2910 19085
rect 3307 19047 3319 19085
rect 2898 19041 3319 19047
rect -1797 18925 -1747 19041
rect 653 18925 703 19041
rect 3352 18925 3402 19124
rect -1797 18919 -1376 18925
rect -1797 18881 -1785 18919
rect -1388 18881 -1376 18919
rect -1797 18875 -1376 18881
rect 282 18919 703 18925
rect 282 18881 294 18919
rect 691 18881 703 18919
rect 282 18875 703 18881
rect 736 18919 1240 18925
rect 736 18881 831 18919
rect 1228 18881 1240 18919
rect 736 18875 1240 18881
rect 2898 18919 3402 18925
rect 2898 18881 2910 18919
rect 3307 18881 3402 18919
rect 2898 18875 3402 18881
rect 3435 19091 3485 19124
rect 5885 19091 5935 19124
rect 3435 19085 3856 19091
rect 3435 19047 3447 19085
rect 3844 19047 3856 19085
rect 3435 19041 3856 19047
rect 5514 19085 5935 19091
rect 5514 19047 5526 19085
rect 5923 19047 5935 19085
rect 5514 19041 5935 19047
rect 6051 19091 6101 19124
rect 8501 19091 8551 19124
rect 6051 19085 6472 19091
rect 6051 19047 6063 19085
rect 6460 19047 6472 19085
rect 6051 19041 6472 19047
rect 8130 19085 8551 19091
rect 8130 19047 8142 19085
rect 8539 19047 8551 19085
rect 8130 19041 8551 19047
rect 3435 18925 3485 19041
rect 5885 18925 5935 19041
rect 8584 18925 8634 19124
rect 3435 18919 3856 18925
rect 3435 18881 3447 18919
rect 3844 18881 3856 18919
rect 3435 18875 3856 18881
rect 5514 18919 5935 18925
rect 5514 18881 5526 18919
rect 5923 18881 5935 18919
rect 5514 18875 5935 18881
rect 5968 18919 6472 18925
rect 5968 18881 6063 18919
rect 6460 18881 6472 18919
rect 5968 18875 6472 18881
rect 8130 18919 8634 18925
rect 8130 18881 8142 18919
rect 8539 18881 8634 18919
rect 8130 18875 8634 18881
rect -6844 18760 -6792 18770
rect -7029 18753 -6844 18759
rect -4765 18760 -4713 18770
rect -6792 18753 -6608 18759
rect -7029 18715 -7017 18753
rect -6620 18715 -6608 18753
rect -7029 18709 -6844 18715
rect -6792 18709 -6608 18715
rect -4950 18753 -4765 18759
rect -4713 18753 -4529 18759
rect -4950 18715 -4938 18753
rect -4541 18715 -4529 18753
rect -4950 18709 -4765 18715
rect -6844 18698 -6792 18708
rect -4713 18709 -4529 18715
rect -4765 18698 -4713 18708
rect -7017 18594 -6965 18604
rect -7029 18543 -7017 18593
rect -4593 18594 -4541 18604
rect -6965 18587 -6608 18593
rect -6620 18549 -6608 18587
rect -6965 18543 -6608 18549
rect -4950 18587 -4593 18593
rect -4496 18593 -4446 18875
rect -4401 18760 -4349 18770
rect -4413 18709 -4401 18759
rect -1977 18760 -1925 18770
rect -4349 18753 -3992 18759
rect -4004 18715 -3992 18753
rect -4349 18709 -3992 18715
rect -2334 18753 -1977 18759
rect -1880 18759 -1830 18875
rect 736 18759 786 18875
rect 831 18760 883 18770
rect -2334 18715 -2322 18753
rect -2334 18709 -1977 18715
rect -4401 18698 -4349 18708
rect -1925 18709 -1913 18759
rect -1880 18753 -1376 18759
rect -1880 18715 -1785 18753
rect -1388 18715 -1376 18753
rect -1880 18709 -1376 18715
rect 282 18753 786 18759
rect 282 18715 294 18753
rect 691 18715 786 18753
rect 282 18709 786 18715
rect 819 18709 831 18759
rect 3255 18760 3307 18770
rect 883 18753 1240 18759
rect 1228 18715 1240 18753
rect -1977 18698 -1925 18708
rect -1880 18593 -1830 18709
rect -1785 18594 -1733 18604
rect -4950 18549 -4938 18587
rect -4950 18543 -4593 18549
rect -7017 18532 -6965 18542
rect -4541 18543 -4529 18593
rect -4496 18587 -3992 18593
rect -4496 18549 -4401 18587
rect -4004 18549 -3992 18587
rect -4496 18543 -3992 18549
rect -2334 18587 -1830 18593
rect -2334 18549 -2322 18587
rect -1925 18549 -1830 18587
rect -2334 18543 -1830 18549
rect -1797 18543 -1785 18593
rect 639 18594 691 18604
rect -1733 18587 -1376 18593
rect -1388 18549 -1376 18587
rect -4593 18532 -4541 18542
rect -7744 18369 -7734 18435
rect -7668 18421 -6604 18435
rect -4496 18427 -4446 18543
rect -4401 18428 -4349 18438
rect -7668 18383 -7017 18421
rect -6620 18383 -6604 18421
rect -7668 18369 -6604 18383
rect -4950 18421 -4446 18427
rect -4950 18383 -4938 18421
rect -4541 18383 -4446 18421
rect -4950 18377 -4446 18383
rect -4413 18377 -4401 18427
rect -1977 18428 -1925 18438
rect -4349 18421 -3992 18427
rect -4004 18383 -3992 18421
rect -7112 18095 -7062 18369
rect -7017 18262 -6965 18272
rect -7029 18211 -7017 18261
rect -4593 18262 -4541 18272
rect -6965 18255 -6608 18261
rect -6620 18217 -6608 18255
rect -6965 18211 -6608 18217
rect -4950 18255 -4593 18261
rect -4496 18261 -4446 18377
rect -4349 18377 -3992 18383
rect -2334 18421 -1977 18427
rect -1880 18427 -1830 18543
rect -1733 18543 -1376 18549
rect 282 18587 639 18593
rect 736 18593 786 18709
rect 883 18709 1240 18715
rect 2898 18753 3255 18759
rect 3352 18759 3402 18875
rect 5968 18759 6018 18875
rect 6063 18760 6115 18770
rect 2898 18715 2910 18753
rect 2898 18709 3255 18715
rect 831 18698 883 18708
rect 3307 18709 3319 18759
rect 3352 18753 3856 18759
rect 3352 18715 3447 18753
rect 3844 18715 3856 18753
rect 3352 18709 3856 18715
rect 5514 18753 6018 18759
rect 5514 18715 5526 18753
rect 5923 18715 6018 18753
rect 5514 18709 6018 18715
rect 6051 18709 6063 18759
rect 8487 18760 8539 18770
rect 6115 18753 6472 18759
rect 6460 18715 6472 18753
rect 3255 18698 3307 18708
rect 3352 18593 3402 18709
rect 3447 18594 3499 18604
rect 282 18549 294 18587
rect 282 18543 639 18549
rect -1785 18532 -1733 18542
rect 691 18543 703 18593
rect 736 18587 1240 18593
rect 736 18549 831 18587
rect 1228 18549 1240 18587
rect 736 18543 1240 18549
rect 2898 18587 3402 18593
rect 2898 18549 2910 18587
rect 3307 18549 3402 18587
rect 2898 18543 3402 18549
rect 3435 18543 3447 18593
rect 5871 18594 5923 18604
rect 3499 18587 3856 18593
rect 3844 18549 3856 18587
rect 639 18532 691 18542
rect 736 18427 786 18543
rect 831 18428 883 18438
rect -2334 18383 -2322 18421
rect -2334 18377 -1977 18383
rect -4401 18366 -4349 18376
rect -1925 18377 -1913 18427
rect -1880 18421 -1376 18427
rect -1880 18383 -1785 18421
rect -1388 18383 -1376 18421
rect -1880 18377 -1376 18383
rect 282 18421 786 18427
rect 282 18383 294 18421
rect 691 18383 786 18421
rect 282 18377 786 18383
rect 819 18377 831 18427
rect 3255 18428 3307 18438
rect 883 18421 1240 18427
rect 1228 18383 1240 18421
rect -1977 18366 -1925 18376
rect -1880 18261 -1830 18377
rect -1785 18262 -1733 18272
rect -4950 18217 -4938 18255
rect -4950 18211 -4593 18217
rect -7017 18200 -6965 18210
rect -4541 18211 -4529 18261
rect -4496 18255 -3992 18261
rect -4496 18217 -4401 18255
rect -4004 18217 -3992 18255
rect -4496 18211 -3992 18217
rect -2334 18255 -1830 18261
rect -2334 18217 -2322 18255
rect -1925 18217 -1830 18255
rect -2334 18211 -1830 18217
rect -1797 18211 -1785 18261
rect 639 18262 691 18272
rect -1733 18255 -1376 18261
rect -1388 18217 -1376 18255
rect -4593 18200 -4541 18210
rect -4496 18095 -4446 18211
rect -1880 18095 -1830 18211
rect -1733 18211 -1376 18217
rect 282 18255 639 18261
rect 736 18261 786 18377
rect 883 18377 1240 18383
rect 2898 18421 3255 18427
rect 3352 18427 3402 18543
rect 3499 18543 3856 18549
rect 5514 18587 5871 18593
rect 5968 18593 6018 18709
rect 6115 18709 6472 18715
rect 8130 18753 8487 18759
rect 8130 18715 8142 18753
rect 8130 18709 8487 18715
rect 6063 18698 6115 18708
rect 8539 18709 8551 18759
rect 8487 18698 8539 18708
rect 8584 18593 8634 18875
rect 5514 18549 5526 18587
rect 5514 18543 5871 18549
rect 3447 18532 3499 18542
rect 5923 18543 5935 18593
rect 5968 18587 6472 18593
rect 5968 18549 6063 18587
rect 6460 18549 6472 18587
rect 5968 18543 6472 18549
rect 8130 18587 8634 18593
rect 8130 18549 8142 18587
rect 8539 18549 8634 18587
rect 8130 18543 8634 18549
rect 5871 18532 5923 18542
rect 5968 18427 6018 18543
rect 6063 18428 6115 18438
rect 2898 18383 2910 18421
rect 2898 18377 3255 18383
rect 831 18366 883 18376
rect 3307 18377 3319 18427
rect 3352 18421 3856 18427
rect 3352 18383 3447 18421
rect 3844 18383 3856 18421
rect 3352 18377 3856 18383
rect 5514 18421 6018 18427
rect 5514 18383 5526 18421
rect 5923 18383 6018 18421
rect 5514 18377 6018 18383
rect 6051 18377 6063 18427
rect 8487 18428 8539 18438
rect 6115 18421 6472 18427
rect 6460 18383 6472 18421
rect 3255 18366 3307 18376
rect 3352 18261 3402 18377
rect 3447 18262 3499 18272
rect 282 18217 294 18255
rect 282 18211 639 18217
rect -1785 18200 -1733 18210
rect 691 18211 703 18261
rect 736 18255 1240 18261
rect 736 18217 831 18255
rect 1228 18217 1240 18255
rect 736 18211 1240 18217
rect 2898 18255 3402 18261
rect 2898 18217 2910 18255
rect 3307 18217 3402 18255
rect 2898 18211 3402 18217
rect 3435 18211 3447 18261
rect 5871 18262 5923 18272
rect 3499 18255 3856 18261
rect 3844 18217 3856 18255
rect 639 18200 691 18210
rect 736 18095 786 18211
rect 3352 18095 3402 18211
rect 3499 18211 3856 18217
rect 5514 18255 5871 18261
rect 5514 18217 5526 18255
rect 5514 18211 5871 18217
rect 3447 18200 3499 18210
rect 5923 18211 5935 18261
rect 5871 18200 5923 18210
rect 5968 18095 6018 18377
rect 6115 18377 6472 18383
rect 8130 18421 8487 18427
rect 8130 18383 8142 18421
rect 8130 18377 8487 18383
rect 6063 18366 6115 18376
rect 8539 18377 8551 18427
rect 8487 18366 8539 18376
rect 6236 18262 6288 18272
rect 6051 18255 6236 18261
rect 8315 18262 8367 18272
rect 6288 18255 6472 18261
rect 6051 18217 6063 18255
rect 6460 18217 6472 18255
rect 6051 18211 6236 18217
rect 6288 18211 6472 18217
rect 8130 18255 8315 18261
rect 8367 18255 8551 18261
rect 8130 18217 8142 18255
rect 8539 18217 8551 18255
rect 8130 18211 8315 18217
rect 6236 18200 6288 18210
rect 8367 18211 8551 18217
rect 8315 18200 8367 18210
rect -7112 18089 -6608 18095
rect -7112 18051 -7017 18089
rect -6620 18051 -6608 18089
rect -7112 18045 -6608 18051
rect -4950 18089 -4446 18095
rect -4950 18051 -4938 18089
rect -4541 18051 -4446 18089
rect -4950 18045 -4446 18051
rect -7017 17930 -6965 17940
rect -7029 17879 -7017 17929
rect -4593 17930 -4541 17940
rect -6965 17923 -6608 17929
rect -6620 17885 -6608 17923
rect -6965 17879 -6608 17885
rect -4950 17923 -4593 17929
rect -4950 17885 -4938 17923
rect -4950 17879 -4593 17885
rect -7017 17868 -6965 17878
rect -4541 17879 -4529 17929
rect -4593 17868 -4541 17878
rect -4496 17846 -4446 18045
rect -4413 18089 -3992 18095
rect -4413 18051 -4401 18089
rect -4004 18051 -3992 18089
rect -4413 18045 -3992 18051
rect -2334 18089 -1913 18095
rect -2334 18051 -2322 18089
rect -1925 18051 -1913 18089
rect -2334 18045 -1913 18051
rect -1880 18089 -1376 18095
rect -1880 18051 -1785 18089
rect -1388 18051 -1376 18089
rect -1880 18045 -1376 18051
rect 282 18089 786 18095
rect 282 18051 294 18089
rect 691 18051 786 18089
rect 282 18045 786 18051
rect -4413 17929 -4363 18045
rect -1963 17929 -1913 18045
rect -4413 17923 -3992 17929
rect -4413 17885 -4401 17923
rect -4004 17885 -3992 17923
rect -4413 17879 -3992 17885
rect -2334 17923 -1913 17929
rect -2334 17885 -2322 17923
rect -1925 17885 -1913 17923
rect -2334 17879 -1913 17885
rect -4413 17846 -4363 17879
rect -2178 17846 -2044 17879
rect -1963 17846 -1913 17879
rect -1797 17923 -1376 17929
rect -1797 17885 -1785 17923
rect -1388 17885 -1376 17923
rect -1797 17879 -1376 17885
rect 282 17923 703 17929
rect 282 17885 294 17923
rect 691 17885 703 17923
rect 282 17879 703 17885
rect -1797 17846 -1747 17879
rect 653 17846 703 17879
rect 736 17846 786 18045
rect 819 18089 1240 18095
rect 819 18051 831 18089
rect 1228 18051 1240 18089
rect 819 18045 1240 18051
rect 2898 18089 3319 18095
rect 2898 18051 2910 18089
rect 3307 18051 3319 18089
rect 2898 18045 3319 18051
rect 3352 18089 3856 18095
rect 3352 18051 3447 18089
rect 3844 18051 3856 18089
rect 3352 18045 3856 18051
rect 5514 18089 6472 18095
rect 5514 18051 5526 18089
rect 5923 18051 6063 18089
rect 6460 18051 6472 18089
rect 5514 18045 6472 18051
rect 8130 18089 8551 18095
rect 8130 18051 8142 18089
rect 8539 18051 8551 18089
rect 8130 18045 8551 18051
rect 819 17929 869 18045
rect 3269 17929 3319 18045
rect 5968 18012 6018 18045
rect 8501 18012 8551 18045
rect 5968 17962 8551 18012
rect 5968 17929 6018 17962
rect 8501 17929 8551 17962
rect 819 17923 1240 17929
rect 819 17885 831 17923
rect 1228 17885 1240 17923
rect 819 17879 1240 17885
rect 2898 17923 3319 17929
rect 2898 17885 2910 17923
rect 3307 17885 3319 17923
rect 2898 17879 3319 17885
rect 819 17846 869 17879
rect 3269 17846 3319 17879
rect 3435 17923 3856 17929
rect 3435 17885 3447 17923
rect 3844 17885 3856 17923
rect 3435 17879 3856 17885
rect 5514 17923 5935 17929
rect 5514 17885 5526 17923
rect 5923 17885 5935 17923
rect 5514 17879 5935 17885
rect 3435 17846 3485 17879
rect 5885 17846 5935 17879
rect 5968 17923 6472 17929
rect 5968 17885 6063 17923
rect 6460 17885 6472 17923
rect 5968 17879 6472 17885
rect 8130 17923 8551 17929
rect 8130 17885 8142 17923
rect 8539 17885 8551 17923
rect 8130 17879 8551 17885
rect 5968 17846 6018 17879
rect -4496 17796 6018 17846
rect -16705 17647 -16659 17653
rect -14377 17647 -14331 17653
rect -12319 17647 -12273 17653
rect -10261 17647 -10215 17653
rect -7941 17647 -7895 17653
rect -16711 17641 -7889 17647
rect -16711 17601 -16699 17641
rect -16705 15704 -16699 17601
rect -16711 15664 -16699 15704
rect -16665 17601 -7935 17607
rect -16665 15704 -16659 17601
rect -16523 17547 -16477 17559
rect -16523 17513 -16517 17547
rect -16483 17513 -16477 17547
rect -16523 17466 -16477 17513
rect -16523 17454 -16389 17466
rect -14377 17454 -14331 17601
rect -12319 17454 -12273 17601
rect -10261 17454 -10215 17601
rect -8115 17547 -8069 17559
rect -8115 17513 -8109 17547
rect -8075 17513 -8069 17547
rect -8115 17466 -8069 17513
rect -8209 17454 -8069 17466
rect -16523 17278 -16517 17454
rect -16483 17278 -16438 17454
rect -16386 17278 -16376 17454
rect -14390 17278 -14380 17454
rect -14328 17278 -14318 17454
rect -12319 17278 -12313 17454
rect -12279 17278 -12273 17454
rect -10274 17278 -10264 17454
rect -10212 17278 -10202 17454
rect -8216 17278 -8206 17454
rect -8154 17278 -8109 17454
rect -8075 17278 -8069 17454
rect -16523 17266 -16389 17278
rect -14377 17266 -14331 17278
rect -12319 17225 -12273 17278
rect -10261 17266 -10215 17278
rect -8209 17266 -8069 17278
rect -15887 17219 -14879 17225
rect -15887 17185 -15875 17219
rect -14891 17185 -14879 17219
rect -15887 17151 -14879 17185
rect -13829 17219 -10763 17225
rect -13829 17185 -13817 17219
rect -12833 17185 -11759 17219
rect -10775 17185 -10763 17219
rect -13829 17179 -10763 17185
rect -9713 17219 -8705 17225
rect -9713 17185 -9701 17219
rect -8717 17185 -8705 17219
rect -9713 17151 -8705 17185
rect -16611 17105 -7981 17151
rect -16611 16783 -16565 17105
rect -15885 17074 -15875 17077
rect -15887 17028 -15875 17074
rect -14891 17074 -14881 17077
rect -9711 17074 -9701 17077
rect -14891 17068 -9701 17074
rect -8717 17074 -8707 17077
rect -14891 17034 -13817 17068
rect -12833 17034 -11759 17068
rect -10775 17034 -9701 17068
rect -15885 17025 -15875 17028
rect -14891 17028 -9701 17034
rect -14891 17025 -14881 17028
rect -9711 17025 -9701 17028
rect -8717 17028 -8705 17074
rect -8717 17025 -8707 17028
rect -16523 16975 -16477 16987
rect -16435 16975 -16389 16987
rect -14377 16975 -14331 16987
rect -12319 16975 -12273 16987
rect -10261 16975 -10215 16987
rect -8203 16975 -8157 16987
rect -16527 16799 -16517 16975
rect -16395 16799 -16385 16975
rect -14390 16799 -14380 16975
rect -14328 16799 -14318 16975
rect -12332 16799 -12322 16975
rect -12270 16799 -12260 16975
rect -10274 16799 -10264 16975
rect -10212 16799 -10202 16975
rect -8203 16799 -8197 16975
rect -8163 16799 -8157 16975
rect -16620 16777 -16556 16783
rect -16620 16725 -16614 16777
rect -16562 16725 -16556 16777
rect -16620 16719 -16556 16725
rect -16523 16678 -16477 16799
rect -16435 16678 -16389 16799
rect -14377 16787 -14331 16799
rect -12319 16787 -12273 16799
rect -10261 16787 -10215 16799
rect -15887 16740 -14879 16746
rect -15887 16706 -15875 16740
rect -14891 16706 -14879 16740
rect -16523 16669 -16438 16678
rect -16523 16635 -16517 16669
rect -16483 16635 -16438 16669
rect -16523 16626 -16438 16635
rect -16386 16626 -16376 16678
rect -15887 16669 -14879 16706
rect -13829 16740 -12821 16746
rect -13829 16706 -13817 16740
rect -12833 16706 -12821 16740
rect -13829 16700 -12821 16706
rect -11771 16740 -10763 16746
rect -11771 16706 -11759 16740
rect -10775 16706 -10763 16740
rect -11771 16700 -10763 16706
rect -9713 16740 -8705 16746
rect -9713 16706 -9701 16740
rect -8717 16706 -8705 16740
rect -9713 16669 -8705 16706
rect -8203 16678 -8157 16799
rect -8115 16975 -8069 16987
rect -8115 16799 -8109 16975
rect -8075 16799 -8069 16975
rect -8115 16678 -8069 16799
rect -8027 16783 -7981 17105
rect -8036 16777 -7972 16783
rect -8036 16725 -8030 16777
rect -7978 16725 -7972 16777
rect -8036 16719 -7972 16725
rect -15887 16635 -8705 16669
rect -16620 16579 -16556 16585
rect -16620 16527 -16614 16579
rect -16562 16527 -16556 16579
rect -16620 16521 -16556 16527
rect -16611 16199 -16565 16521
rect -16523 16505 -16477 16626
rect -16523 16329 -16517 16505
rect -16483 16329 -16477 16505
rect -16523 16317 -16477 16329
rect -16435 16505 -16389 16626
rect -15887 16598 -14879 16635
rect -15887 16564 -15875 16598
rect -14891 16564 -14879 16598
rect -15887 16558 -14879 16564
rect -13829 16598 -12821 16604
rect -13829 16564 -13817 16598
rect -12833 16564 -12821 16598
rect -13829 16558 -12821 16564
rect -11771 16598 -10763 16604
rect -11771 16564 -11759 16598
rect -10775 16564 -10763 16598
rect -11771 16558 -10763 16564
rect -9713 16598 -8705 16635
rect -8216 16626 -8206 16678
rect -8154 16669 -8069 16678
rect -8154 16635 -8109 16669
rect -8075 16635 -8069 16669
rect -8154 16626 -8069 16635
rect -9713 16564 -9701 16598
rect -8717 16564 -8705 16598
rect -9713 16558 -8705 16564
rect -14377 16505 -14331 16517
rect -12319 16505 -12273 16517
rect -10261 16505 -10215 16517
rect -8203 16505 -8157 16626
rect -16435 16329 -16429 16505
rect -16395 16329 -16389 16505
rect -14390 16329 -14380 16505
rect -14328 16329 -14318 16505
rect -12332 16329 -12322 16505
rect -12270 16329 -12260 16505
rect -10274 16329 -10264 16505
rect -10212 16329 -10202 16505
rect -8203 16329 -8197 16505
rect -8163 16329 -8157 16505
rect -16435 16317 -16389 16329
rect -14377 16317 -14331 16329
rect -12319 16317 -12273 16329
rect -10261 16317 -10215 16329
rect -8203 16317 -8157 16329
rect -8115 16505 -8069 16626
rect -8036 16579 -7972 16585
rect -8036 16527 -8030 16579
rect -7978 16527 -7972 16579
rect -8036 16521 -7972 16527
rect -8115 16329 -8109 16505
rect -8075 16329 -8069 16505
rect -8027 16397 -7981 16521
rect -8030 16391 -7978 16397
rect -8030 16333 -7978 16339
rect -8115 16317 -8069 16329
rect -15885 16276 -15875 16279
rect -15887 16230 -15875 16276
rect -14891 16276 -14881 16279
rect -9711 16276 -9701 16279
rect -14891 16270 -9701 16276
rect -8717 16276 -8707 16279
rect -14891 16236 -13817 16270
rect -12833 16236 -11759 16270
rect -10775 16236 -9701 16270
rect -15885 16227 -15875 16230
rect -14891 16230 -9701 16236
rect -14891 16227 -14881 16230
rect -9711 16227 -9701 16230
rect -8717 16230 -8705 16276
rect -8717 16227 -8707 16230
rect -8027 16199 -7981 16333
rect -16611 16153 -7981 16199
rect -15887 16119 -14879 16153
rect -15887 16085 -15875 16119
rect -14891 16085 -14879 16119
rect -15887 16079 -14879 16085
rect -13829 16119 -10763 16125
rect -13829 16085 -13817 16119
rect -12833 16085 -11759 16119
rect -10775 16085 -10763 16119
rect -13829 16079 -10763 16085
rect -9713 16119 -8705 16153
rect -9713 16085 -9701 16119
rect -8717 16085 -8705 16119
rect -9713 16079 -8705 16085
rect -16523 16026 -16389 16038
rect -14377 16026 -14331 16038
rect -12319 16026 -12273 16079
rect -10261 16026 -10215 16038
rect -8203 16026 -8069 16038
rect -16523 15850 -16517 16026
rect -16483 15850 -16438 16026
rect -16386 15850 -16376 16026
rect -14390 15850 -14380 16026
rect -14328 15850 -14318 16026
rect -12319 15850 -12313 16026
rect -12279 15850 -12273 16026
rect -10274 15850 -10264 16026
rect -10212 15850 -10202 16026
rect -8216 15850 -8206 16026
rect -8154 15850 -8109 16026
rect -8075 15850 -8069 16026
rect -16523 15838 -16389 15850
rect -16523 15791 -16477 15838
rect -16523 15757 -16517 15791
rect -16483 15757 -16477 15791
rect -16523 15745 -16477 15757
rect -14377 15704 -14331 15850
rect -12319 15704 -12273 15850
rect -10261 15704 -10215 15850
rect -8203 15838 -8069 15850
rect -8115 15791 -8069 15838
rect -8115 15757 -8109 15791
rect -8075 15757 -8069 15791
rect -8115 15745 -8069 15757
rect -7941 15704 -7935 17601
rect -16665 15698 -7935 15704
rect -7901 17601 -7889 17641
rect -7901 15704 -7895 17601
rect -7676 17558 -7630 17564
rect -5356 17558 -5310 17564
rect -3036 17558 -2990 17564
rect -7682 17552 -2984 17558
rect -7682 17512 -7670 17552
rect -7901 15685 -7889 15704
rect -7676 15698 -7670 17512
rect -7682 15685 -7670 15698
rect -7636 17512 -3030 17518
rect -7636 15698 -7630 17512
rect -7502 17453 -7456 17465
rect -7502 17419 -7496 17453
rect -7462 17419 -7456 17453
rect -7502 17372 -7456 17419
rect -7502 17360 -7368 17372
rect -5356 17360 -5310 17512
rect -3210 17453 -3164 17465
rect -3210 17419 -3204 17453
rect -3170 17419 -3164 17453
rect -3298 17360 -3252 17372
rect -7502 17184 -7496 17360
rect -7462 17184 -7417 17360
rect -7365 17184 -7355 17360
rect -5369 17184 -5359 17360
rect -5307 17184 -5297 17360
rect -3298 17184 -3292 17360
rect -3258 17184 -3252 17360
rect -7502 17172 -7368 17184
rect -5356 17172 -5310 17184
rect -3298 17131 -3252 17184
rect -3210 17360 -3164 17419
rect -3210 17184 -3204 17360
rect -3170 17184 -3164 17360
rect -3210 17131 -3164 17184
rect -7589 17125 -3077 17131
rect -7589 17091 -6854 17125
rect -5870 17091 -4796 17125
rect -3812 17091 -3077 17125
rect -7589 17085 -3077 17091
rect -7589 16726 -7543 17085
rect -7502 17021 -7456 17033
rect -7502 16987 -7496 17021
rect -7462 16987 -7456 17021
rect -7502 16940 -7456 16987
rect -3210 17021 -3164 17033
rect -3210 16987 -3204 17021
rect -3170 16987 -3164 17021
rect -3210 16940 -3164 16987
rect -7502 16928 -7368 16940
rect -5356 16928 -5310 16940
rect -3298 16928 -3164 16940
rect -7502 16752 -7496 16928
rect -7462 16752 -7408 16928
rect -7374 16752 -7368 16928
rect -5369 16752 -5359 16928
rect -5307 16752 -5297 16928
rect -3311 16752 -3301 16928
rect -3249 16752 -3204 16928
rect -3170 16752 -3164 16928
rect -7502 16740 -7368 16752
rect -5356 16740 -5310 16752
rect -3298 16740 -3164 16752
rect -7598 16720 -7534 16726
rect -7598 16668 -7592 16720
rect -7540 16668 -7534 16720
rect -7598 16662 -7534 16668
rect -7414 16628 -7368 16740
rect -3123 16726 -3077 17085
rect -3132 16720 -3068 16726
rect -6866 16693 -5858 16699
rect -6866 16659 -6854 16693
rect -5870 16659 -5858 16693
rect -6866 16628 -5858 16659
rect -4808 16693 -3800 16699
rect -4808 16659 -4796 16693
rect -3812 16659 -3800 16693
rect -3132 16668 -3126 16720
rect -3074 16668 -3068 16720
rect -3132 16662 -3068 16668
rect -4808 16628 -3800 16659
rect -7414 16582 -3252 16628
rect -6866 16551 -5858 16582
rect -7598 16542 -7534 16548
rect -7598 16490 -7592 16542
rect -7540 16490 -7534 16542
rect -6866 16517 -6854 16551
rect -5870 16517 -5858 16551
rect -6866 16511 -5858 16517
rect -4808 16551 -3800 16582
rect -4808 16517 -4796 16551
rect -3812 16517 -3800 16551
rect -4808 16511 -3800 16517
rect -7598 16484 -7534 16490
rect -7589 16125 -7543 16484
rect -3298 16470 -3252 16582
rect -3132 16542 -3068 16548
rect -3132 16490 -3126 16542
rect -3074 16490 -3068 16542
rect -3132 16484 -3068 16490
rect -7502 16458 -7368 16470
rect -5356 16458 -5310 16470
rect -3298 16458 -3164 16470
rect -7502 16282 -7496 16458
rect -7462 16282 -7417 16458
rect -7365 16282 -7355 16458
rect -5369 16282 -5359 16458
rect -5307 16282 -5297 16458
rect -3302 16282 -3292 16458
rect -3240 16282 -3204 16458
rect -3170 16282 -3164 16458
rect -7502 16270 -7368 16282
rect -5356 16270 -5310 16282
rect -3298 16270 -3164 16282
rect -7502 16223 -7456 16270
rect -7502 16189 -7496 16223
rect -7462 16189 -7456 16223
rect -7502 16177 -7456 16189
rect -3210 16223 -3164 16270
rect -3210 16189 -3204 16223
rect -3170 16189 -3164 16223
rect -3210 16177 -3164 16189
rect -3123 16125 -3077 16484
rect -7589 16119 -3077 16125
rect -7589 16085 -6854 16119
rect -5870 16085 -4796 16119
rect -3812 16085 -3077 16119
rect -7589 16079 -3077 16085
rect -7502 16026 -7456 16079
rect -7502 15850 -7496 16026
rect -7462 15850 -7456 16026
rect -7502 15791 -7456 15850
rect -7414 16026 -7368 16079
rect -5356 16026 -5310 16038
rect -3298 16026 -3164 16038
rect -7414 15850 -7408 16026
rect -7374 15850 -7368 16026
rect -5369 15850 -5359 16026
rect -5307 15850 -5297 16026
rect -3311 15850 -3301 16026
rect -3249 15850 -3204 16026
rect -3170 15850 -3164 16026
rect -7414 15838 -7368 15850
rect -7502 15757 -7496 15791
rect -7462 15757 -7456 15791
rect -7502 15745 -7456 15757
rect -5356 15698 -5310 15850
rect -3298 15838 -3164 15850
rect -3210 15791 -3164 15838
rect -3210 15757 -3204 15791
rect -3170 15757 -3164 15791
rect -3210 15745 -3164 15757
rect -3036 15698 -3030 17512
rect -7636 15692 -3030 15698
rect -2996 17512 -2984 17552
rect -2996 15698 -2990 17512
rect -2178 17409 -2044 17796
rect -215 17627 -169 17633
rect 4272 17627 4318 17633
rect 8647 17627 8693 17633
rect -221 17621 8699 17627
rect -1276 17614 -1230 17620
rect -384 17614 -338 17620
rect -1282 17608 -332 17614
rect -1282 17568 -1270 17608
rect -2188 17275 -2178 17409
rect -2044 17275 -2034 17409
rect -1276 16826 -1270 17568
rect -1282 16786 -1270 16826
rect -1236 17568 -378 17574
rect -1236 16826 -1230 17568
rect -1176 17524 -1130 17536
rect -1176 17490 -1170 17524
rect -1136 17490 -1130 17524
rect -1176 17452 -1130 17490
rect -990 17524 -882 17530
rect -990 17490 -978 17524
rect -894 17490 -882 17524
rect -990 17484 -882 17490
rect -1176 17440 -1042 17452
rect -1176 17264 -1170 17440
rect -1136 17264 -1082 17440
rect -1048 17264 -1042 17440
rect -1176 17252 -1042 17264
rect -1088 17223 -1042 17252
rect -830 17440 -784 17568
rect -732 17524 -624 17530
rect -732 17490 -720 17524
rect -636 17490 -624 17524
rect -732 17484 -624 17490
rect -484 17524 -438 17536
rect -484 17490 -478 17524
rect -444 17490 -438 17524
rect -484 17452 -438 17490
rect -830 17264 -824 17440
rect -790 17264 -784 17440
rect -1101 17171 -1091 17223
rect -1039 17171 -1029 17223
rect -990 17214 -882 17221
rect -990 17180 -978 17214
rect -894 17180 -882 17214
rect -990 17174 -882 17180
rect -1088 17142 -1042 17171
rect -1176 17130 -1042 17142
rect -1176 16954 -1170 17130
rect -1136 16954 -1082 17130
rect -1048 16954 -1042 17130
rect -1176 16942 -1042 16954
rect -830 17130 -784 17264
rect -572 17440 -438 17452
rect -572 17264 -566 17440
rect -532 17264 -478 17440
rect -444 17264 -438 17440
rect -572 17252 -438 17264
rect -572 17223 -526 17252
rect -732 17214 -624 17220
rect -732 17180 -720 17214
rect -636 17180 -624 17214
rect -732 17174 -624 17180
rect -585 17171 -575 17223
rect -523 17171 -513 17223
rect -830 16954 -824 17130
rect -790 16954 -784 17130
rect -1176 16904 -1130 16942
rect -988 16910 -978 16913
rect -1176 16870 -1170 16904
rect -1136 16870 -1130 16904
rect -1176 16858 -1130 16870
rect -990 16864 -978 16910
rect -894 16910 -884 16913
rect -988 16861 -978 16864
rect -894 16864 -882 16910
rect -894 16861 -884 16864
rect -830 16826 -784 16954
rect -572 17142 -526 17171
rect -572 17130 -438 17142
rect -572 16954 -566 17130
rect -532 16954 -478 17130
rect -444 16954 -438 17130
rect -572 16942 -438 16954
rect -732 16904 -624 16910
rect -732 16870 -720 16904
rect -636 16870 -624 16904
rect -732 16864 -624 16870
rect -484 16904 -438 16942
rect -484 16870 -478 16904
rect -444 16870 -438 16904
rect -484 16858 -438 16870
rect -384 16826 -378 17568
rect -1236 16820 -378 16826
rect -344 17568 -332 17608
rect -221 17581 -209 17621
rect -344 16826 -338 17568
rect -344 16786 -332 16826
rect -1282 16780 -332 16786
rect -1276 16774 -1230 16780
rect -384 16774 -338 16780
rect -215 15965 -209 17581
rect -221 15925 -209 15965
rect -175 17581 8653 17587
rect -175 15965 -169 17581
rect -98 17536 -52 17548
rect -98 17502 -92 17536
rect -58 17502 -52 17536
rect -98 17464 -52 17502
rect -98 17452 148 17464
rect 4160 17452 4206 17464
rect 4272 17452 4318 17581
rect 7289 17542 8370 17543
rect 5320 17536 8370 17542
rect 5320 17502 5332 17536
rect 7316 17502 8370 17536
rect 5320 17497 8370 17502
rect 5320 17496 7328 17497
rect 8336 17464 8370 17497
rect 8530 17536 8576 17548
rect 8530 17502 8536 17536
rect 8570 17502 8576 17536
rect 8530 17464 8576 17502
rect -98 17276 -92 17452
rect -58 17276 -4 17452
rect 30 17276 43 17452
rect 95 17276 108 17452
rect 142 17276 148 17452
rect 4141 17276 4151 17452
rect 4215 17276 4225 17452
rect 4272 17276 4278 17452
rect 4312 17276 4318 17452
rect -98 17264 148 17276
rect 4160 17264 4206 17276
rect -98 17142 -52 17154
rect -98 17108 -92 17142
rect -58 17108 -52 17142
rect -98 17070 -52 17108
rect 4272 17070 4318 17276
rect 8330 17452 8576 17464
rect 8330 17276 8336 17452
rect 8370 17276 8448 17452
rect 8482 17276 8536 17452
rect 8570 17276 8576 17452
rect 8330 17264 8576 17276
rect 8530 17142 8576 17154
rect 8530 17108 8536 17142
rect 8570 17108 8576 17142
rect 8530 17070 8576 17108
rect -98 17058 148 17070
rect -98 16882 -92 17058
rect -58 16882 -4 17058
rect 30 16882 43 17058
rect 95 16882 108 17058
rect 142 16882 148 17058
rect -98 16870 148 16882
rect 4160 17058 4318 17070
rect 4160 16882 4166 17058
rect 4200 16882 4278 17058
rect 4312 16882 4318 17058
rect 4160 16870 4318 16882
rect 8330 17058 8576 17070
rect 8330 16882 8336 17058
rect 8370 16882 8383 17058
rect 8435 16882 8448 17058
rect 8482 16882 8536 17058
rect 8570 16882 8576 17058
rect 8330 16870 8576 16882
rect 4161 16676 4318 16870
rect -98 16664 148 16676
rect -98 16488 -92 16664
rect -58 16488 -4 16664
rect 30 16488 43 16664
rect 95 16488 108 16664
rect 142 16488 148 16664
rect -98 16476 148 16488
rect 4160 16664 4318 16676
rect 4160 16488 4166 16664
rect 4200 16488 4278 16664
rect 4312 16488 4318 16664
rect 4160 16476 4318 16488
rect 8330 16664 8576 16676
rect 8330 16488 8336 16664
rect 8370 16488 8383 16664
rect 8435 16488 8448 16664
rect 8482 16488 8536 16664
rect 8570 16488 8576 16664
rect 8330 16476 8576 16488
rect -98 16438 -52 16476
rect -98 16404 -92 16438
rect -58 16404 -52 16438
rect -98 16392 -52 16404
rect -98 16270 148 16282
rect -102 16094 -92 16270
rect -40 16094 -4 16270
rect 30 16094 108 16270
rect 142 16094 148 16270
rect -98 16082 148 16094
rect 4160 16270 4206 16476
rect 8530 16438 8576 16476
rect 8530 16404 8536 16438
rect 8570 16404 8576 16438
rect 8530 16392 8576 16404
rect 4272 16270 4318 16282
rect 8330 16270 8576 16282
rect 4160 16094 4166 16270
rect 4200 16094 4206 16270
rect 4253 16094 4263 16270
rect 4327 16094 4337 16270
rect 8330 16094 8336 16270
rect 8370 16094 8383 16270
rect 8435 16094 8448 16270
rect 8482 16094 8536 16270
rect 8570 16094 8576 16270
rect -98 16044 -52 16082
rect -98 16010 -92 16044
rect -58 16010 -52 16044
rect -98 15998 -52 16010
rect 108 16051 142 16082
rect 108 16050 1217 16051
rect 108 16044 3158 16050
rect 108 16010 1162 16044
rect 3146 16010 3158 16044
rect 108 16005 3158 16010
rect 1150 16004 3158 16005
rect 4160 15965 4206 16094
rect 4272 16082 4318 16094
rect 8330 16082 8576 16094
rect 8530 16044 8576 16082
rect 8530 16010 8536 16044
rect 8570 16010 8576 16044
rect 8530 15998 8576 16010
rect 8647 15965 8653 17581
rect -175 15959 8653 15965
rect 8687 17581 8699 17621
rect 8687 15965 8693 17581
rect 8687 15925 8699 15965
rect -221 15919 8699 15925
rect -215 15913 -169 15919
rect -1226 15869 -1180 15875
rect 856 15869 1662 15919
rect 4160 15913 4206 15919
rect 2588 15869 2634 15875
rect -1232 15863 2640 15869
rect -1232 15823 -1220 15863
rect -7901 15664 -7670 15685
rect -16711 15658 -7670 15664
rect -2996 15658 -2984 15698
rect -16705 15652 -16659 15658
rect -14377 15652 -14331 15658
rect -12319 15652 -12273 15658
rect -12489 15598 -12443 15604
rect -12144 15598 -11338 15658
rect -10261 15652 -10215 15658
rect -7949 15652 -2984 15658
rect -7949 15604 -7540 15652
rect -7966 15598 -7540 15604
rect -12495 15592 -7540 15598
rect -12495 15552 -12483 15592
rect -7926 15589 -7540 15592
rect -7926 15583 -7522 15589
rect -6595 15583 -5789 15652
rect -5356 15646 -5310 15652
rect -3036 15646 -2990 15652
rect -3076 15583 -3030 15589
rect -7926 15577 -3024 15583
rect -12489 14702 -12483 15552
rect -12495 14662 -12483 14702
rect -12449 15552 -7960 15558
rect -12449 14702 -12443 15552
rect -11736 15511 -11726 15514
rect -11738 15465 -11726 15511
rect -10742 15511 -10732 15514
rect -11736 15462 -11726 15465
rect -10742 15465 -10730 15511
rect -10742 15462 -10732 15465
rect -12374 15412 -12328 15424
rect -12374 15236 -12368 15412
rect -12334 15236 -12328 15412
rect -12374 15153 -12328 15236
rect -12286 15412 -12240 15424
rect -10234 15412 -10176 15552
rect -9678 15511 -9668 15514
rect -9680 15465 -9668 15511
rect -8684 15511 -8674 15514
rect -9678 15462 -9668 15465
rect -8684 15465 -8672 15511
rect -8684 15462 -8674 15465
rect -8170 15412 -8124 15424
rect -12286 15236 -12280 15412
rect -12246 15236 -12240 15412
rect -10241 15236 -10231 15412
rect -10179 15236 -10169 15412
rect -8170 15236 -8164 15412
rect -8130 15236 -8124 15412
rect -12387 15101 -12377 15153
rect -12325 15150 -12315 15153
rect -12286 15150 -12240 15236
rect -10228 15224 -10182 15236
rect -8170 15150 -8124 15236
rect -8082 15412 -8036 15424
rect -8082 15236 -8076 15412
rect -8042 15236 -8036 15412
rect -8082 15150 -8036 15236
rect -12325 15144 -8036 15150
rect -12325 15110 -8076 15144
rect -8042 15110 -8036 15144
rect -12325 15104 -8036 15110
rect -12325 15101 -12315 15104
rect -12374 15018 -12328 15101
rect -12374 14842 -12368 15018
rect -12334 14842 -12328 15018
rect -12374 14830 -12328 14842
rect -12286 15018 -12240 15104
rect -10228 15018 -10182 15030
rect -8170 15018 -8124 15104
rect -12286 14842 -12280 15018
rect -12246 14842 -12240 15018
rect -10241 14842 -10231 15018
rect -10179 14842 -10169 15018
rect -8170 14842 -8164 15018
rect -8130 14842 -8124 15018
rect -12286 14830 -12240 14842
rect -11738 14783 -10730 14789
rect -11738 14749 -11726 14783
rect -10742 14749 -10730 14783
rect -11738 14743 -10730 14749
rect -10234 14702 -10176 14842
rect -8170 14830 -8124 14842
rect -8082 15018 -8036 15104
rect -8082 14842 -8076 15018
rect -8042 14842 -8036 15018
rect -8082 14830 -8036 14842
rect -9680 14783 -8672 14789
rect -9680 14749 -9668 14783
rect -8684 14749 -8672 14783
rect -9680 14743 -8672 14749
rect -7966 14702 -7960 15552
rect -12449 14696 -7960 14702
rect -7926 15494 -7562 15577
rect -7926 14702 -7920 15494
rect -7926 14662 -7914 14702
rect -12495 14656 -7914 14662
rect -12489 14650 -12443 14656
rect -7966 14650 -7920 14656
rect -7847 14457 -7631 15494
rect -7568 14765 -7562 15494
rect -7574 14725 -7562 14765
rect -7528 15537 -3070 15543
rect -7528 14765 -7522 15537
rect -7468 15483 -7422 15489
rect -7380 15483 -7334 15489
rect -7468 15477 -7334 15483
rect -7472 15301 -7462 15477
rect -7410 15301 -7374 15477
rect -7340 15301 -7334 15477
rect -5322 15477 -5276 15489
rect -5322 15465 -5316 15477
rect -5282 15465 -5276 15477
rect -3264 15483 -3218 15489
rect -3176 15483 -3130 15489
rect -3264 15477 -3130 15483
rect -7468 15288 -7334 15301
rect -5335 15289 -5325 15465
rect -5273 15289 -5263 15465
rect -3264 15301 -3258 15477
rect -3224 15423 -3170 15477
rect -3136 15423 -3130 15477
rect -3224 15351 -3179 15423
rect -3127 15351 -3117 15423
rect -3224 15301 -3170 15351
rect -3136 15301 -3130 15351
rect -3264 15289 -3130 15301
rect -7468 15241 -7422 15288
rect -7468 15207 -7462 15241
rect -7428 15207 -7422 15241
rect -7468 15195 -7422 15207
rect -7380 15174 -7334 15288
rect -6832 15242 -3766 15248
rect -3264 15242 -3218 15289
rect -6832 15208 -6820 15242
rect -5836 15208 -4762 15242
rect -3778 15208 -3218 15242
rect -6832 15202 -3218 15208
rect -3176 15242 -3130 15289
rect -3176 15208 -3170 15242
rect -3136 15208 -3130 15242
rect -3796 15196 -3264 15202
rect -3176 15196 -3130 15208
rect -7380 15128 -4728 15174
rect -7468 15094 -7422 15106
rect -4774 15100 -4728 15128
rect -7468 15060 -7462 15094
rect -7428 15060 -7422 15094
rect -7468 15013 -7422 15060
rect -7380 15094 -5276 15100
rect -7380 15060 -6820 15094
rect -5836 15060 -5276 15094
rect -7380 15054 -5276 15060
rect -4774 15094 -3766 15100
rect -4774 15060 -4762 15094
rect -3778 15060 -3766 15094
rect -4774 15054 -3766 15060
rect -3176 15094 -3130 15106
rect -3176 15060 -3170 15094
rect -3136 15060 -3130 15094
rect -7380 15013 -7334 15054
rect -7468 15001 -7334 15013
rect -5322 15001 -5276 15054
rect -3176 15013 -3130 15060
rect -3264 15001 -3130 15013
rect -7468 14825 -7462 15001
rect -7428 14825 -7374 15001
rect -7340 14825 -7334 15001
rect -5335 14825 -5325 15001
rect -5273 14825 -5263 15001
rect -3264 14825 -3258 15001
rect -3224 14942 -3170 15001
rect -3136 14942 -3130 15001
rect -3224 14882 -3180 14942
rect -3128 14882 -3118 14942
rect -3224 14825 -3170 14882
rect -3136 14825 -3130 14882
rect -7468 14813 -7334 14825
rect -7380 14765 -7334 14813
rect -5322 14765 -5276 14825
rect -3264 14813 -3130 14825
rect -3076 14765 -3070 15537
rect -7528 14759 -3070 14765
rect -3036 15537 -3024 15577
rect -3036 14765 -3030 15537
rect -3036 14725 -3024 14765
rect -1226 14743 -1220 15823
rect -7574 14719 -3024 14725
rect -7568 14713 -7522 14719
rect -3076 14713 -3030 14719
rect -1232 14703 -1220 14743
rect -1186 15823 2594 15829
rect -1186 15723 -1180 15823
rect 2588 15723 2594 15823
rect -1186 15717 -653 15723
rect -1186 15679 -1062 15717
rect -665 15679 -653 15717
rect -1186 15673 -653 15679
rect 225 15717 1183 15723
rect 225 15679 237 15717
rect 634 15679 774 15717
rect 1171 15679 1183 15717
rect 225 15673 1183 15679
rect 2061 15717 2594 15723
rect 2061 15679 2073 15717
rect 2470 15679 2594 15717
rect 2061 15673 2594 15679
rect -1186 15391 -1180 15673
rect -1062 15558 -1010 15568
rect -1074 15507 -1062 15557
rect 774 15558 826 15568
rect -1010 15551 -653 15557
rect -665 15513 -653 15551
rect -1010 15507 -653 15513
rect 225 15551 729 15557
rect 225 15513 237 15551
rect 634 15513 729 15551
rect 225 15507 729 15513
rect 762 15507 774 15557
rect 2420 15558 2472 15568
rect 826 15551 1183 15557
rect 1171 15513 1183 15551
rect -1062 15496 -1010 15506
rect 582 15392 634 15402
rect -1186 15385 -653 15391
rect -1186 15347 -1062 15385
rect -665 15347 -653 15385
rect -1186 15341 -653 15347
rect 225 15385 582 15391
rect 679 15391 729 15507
rect 826 15507 1183 15513
rect 2061 15551 2420 15557
rect 2061 15513 2073 15551
rect 2061 15507 2420 15513
rect 774 15496 826 15506
rect 2472 15507 2482 15557
rect 2420 15496 2472 15506
rect 2063 15391 2073 15392
rect 225 15347 237 15385
rect 225 15341 582 15347
rect -1186 15225 -1102 15341
rect 634 15341 646 15391
rect 679 15385 1183 15391
rect 679 15347 774 15385
rect 1171 15347 1183 15385
rect 679 15341 1183 15347
rect 2061 15341 2073 15391
rect 2193 15391 2203 15392
rect 2193 15385 2560 15391
rect 2470 15347 2560 15385
rect 582 15330 634 15340
rect 582 15226 634 15236
rect -1186 15219 -653 15225
rect -1186 15181 -1062 15219
rect -665 15181 -653 15219
rect -1186 15175 -653 15181
rect 225 15219 582 15225
rect 679 15225 729 15341
rect 2063 15340 2073 15341
rect 2193 15341 2560 15347
rect 2193 15340 2203 15341
rect 2063 15225 2073 15226
rect 225 15181 237 15219
rect 225 15175 582 15181
rect -1186 14893 -1180 15175
rect 634 15175 646 15225
rect 679 15219 1183 15225
rect 679 15181 774 15219
rect 1171 15181 1183 15219
rect 679 15175 1183 15181
rect 2061 15175 2073 15225
rect 2193 15225 2203 15226
rect 2510 15225 2560 15341
rect 2193 15219 2560 15225
rect 2470 15181 2560 15219
rect 582 15164 634 15174
rect -1062 15060 -1010 15070
rect -1074 15009 -1062 15059
rect 679 15059 729 15175
rect 2063 15174 2073 15175
rect 2193 15175 2560 15181
rect 2193 15174 2203 15175
rect 764 15059 774 15060
rect -1010 15053 -653 15059
rect -665 15015 -653 15053
rect -1010 15009 -653 15015
rect 225 15053 729 15059
rect 225 15015 237 15053
rect 634 15015 729 15053
rect 225 15009 729 15015
rect 762 15009 774 15059
rect 826 15059 836 15060
rect 2408 15059 2418 15060
rect 826 15053 1183 15059
rect 1171 15015 1183 15053
rect 764 15008 774 15009
rect 826 15009 1183 15015
rect 2061 15053 2418 15059
rect 2470 15059 2480 15060
rect 2061 15015 2073 15053
rect 2061 15009 2418 15015
rect 826 15008 836 15009
rect 2408 15008 2418 15009
rect 2470 15009 2482 15059
rect 2470 15008 2480 15009
rect -1062 14998 -1010 15008
rect 2588 14893 2594 15673
rect -1186 14887 -653 14893
rect -1186 14849 -1062 14887
rect -665 14849 -653 14887
rect -1186 14843 -653 14849
rect 225 14887 1183 14893
rect 225 14849 237 14887
rect 634 14849 774 14887
rect 1171 14849 1183 14887
rect 225 14843 1183 14849
rect 2061 14887 2594 14893
rect 2061 14849 2073 14887
rect 2470 14849 2594 14887
rect 2061 14843 2594 14849
rect -1186 14743 -1180 14843
rect 2588 14743 2594 14843
rect -1186 14737 2594 14743
rect 2628 15823 2640 15863
rect 2628 14743 2634 15823
rect 2709 15821 4264 15885
rect 4328 15821 4338 15885
rect 2709 15310 2773 15821
rect 2859 15784 2905 15790
rect 4659 15784 5632 15919
rect 8647 15913 8693 15919
rect 8647 15784 8693 15790
rect 2853 15778 8699 15784
rect 2853 15738 2865 15778
rect 2709 15240 2773 15246
rect 2859 14826 2865 15738
rect 2853 14786 2865 14826
rect 2899 15738 8653 15744
rect 2899 14826 2905 15738
rect 2933 15664 8379 15710
rect 2933 14900 2979 15664
rect 3795 15624 3805 15627
rect 3793 15578 3805 15624
rect 5089 15624 5099 15627
rect 3795 15575 3805 15578
rect 5089 15578 5101 15624
rect 5089 15575 5099 15578
rect 3007 15534 3154 15546
rect 3007 15378 3013 15534
rect 3047 15378 3092 15534
rect 3144 15378 3154 15534
rect 3007 15366 3154 15378
rect 5753 15534 5799 15664
rect 8369 15650 8379 15664
rect 8439 15664 8619 15710
rect 8439 15650 8449 15664
rect 6453 15624 6463 15629
rect 6451 15578 6463 15624
rect 7747 15624 7757 15629
rect 6453 15573 6463 15578
rect 7747 15578 7759 15624
rect 7747 15573 7757 15578
rect 5753 15378 5759 15534
rect 5793 15378 5799 15534
rect 5753 15366 5799 15378
rect 8398 15534 8545 15546
rect 8398 15378 8408 15534
rect 8460 15378 8505 15534
rect 8539 15378 8545 15534
rect 8398 15366 8545 15378
rect 3007 15328 3053 15366
rect 6453 15334 6463 15337
rect 3007 15294 3013 15328
rect 3047 15294 3053 15328
rect 3007 15282 3053 15294
rect 3793 15328 5647 15334
rect 3793 15294 3805 15328
rect 5089 15294 5647 15328
rect 3793 15288 5647 15294
rect 6451 15288 6463 15334
rect 7747 15334 7757 15337
rect 5601 15263 5647 15288
rect 6453 15285 6463 15288
rect 7747 15288 7759 15334
rect 8499 15328 8545 15366
rect 8499 15294 8505 15328
rect 8539 15294 8545 15328
rect 7747 15285 7757 15288
rect 8499 15282 8545 15294
rect 5601 15217 5951 15263
rect 3007 15186 3053 15198
rect 3795 15192 3805 15195
rect 3007 15152 3013 15186
rect 3047 15152 3053 15186
rect 3007 15114 3053 15152
rect 3793 15146 3805 15192
rect 5089 15192 5099 15195
rect 5905 15192 5951 15217
rect 3795 15143 3805 15146
rect 5089 15146 5101 15192
rect 5905 15186 7759 15192
rect 5905 15152 6463 15186
rect 7747 15152 7759 15186
rect 5905 15146 7759 15152
rect 8499 15186 8545 15198
rect 8499 15152 8505 15186
rect 8539 15152 8545 15186
rect 5089 15143 5099 15146
rect 8499 15114 8545 15152
rect 3007 15102 3154 15114
rect 3007 14946 3013 15102
rect 3047 14946 3092 15102
rect 3144 14946 3154 15102
rect 3007 14934 3154 14946
rect 5753 15102 5799 15114
rect 5753 14946 5759 15102
rect 5793 14946 5799 15102
rect 5753 14900 5799 14946
rect 8398 15102 8545 15114
rect 8398 14946 8408 15102
rect 8460 14946 8505 15102
rect 8539 14946 8545 15102
rect 8398 14934 8545 14946
rect 8573 14900 8619 15664
rect 2933 14854 8619 14900
rect 8647 14826 8653 15738
rect 2899 14820 8653 14826
rect 8687 15738 8699 15778
rect 8687 14826 8693 15738
rect 8687 14786 8699 14826
rect 2853 14780 8699 14786
rect 2859 14774 2905 14780
rect 8647 14774 8693 14780
rect 2628 14703 2640 14743
rect -1232 14697 2640 14703
rect -1226 14691 -1180 14697
rect 2588 14691 2634 14697
rect -7847 14456 5584 14457
rect -7847 14240 5594 14456
rect 842 12250 1292 12256
rect 842 12216 854 12250
rect 1022 12216 1112 12250
rect 1280 12216 1292 12250
rect 842 12210 1292 12216
rect 1734 12250 2184 12256
rect 1734 12216 1746 12250
rect 1914 12216 2004 12250
rect 2172 12216 2184 12250
rect 1734 12210 2184 12216
rect 2626 12250 3076 12256
rect 2626 12216 2638 12250
rect 2806 12216 2896 12250
rect 3064 12216 3076 12250
rect 2626 12210 3076 12216
rect 3518 12250 3968 12256
rect 3518 12216 3530 12250
rect 3698 12216 3788 12250
rect 3956 12216 3968 12250
rect 3518 12210 3968 12216
rect 4332 12201 4617 12207
rect 698 12166 744 12178
rect 786 12166 832 12178
rect 1044 12166 1090 12178
rect 1302 12166 1348 12178
rect 698 11390 704 12166
rect 738 11390 744 12166
rect 773 11390 783 12166
rect 835 11390 845 12166
rect 1031 11390 1041 12166
rect 1093 11390 1103 12166
rect 1302 11390 1308 12166
rect 1342 11390 1348 12166
rect 698 11310 744 11390
rect 786 11310 832 11390
rect 1044 11378 1090 11390
rect 1302 11310 1348 11390
rect 1390 12166 1436 12178
rect 1390 11390 1396 12166
rect 1430 11390 1436 12166
rect 1390 11310 1436 11390
rect 698 11298 1436 11310
rect 698 11264 704 11298
rect 738 11264 1396 11298
rect 1430 11264 1436 11298
rect 698 11252 1436 11264
rect 698 11172 744 11252
rect 594 10471 647 10483
rect 594 10291 604 10471
rect 638 10291 647 10471
rect 698 10396 704 11172
rect 738 10396 744 11172
rect 698 10384 744 10396
rect 786 11172 832 11252
rect 1044 11172 1090 11184
rect 1302 11172 1348 11252
rect 786 10396 792 11172
rect 826 10396 832 11172
rect 1031 10396 1041 11172
rect 1093 10396 1103 11172
rect 1302 10396 1308 11172
rect 1342 10396 1348 11172
rect 786 10384 832 10396
rect 1044 10384 1090 10396
rect 1302 10384 1348 10396
rect 1390 11172 1436 11252
rect 1390 10396 1396 11172
rect 1430 10396 1436 11172
rect 1390 10384 1436 10396
rect 1590 12166 1636 12178
rect 1590 11390 1596 12166
rect 1630 11390 1636 12166
rect 1590 11317 1636 11390
rect 1678 12166 1724 12178
rect 1936 12166 1982 12178
rect 2194 12166 2240 12178
rect 1678 11390 1684 12166
rect 1718 11390 1724 12166
rect 1923 11390 1933 12166
rect 1985 11390 1995 12166
rect 2194 11390 2200 12166
rect 2234 11390 2240 12166
rect 1678 11317 1724 11390
rect 1936 11378 1982 11390
rect 1590 11310 1724 11317
rect 2194 11310 2240 11390
rect 2282 12166 2328 12178
rect 2282 11390 2288 12166
rect 2322 11390 2328 12166
rect 2282 11310 2328 11390
rect 1590 11307 2328 11310
rect 1590 11255 1596 11307
rect 1718 11298 2328 11307
rect 1718 11264 2288 11298
rect 2322 11264 2328 11298
rect 1718 11255 2328 11264
rect 1590 11252 2328 11255
rect 1590 11245 1724 11252
rect 1590 11172 1636 11245
rect 1590 10396 1596 11172
rect 1630 10396 1636 11172
rect 1590 10384 1636 10396
rect 1678 11172 1724 11245
rect 1936 11172 1982 11184
rect 2194 11172 2240 11252
rect 1678 10396 1684 11172
rect 1718 10396 1724 11172
rect 1923 10396 1933 11172
rect 1985 10396 1995 11172
rect 2194 10396 2200 11172
rect 2234 10396 2240 11172
rect 1678 10384 1724 10396
rect 1936 10384 1982 10396
rect 2194 10384 2240 10396
rect 2282 11172 2328 11252
rect 2282 10396 2288 11172
rect 2322 10396 2328 11172
rect 2282 10384 2328 10396
rect 2482 12166 2528 12178
rect 2482 11390 2488 12166
rect 2522 11390 2528 12166
rect 2482 11317 2528 11390
rect 2570 12166 2616 12178
rect 2828 12166 2874 12178
rect 3086 12166 3132 12178
rect 2570 11390 2576 12166
rect 2610 11390 2616 12166
rect 2815 11390 2825 12166
rect 2877 11390 2887 12166
rect 3086 11390 3092 12166
rect 3126 11390 3132 12166
rect 2570 11317 2616 11390
rect 2828 11378 2874 11390
rect 2482 11310 2616 11317
rect 3086 11310 3132 11390
rect 3174 12166 3220 12178
rect 3174 11390 3180 12166
rect 3214 11390 3220 12166
rect 3174 11310 3220 11390
rect 2482 11307 3220 11310
rect 2482 11255 2488 11307
rect 2610 11298 3220 11307
rect 2610 11264 3180 11298
rect 3214 11264 3220 11298
rect 2610 11255 3220 11264
rect 2482 11252 3220 11255
rect 2482 11245 2616 11252
rect 2482 11172 2528 11245
rect 2482 10396 2488 11172
rect 2522 10396 2528 11172
rect 2482 10384 2528 10396
rect 2570 11172 2616 11245
rect 2828 11172 2874 11184
rect 3086 11172 3132 11252
rect 2570 10396 2576 11172
rect 2610 10396 2616 11172
rect 2815 10396 2825 11172
rect 2877 10396 2887 11172
rect 3086 10396 3092 11172
rect 3126 10396 3132 11172
rect 2570 10384 2616 10396
rect 2828 10384 2874 10396
rect 3086 10384 3132 10396
rect 3174 11172 3220 11252
rect 3174 10396 3180 11172
rect 3214 10396 3220 11172
rect 3174 10384 3220 10396
rect 3374 12166 3420 12178
rect 3374 11390 3380 12166
rect 3414 11390 3420 12166
rect 3374 11317 3420 11390
rect 3462 12166 3508 12178
rect 3720 12166 3766 12178
rect 3978 12166 4024 12178
rect 3462 11390 3468 12166
rect 3502 11390 3508 12166
rect 3707 11390 3717 12166
rect 3769 11390 3779 12166
rect 3978 11390 3984 12166
rect 4018 11390 4024 12166
rect 3462 11317 3508 11390
rect 3720 11378 3766 11390
rect 3374 11310 3508 11317
rect 3978 11310 4024 11390
rect 4066 12166 4112 12178
rect 4066 11390 4072 12166
rect 4106 11390 4112 12166
rect 4332 12167 4344 12201
rect 4378 12167 4428 12201
rect 4604 12167 4617 12201
rect 4332 12161 4617 12167
rect 4334 12119 4380 12161
rect 4334 12113 4616 12119
rect 4334 12079 4428 12113
rect 4604 12079 4616 12113
rect 4334 12073 4616 12079
rect 4334 11603 4380 12073
rect 4648 12051 4694 12063
rect 4648 11883 4654 12051
rect 4688 11883 4694 12051
rect 4418 11861 4428 11864
rect 4416 11815 4428 11861
rect 4604 11861 4614 11864
rect 4418 11812 4428 11815
rect 4604 11815 4616 11861
rect 4604 11812 4614 11815
rect 4648 11793 4694 11883
rect 5378 11818 5594 14240
rect 4648 11625 4654 11793
rect 4688 11625 4694 11793
rect 4989 11812 5983 11818
rect 4989 11778 5001 11812
rect 5377 11778 5469 11812
rect 5503 11778 5595 11812
rect 5971 11778 5983 11812
rect 4989 11724 5983 11778
rect 4989 11690 5001 11724
rect 5377 11690 5595 11724
rect 5971 11690 5983 11724
rect 4989 11684 5983 11690
rect 4334 11597 4616 11603
rect 4334 11563 4428 11597
rect 4604 11563 4616 11597
rect 4334 11557 4616 11563
rect 4334 11515 4380 11557
rect 4418 11515 4428 11518
rect 4332 11509 4428 11515
rect 4604 11515 4614 11518
rect 4332 11475 4344 11509
rect 4378 11475 4428 11509
rect 4332 11469 4428 11475
rect 4418 11466 4428 11469
rect 4604 11469 4616 11515
rect 4604 11466 4614 11469
rect 4066 11310 4112 11390
rect 3374 11307 4112 11310
rect 4648 11307 4694 11625
rect 4902 11570 4948 11582
rect 4902 11386 4908 11570
rect 4942 11386 4948 11570
rect 3374 11255 3380 11307
rect 3502 11298 4112 11307
rect 3502 11264 4072 11298
rect 4106 11264 4112 11298
rect 3502 11255 4112 11264
rect 4635 11255 4645 11307
rect 4697 11255 4707 11307
rect 3374 11252 4112 11255
rect 3374 11245 3508 11252
rect 3374 11172 3420 11245
rect 3374 10396 3380 11172
rect 3414 10396 3420 11172
rect 3374 10384 3420 10396
rect 3462 11172 3508 11245
rect 3720 11172 3766 11184
rect 3978 11172 4024 11252
rect 3462 10396 3468 11172
rect 3502 10396 3508 11172
rect 3707 10396 3717 11172
rect 3769 10396 3779 11172
rect 3978 10396 3984 11172
rect 4018 10396 4024 11172
rect 3462 10384 3508 10396
rect 3720 10384 3766 10396
rect 3978 10384 4024 10396
rect 4066 11172 4112 11252
rect 4066 10396 4072 11172
rect 4106 10396 4112 11172
rect 4332 11087 4616 11093
rect 4332 11053 4344 11087
rect 4378 11053 4428 11087
rect 4604 11053 4616 11087
rect 4332 11047 4616 11053
rect 4334 11005 4380 11047
rect 4334 10999 4616 11005
rect 4334 10965 4428 10999
rect 4604 10965 4616 10999
rect 4334 10959 4616 10965
rect 4334 10489 4380 10959
rect 4648 10937 4694 11255
rect 4648 10769 4654 10937
rect 4688 10769 4694 10937
rect 4902 11112 4948 11386
rect 5001 11275 5377 11285
rect 4989 11226 5001 11272
rect 5377 11226 5389 11272
rect 5001 11213 5377 11223
rect 4902 10928 4908 11112
rect 4942 10928 4948 11112
rect 4902 10916 4948 10928
rect 5463 10814 5509 11684
rect 6024 11570 6070 11582
rect 6024 11386 6030 11570
rect 6064 11386 6070 11570
rect 6024 11374 6070 11386
rect 5595 11275 5971 11285
rect 5583 11226 5595 11272
rect 5971 11226 5983 11272
rect 5595 11213 5971 11223
rect 6024 11124 6069 11374
rect 6024 11112 6070 11124
rect 6024 10928 6030 11112
rect 6064 10966 6070 11112
rect 6064 10928 9119 10966
rect 6024 10917 9119 10928
rect 6024 10916 6070 10917
rect 4418 10747 4428 10750
rect 4416 10701 4428 10747
rect 4604 10747 4614 10750
rect 4418 10698 4428 10701
rect 4604 10701 4616 10747
rect 4604 10698 4614 10701
rect 4648 10679 4694 10769
rect 4989 10808 5983 10814
rect 4989 10774 5001 10808
rect 5377 10774 5595 10808
rect 5971 10774 5983 10808
rect 4989 10768 5983 10774
rect 5463 10726 5509 10768
rect 4989 10720 5983 10726
rect 4989 10686 5001 10720
rect 5377 10686 5469 10720
rect 5503 10686 5595 10720
rect 5971 10686 5983 10720
rect 4989 10680 5983 10686
rect 4648 10511 4654 10679
rect 4688 10511 4694 10679
rect 4648 10499 4694 10511
rect 4334 10483 4616 10489
rect 4334 10449 4428 10483
rect 4604 10449 4616 10483
rect 4334 10443 4616 10449
rect 4334 10401 4380 10443
rect 4418 10401 4428 10404
rect 4066 10384 4112 10396
rect 4332 10395 4428 10401
rect 4604 10401 4614 10404
rect 4332 10361 4344 10395
rect 4378 10361 4428 10395
rect 4332 10355 4428 10361
rect 4418 10352 4428 10355
rect 4604 10355 4617 10401
rect 4604 10352 4614 10355
rect 842 10346 1292 10352
rect 842 10312 854 10346
rect 1022 10312 1112 10346
rect 1280 10312 1292 10346
rect 842 10306 1292 10312
rect 1734 10346 2184 10352
rect 1734 10312 1746 10346
rect 1914 10312 2004 10346
rect 2172 10312 2184 10346
rect 1734 10306 2184 10312
rect 2626 10346 3076 10352
rect 2626 10312 2638 10346
rect 2806 10312 2896 10346
rect 3064 10312 3076 10346
rect 2626 10306 3076 10312
rect 3518 10346 3968 10352
rect 3518 10312 3530 10346
rect 3698 10312 3788 10346
rect 3956 10312 3968 10346
rect 3518 10306 3968 10312
rect 594 9818 647 10291
rect 745 10007 949 10013
rect 745 9973 757 10007
rect 937 9973 949 10007
rect 745 9967 949 9973
rect 1041 9979 1093 10306
rect 1933 10059 1985 10306
rect 2825 10139 2877 10306
rect 3717 10219 3769 10306
rect 3717 10167 9119 10219
rect 2825 10087 9119 10139
rect 1933 10007 9119 10059
rect 821 9899 874 9967
rect 1041 9927 9119 9979
rect 821 9846 9119 9899
rect 594 9765 9119 9818
rect 668 8022 6830 8067
rect 668 7988 713 8022
rect 747 7988 813 8022
rect 847 7988 913 8022
rect 947 7988 1013 8022
rect 1047 7988 1113 8022
rect 1147 7988 1213 8022
rect 1247 7988 2101 8022
rect 2135 7988 2201 8022
rect 2235 7988 2301 8022
rect 2335 7988 2401 8022
rect 2435 7988 2501 8022
rect 2535 7988 2601 8022
rect 2635 7988 3489 8022
rect 3523 7988 3589 8022
rect 3623 7988 3689 8022
rect 3723 7988 3789 8022
rect 3823 7988 3889 8022
rect 3923 7988 3989 8022
rect 4023 7988 4877 8022
rect 4911 7988 4977 8022
rect 5011 7988 5077 8022
rect 5111 7988 5177 8022
rect 5211 7988 5277 8022
rect 5311 7988 5377 8022
rect 5411 7988 6265 8022
rect 6299 7988 6365 8022
rect 6399 7988 6465 8022
rect 6499 7988 6565 8022
rect 6599 7988 6665 8022
rect 6699 7988 6765 8022
rect 6799 7988 6830 8022
rect 668 7922 6830 7988
rect 668 7888 713 7922
rect 747 7888 813 7922
rect 847 7888 913 7922
rect 947 7888 1013 7922
rect 1047 7888 1113 7922
rect 1147 7888 1213 7922
rect 1247 7911 2101 7922
rect 1247 7888 1278 7911
rect 668 7822 1278 7888
rect 668 7788 713 7822
rect 747 7788 813 7822
rect 847 7788 913 7822
rect 947 7788 1013 7822
rect 1047 7788 1113 7822
rect 1147 7788 1213 7822
rect 1247 7788 1278 7822
rect 668 7772 1278 7788
rect 667 7722 1278 7772
rect 667 7688 713 7722
rect 747 7688 813 7722
rect 847 7688 913 7722
rect 947 7688 1013 7722
rect 1047 7688 1113 7722
rect 1147 7688 1213 7722
rect 1247 7688 1278 7722
rect 667 7622 1278 7688
rect 667 7588 713 7622
rect 747 7588 813 7622
rect 847 7588 913 7622
rect 947 7588 1013 7622
rect 1047 7588 1113 7622
rect 1147 7588 1213 7622
rect 1247 7588 1278 7622
rect 667 7522 1278 7588
rect 667 7488 713 7522
rect 747 7488 813 7522
rect 847 7488 913 7522
rect 947 7488 1013 7522
rect 1047 7488 1113 7522
rect 1147 7488 1213 7522
rect 1247 7488 1278 7522
rect 667 7457 1278 7488
rect 667 7092 823 7457
rect 1643 7366 1691 7911
rect 2056 7888 2101 7911
rect 2135 7888 2201 7922
rect 2235 7888 2301 7922
rect 2335 7888 2401 7922
rect 2435 7888 2501 7922
rect 2535 7888 2601 7922
rect 2635 7911 3489 7922
rect 2635 7888 2666 7911
rect 2056 7822 2666 7888
rect 2056 7788 2101 7822
rect 2135 7788 2201 7822
rect 2235 7788 2301 7822
rect 2335 7788 2401 7822
rect 2435 7788 2501 7822
rect 2535 7788 2601 7822
rect 2635 7788 2666 7822
rect 2056 7722 2666 7788
rect 2056 7688 2101 7722
rect 2135 7688 2201 7722
rect 2235 7688 2301 7722
rect 2335 7688 2401 7722
rect 2435 7688 2501 7722
rect 2535 7688 2601 7722
rect 2635 7688 2666 7722
rect 2056 7622 2666 7688
rect 2056 7588 2101 7622
rect 2135 7588 2201 7622
rect 2235 7588 2301 7622
rect 2335 7588 2401 7622
rect 2435 7588 2501 7622
rect 2535 7588 2601 7622
rect 2635 7588 2666 7622
rect 2056 7522 2666 7588
rect 2056 7488 2101 7522
rect 2135 7488 2201 7522
rect 2235 7488 2301 7522
rect 2335 7488 2401 7522
rect 2435 7488 2501 7522
rect 2535 7488 2601 7522
rect 2635 7488 2666 7522
rect 2056 7457 2666 7488
rect 3031 7366 3079 7911
rect 3444 7888 3489 7911
rect 3523 7888 3589 7922
rect 3623 7888 3689 7922
rect 3723 7888 3789 7922
rect 3823 7888 3889 7922
rect 3923 7888 3989 7922
rect 4023 7911 4877 7922
rect 4023 7888 4054 7911
rect 3444 7822 4054 7888
rect 3444 7788 3489 7822
rect 3523 7788 3589 7822
rect 3623 7788 3689 7822
rect 3723 7788 3789 7822
rect 3823 7788 3889 7822
rect 3923 7788 3989 7822
rect 4023 7788 4054 7822
rect 3444 7722 4054 7788
rect 3444 7688 3489 7722
rect 3523 7688 3589 7722
rect 3623 7688 3689 7722
rect 3723 7688 3789 7722
rect 3823 7688 3889 7722
rect 3923 7688 3989 7722
rect 4023 7688 4054 7722
rect 3444 7622 4054 7688
rect 3444 7588 3489 7622
rect 3523 7588 3589 7622
rect 3623 7588 3689 7622
rect 3723 7588 3789 7622
rect 3823 7588 3889 7622
rect 3923 7588 3989 7622
rect 4023 7588 4054 7622
rect 3444 7522 4054 7588
rect 3444 7488 3489 7522
rect 3523 7488 3589 7522
rect 3623 7488 3689 7522
rect 3723 7488 3789 7522
rect 3823 7488 3889 7522
rect 3923 7488 3989 7522
rect 4023 7488 4054 7522
rect 3444 7457 4054 7488
rect 4419 7366 4467 7911
rect 4832 7888 4877 7911
rect 4911 7888 4977 7922
rect 5011 7888 5077 7922
rect 5111 7888 5177 7922
rect 5211 7888 5277 7922
rect 5311 7888 5377 7922
rect 5411 7911 6265 7922
rect 5411 7888 5442 7911
rect 4832 7822 5442 7888
rect 4832 7788 4877 7822
rect 4911 7788 4977 7822
rect 5011 7788 5077 7822
rect 5111 7788 5177 7822
rect 5211 7788 5277 7822
rect 5311 7788 5377 7822
rect 5411 7788 5442 7822
rect 4832 7722 5442 7788
rect 4832 7688 4877 7722
rect 4911 7688 4977 7722
rect 5011 7688 5077 7722
rect 5111 7688 5177 7722
rect 5211 7688 5277 7722
rect 5311 7688 5377 7722
rect 5411 7688 5442 7722
rect 4832 7622 5442 7688
rect 4832 7588 4877 7622
rect 4911 7588 4977 7622
rect 5011 7588 5077 7622
rect 5111 7588 5177 7622
rect 5211 7588 5277 7622
rect 5311 7588 5377 7622
rect 5411 7588 5442 7622
rect 4832 7522 5442 7588
rect 4832 7488 4877 7522
rect 4911 7488 4977 7522
rect 5011 7488 5077 7522
rect 5111 7488 5177 7522
rect 5211 7488 5277 7522
rect 5311 7488 5377 7522
rect 5411 7488 5442 7522
rect 4832 7457 5442 7488
rect 5807 7366 5855 7911
rect 6220 7888 6265 7911
rect 6299 7888 6365 7922
rect 6399 7888 6465 7922
rect 6499 7888 6565 7922
rect 6599 7888 6665 7922
rect 6699 7888 6765 7922
rect 6799 7888 6830 7922
rect 6220 7822 6830 7888
rect 6220 7788 6265 7822
rect 6299 7788 6365 7822
rect 6399 7788 6465 7822
rect 6499 7788 6565 7822
rect 6599 7788 6665 7822
rect 6699 7788 6765 7822
rect 6799 7788 6830 7822
rect 6220 7773 6830 7788
rect 6220 7722 6831 7773
rect 6220 7688 6265 7722
rect 6299 7688 6365 7722
rect 6399 7688 6465 7722
rect 6499 7688 6565 7722
rect 6599 7688 6665 7722
rect 6699 7688 6765 7722
rect 6799 7688 6831 7722
rect 6220 7622 6831 7688
rect 6220 7588 6265 7622
rect 6299 7588 6365 7622
rect 6399 7588 6465 7622
rect 6499 7588 6565 7622
rect 6599 7588 6665 7622
rect 6699 7588 6765 7622
rect 6799 7588 6831 7622
rect 6220 7522 6831 7588
rect 6220 7488 6265 7522
rect 6299 7488 6365 7522
rect 6399 7488 6465 7522
rect 6499 7488 6565 7522
rect 6599 7488 6665 7522
rect 6699 7488 6765 7522
rect 6799 7488 6831 7522
rect 6220 7457 6831 7488
rect 1369 7353 6128 7366
rect 1369 7281 1382 7353
rect 1454 7281 1518 7353
rect 1617 7281 2770 7353
rect 2842 7281 2906 7353
rect 3005 7281 3105 7353
rect 3204 7281 3268 7353
rect 3340 7281 4158 7353
rect 4230 7281 4294 7353
rect 4393 7281 4493 7353
rect 4592 7281 4656 7353
rect 4728 7281 5546 7353
rect 5618 7281 5682 7353
rect 5781 7281 5881 7353
rect 5980 7281 6044 7353
rect 6116 7281 6128 7353
rect 1369 7268 6128 7281
rect 1369 7217 1467 7268
rect 1369 7118 1382 7217
rect 1454 7118 1467 7217
rect 1369 7092 1467 7118
rect 667 7044 1467 7092
rect 667 6679 823 7044
rect 1369 7018 1467 7044
rect 1369 6919 1382 7018
rect 1454 6919 1467 7018
rect 1369 6855 1467 6919
rect 1369 6783 1382 6855
rect 1454 6783 1467 6855
rect 667 6634 1278 6679
rect 667 6600 713 6634
rect 747 6600 813 6634
rect 847 6600 913 6634
rect 947 6600 1013 6634
rect 1047 6600 1113 6634
rect 1147 6600 1213 6634
rect 1247 6600 1278 6634
rect 667 6534 1278 6600
rect 667 6500 713 6534
rect 747 6500 813 6534
rect 847 6500 913 6534
rect 947 6500 1013 6534
rect 1047 6500 1113 6534
rect 1147 6500 1213 6534
rect 1247 6500 1278 6534
rect 667 6434 1278 6500
rect 667 6400 713 6434
rect 747 6400 813 6434
rect 847 6400 913 6434
rect 947 6400 1013 6434
rect 1047 6400 1113 6434
rect 1147 6400 1213 6434
rect 1247 6400 1278 6434
rect 667 6334 1278 6400
rect 667 6300 713 6334
rect 747 6300 813 6334
rect 847 6300 913 6334
rect 947 6300 1013 6334
rect 1047 6300 1113 6334
rect 1147 6300 1213 6334
rect 1247 6300 1278 6334
rect 667 6234 1278 6300
rect 667 6200 713 6234
rect 747 6200 813 6234
rect 847 6200 913 6234
rect 947 6200 1013 6234
rect 1047 6200 1113 6234
rect 1147 6200 1213 6234
rect 1247 6200 1278 6234
rect 667 6134 1278 6200
rect 667 6100 713 6134
rect 747 6100 813 6134
rect 847 6100 913 6134
rect 947 6100 1013 6134
rect 1047 6100 1113 6134
rect 1147 6100 1213 6134
rect 1247 6100 1278 6134
rect 667 6069 1278 6100
rect 667 5704 823 6069
rect 1369 5965 1467 6783
rect 6030 7217 6128 7268
rect 6030 7118 6044 7217
rect 6116 7118 6128 7217
rect 6030 7092 6128 7118
rect 6675 7092 6831 7457
rect 6030 7044 6831 7092
rect 6030 7018 6128 7044
rect 6030 6919 6044 7018
rect 6116 6919 6128 7018
rect 6030 6855 6128 6919
rect 6030 6783 6044 6855
rect 6116 6783 6128 6855
rect 1369 5893 1382 5965
rect 1454 5893 1467 5965
rect 1369 5829 1467 5893
rect 1369 5730 1382 5829
rect 1454 5730 1467 5829
rect 1369 5706 1467 5730
rect 1369 5704 1415 5706
rect 667 5656 1415 5704
rect 667 5291 823 5656
rect 1369 5654 1415 5656
rect 1369 5630 1467 5654
rect 1369 5531 1382 5630
rect 1454 5531 1467 5630
rect 1369 5467 1467 5531
rect 1369 5395 1382 5467
rect 1454 5395 1467 5467
rect 667 5246 1278 5291
rect 667 5212 713 5246
rect 747 5212 813 5246
rect 847 5212 913 5246
rect 947 5212 1013 5246
rect 1047 5212 1113 5246
rect 1147 5212 1213 5246
rect 1247 5212 1278 5246
rect 667 5146 1278 5212
rect 667 5112 713 5146
rect 747 5112 813 5146
rect 847 5112 913 5146
rect 947 5112 1013 5146
rect 1047 5112 1113 5146
rect 1147 5112 1213 5146
rect 1247 5112 1278 5146
rect 667 5046 1278 5112
rect 667 5012 713 5046
rect 747 5012 813 5046
rect 847 5012 913 5046
rect 947 5012 1013 5046
rect 1047 5012 1113 5046
rect 1147 5012 1213 5046
rect 1247 5012 1278 5046
rect 667 4946 1278 5012
rect 667 4912 713 4946
rect 747 4912 813 4946
rect 847 4912 913 4946
rect 947 4912 1013 4946
rect 1047 4912 1113 4946
rect 1147 4912 1213 4946
rect 1247 4912 1278 4946
rect 667 4846 1278 4912
rect 667 4812 713 4846
rect 747 4812 813 4846
rect 847 4812 913 4846
rect 947 4812 1013 4846
rect 1047 4812 1113 4846
rect 1147 4812 1213 4846
rect 1247 4812 1278 4846
rect 667 4746 1278 4812
rect 667 4712 713 4746
rect 747 4712 813 4746
rect 847 4712 913 4746
rect 947 4712 1013 4746
rect 1047 4712 1113 4746
rect 1147 4712 1213 4746
rect 1247 4712 1278 4746
rect 667 4681 1278 4712
rect 667 4316 823 4681
rect 1369 4577 1467 5395
rect 1369 4505 1382 4577
rect 1454 4505 1467 4577
rect 1369 4441 1467 4505
rect 1369 4342 1382 4441
rect 1454 4342 1467 4441
rect 1369 4318 1467 4342
rect 1369 4316 1415 4318
rect 667 4268 1415 4316
rect 667 3903 823 4268
rect 1369 4266 1415 4268
rect 1369 4242 1467 4266
rect 1369 4143 1382 4242
rect 1454 4143 1467 4242
rect 1369 4079 1467 4143
rect 1369 4007 1382 4079
rect 1454 4007 1467 4079
rect 667 3858 1278 3903
rect 667 3824 713 3858
rect 747 3824 813 3858
rect 847 3824 913 3858
rect 947 3824 1013 3858
rect 1047 3824 1113 3858
rect 1147 3824 1213 3858
rect 1247 3824 1278 3858
rect 667 3758 1278 3824
rect 667 3724 713 3758
rect 747 3724 813 3758
rect 847 3724 913 3758
rect 947 3724 1013 3758
rect 1047 3724 1113 3758
rect 1147 3724 1213 3758
rect 1247 3724 1278 3758
rect 667 3658 1278 3724
rect 667 3624 713 3658
rect 747 3624 813 3658
rect 847 3624 913 3658
rect 947 3624 1013 3658
rect 1047 3624 1113 3658
rect 1147 3624 1213 3658
rect 1247 3624 1278 3658
rect 667 3558 1278 3624
rect 667 3524 713 3558
rect 747 3524 813 3558
rect 847 3524 913 3558
rect 947 3524 1013 3558
rect 1047 3524 1113 3558
rect 1147 3524 1213 3558
rect 1247 3524 1278 3558
rect 667 3458 1278 3524
rect 667 3424 713 3458
rect 747 3424 813 3458
rect 847 3424 913 3458
rect 947 3424 1013 3458
rect 1047 3424 1113 3458
rect 1147 3424 1213 3458
rect 1247 3424 1278 3458
rect 667 3358 1278 3424
rect 667 3324 713 3358
rect 747 3324 813 3358
rect 847 3324 913 3358
rect 947 3324 1013 3358
rect 1047 3324 1113 3358
rect 1147 3324 1213 3358
rect 1247 3324 1278 3358
rect 667 3293 1278 3324
rect 667 2928 823 3293
rect 1369 3189 1467 4007
rect 2056 6634 5442 6679
rect 2056 6600 2101 6634
rect 2135 6600 2201 6634
rect 2235 6600 2301 6634
rect 2335 6600 2401 6634
rect 2435 6600 2501 6634
rect 2535 6600 2601 6634
rect 2635 6600 3489 6634
rect 3523 6600 3589 6634
rect 3623 6600 3689 6634
rect 3723 6600 3789 6634
rect 3823 6600 3889 6634
rect 3923 6600 3989 6634
rect 4023 6600 4877 6634
rect 4911 6600 4977 6634
rect 5011 6600 5077 6634
rect 5111 6600 5177 6634
rect 5211 6600 5277 6634
rect 5311 6600 5377 6634
rect 5411 6600 5442 6634
rect 2056 6547 5442 6600
rect 2056 6534 2666 6547
rect 2056 6500 2101 6534
rect 2135 6500 2201 6534
rect 2235 6500 2301 6534
rect 2335 6500 2401 6534
rect 2435 6500 2501 6534
rect 2535 6500 2601 6534
rect 2635 6500 2666 6534
rect 2056 6434 2235 6500
rect 2501 6434 2666 6500
rect 2056 6400 2101 6434
rect 2135 6400 2201 6434
rect 2535 6400 2601 6434
rect 2635 6400 2666 6434
rect 2056 6334 2235 6400
rect 2501 6334 2666 6400
rect 2056 6300 2101 6334
rect 2135 6300 2201 6334
rect 2535 6300 2601 6334
rect 2635 6300 2666 6334
rect 2056 6234 2235 6300
rect 2501 6234 2666 6300
rect 2056 6200 2101 6234
rect 2135 6200 2201 6234
rect 2235 6200 2301 6234
rect 2335 6200 2401 6234
rect 2435 6200 2501 6234
rect 2535 6200 2601 6234
rect 2635 6200 2666 6234
rect 2056 6134 2666 6200
rect 2056 6100 2101 6134
rect 2135 6100 2201 6134
rect 2235 6100 2301 6134
rect 2335 6100 2401 6134
rect 2435 6100 2501 6134
rect 2535 6100 2601 6134
rect 2635 6100 2666 6134
rect 2056 6069 2666 6100
rect 3444 6534 4054 6547
rect 3444 6500 3489 6534
rect 3523 6500 3589 6534
rect 3623 6500 3689 6534
rect 3723 6500 3789 6534
rect 3823 6500 3889 6534
rect 3923 6500 3989 6534
rect 4023 6500 4054 6534
rect 3444 6434 4054 6500
rect 3444 6400 3489 6434
rect 3523 6400 3589 6434
rect 3623 6400 3689 6434
rect 3723 6400 3789 6434
rect 3823 6400 3889 6434
rect 3923 6400 3989 6434
rect 4023 6400 4054 6434
rect 3444 6334 4054 6400
rect 3444 6300 3489 6334
rect 3523 6300 3589 6334
rect 3623 6300 3689 6334
rect 3723 6300 3789 6334
rect 3823 6300 3889 6334
rect 3923 6300 3989 6334
rect 4023 6300 4054 6334
rect 3444 6234 4054 6300
rect 3444 6200 3489 6234
rect 3523 6200 3589 6234
rect 3623 6200 3689 6234
rect 3723 6200 3789 6234
rect 3823 6200 3889 6234
rect 3923 6200 3989 6234
rect 4023 6200 4054 6234
rect 3444 6134 4054 6200
rect 3444 6100 3489 6134
rect 3523 6100 3589 6134
rect 3623 6100 3689 6134
rect 3723 6100 3789 6134
rect 3823 6100 3889 6134
rect 3923 6100 3989 6134
rect 4023 6100 4054 6134
rect 3444 6069 4054 6100
rect 4832 6534 5442 6547
rect 4832 6500 4877 6534
rect 4911 6500 4977 6534
rect 5011 6500 5077 6534
rect 5111 6500 5177 6534
rect 5211 6500 5277 6534
rect 5311 6500 5377 6534
rect 5411 6500 5442 6534
rect 4832 6434 5442 6500
rect 4832 6400 4877 6434
rect 4911 6400 4977 6434
rect 5011 6400 5077 6434
rect 5111 6400 5177 6434
rect 5211 6400 5277 6434
rect 5311 6400 5377 6434
rect 5411 6400 5442 6434
rect 4832 6334 5442 6400
rect 4832 6300 4877 6334
rect 4911 6300 4977 6334
rect 5011 6300 5077 6334
rect 5111 6300 5177 6334
rect 5211 6300 5277 6334
rect 5311 6300 5377 6334
rect 5411 6300 5442 6334
rect 4832 6234 5442 6300
rect 4832 6200 4877 6234
rect 4911 6200 4977 6234
rect 5011 6200 5077 6234
rect 5111 6200 5177 6234
rect 5211 6200 5277 6234
rect 5311 6200 5377 6234
rect 5411 6200 5442 6234
rect 4832 6134 5442 6200
rect 4832 6100 4877 6134
rect 4911 6100 4977 6134
rect 5011 6100 5077 6134
rect 5111 6100 5177 6134
rect 5211 6100 5277 6134
rect 5311 6100 5377 6134
rect 5411 6100 5442 6134
rect 4832 6069 5442 6100
rect 2056 5291 2188 6069
rect 2758 5965 4740 5977
rect 2758 5893 2770 5965
rect 2842 5893 2906 5965
rect 3005 5893 3105 5965
rect 3204 5893 3268 5965
rect 3340 5893 4158 5965
rect 4230 5893 4294 5965
rect 4393 5893 4493 5965
rect 4592 5893 4656 5965
rect 4728 5893 4740 5965
rect 2758 5881 4740 5893
rect 2758 5829 2854 5881
rect 2758 5730 2770 5829
rect 2842 5730 2854 5829
rect 2758 5706 2854 5730
rect 2810 5654 2854 5706
rect 2758 5630 2854 5654
rect 2758 5531 2770 5630
rect 2842 5531 2854 5630
rect 2758 5467 2854 5531
rect 3262 5630 3346 5881
rect 3262 5531 3268 5630
rect 3340 5531 3346 5630
rect 3262 5473 3346 5531
rect 4152 5630 4236 5881
rect 4152 5531 4158 5630
rect 4230 5531 4236 5630
rect 4152 5473 4236 5531
rect 4644 5829 4740 5881
rect 4644 5730 4656 5829
rect 4728 5730 4740 5829
rect 4644 5706 4740 5730
rect 4644 5654 4688 5706
rect 4644 5630 4740 5654
rect 4644 5531 4656 5630
rect 4728 5531 4740 5630
rect 2758 5395 2770 5467
rect 2842 5395 2854 5467
rect 2056 5246 2666 5291
rect 2056 5212 2101 5246
rect 2135 5212 2201 5246
rect 2235 5212 2301 5246
rect 2335 5212 2401 5246
rect 2435 5212 2501 5246
rect 2535 5212 2601 5246
rect 2635 5212 2666 5246
rect 2056 5146 2666 5212
rect 2056 5112 2101 5146
rect 2135 5112 2201 5146
rect 2235 5112 2301 5146
rect 2335 5112 2401 5146
rect 2435 5112 2501 5146
rect 2535 5112 2601 5146
rect 2635 5112 2666 5146
rect 2056 5046 2666 5112
rect 2056 5012 2101 5046
rect 2135 5012 2201 5046
rect 2235 5012 2301 5046
rect 2335 5012 2401 5046
rect 2435 5012 2501 5046
rect 2535 5012 2601 5046
rect 2635 5012 2666 5046
rect 2056 4946 2666 5012
rect 2056 4912 2101 4946
rect 2135 4912 2201 4946
rect 2235 4912 2301 4946
rect 2335 4912 2401 4946
rect 2435 4912 2501 4946
rect 2535 4912 2601 4946
rect 2635 4912 2666 4946
rect 2056 4846 2666 4912
rect 2056 4812 2101 4846
rect 2135 4812 2201 4846
rect 2235 4812 2301 4846
rect 2335 4812 2401 4846
rect 2435 4812 2501 4846
rect 2535 4812 2601 4846
rect 2635 4812 2666 4846
rect 2056 4746 2666 4812
rect 2056 4712 2101 4746
rect 2135 4712 2201 4746
rect 2235 4712 2301 4746
rect 2335 4712 2401 4746
rect 2435 4712 2501 4746
rect 2535 4712 2601 4746
rect 2635 4712 2666 4746
rect 2056 4681 2666 4712
rect 2056 3903 2188 4681
rect 2758 4577 2854 5395
rect 3093 5467 4405 5473
rect 3093 5395 3105 5467
rect 3204 5395 3268 5467
rect 3340 5395 4158 5467
rect 4230 5395 4294 5467
rect 4393 5395 4405 5467
rect 3093 5389 4405 5395
rect 4644 5467 4740 5531
rect 4644 5395 4656 5467
rect 4728 5395 4740 5467
rect 3262 4583 3346 5389
rect 3444 5246 4054 5291
rect 3444 5212 3489 5246
rect 3523 5212 3589 5246
rect 3623 5212 3689 5246
rect 3723 5212 3789 5246
rect 3823 5212 3889 5246
rect 3923 5212 3989 5246
rect 4023 5212 4054 5246
rect 3444 5146 4054 5212
rect 3444 5112 3489 5146
rect 3523 5112 3589 5146
rect 3623 5112 3689 5146
rect 3723 5118 3789 5146
rect 3823 5112 3889 5146
rect 3923 5112 3989 5146
rect 4023 5112 4054 5146
rect 3444 5046 3689 5112
rect 3793 5046 4054 5112
rect 3444 5012 3489 5046
rect 3523 5012 3589 5046
rect 3623 5012 3689 5046
rect 3823 5012 3889 5046
rect 3923 5012 3989 5046
rect 4023 5012 4054 5046
rect 3444 4946 3689 5012
rect 3793 4946 4054 5012
rect 3444 4912 3489 4946
rect 3523 4912 3589 4946
rect 3623 4912 3689 4946
rect 3823 4912 3889 4946
rect 3923 4912 3989 4946
rect 4023 4912 4054 4946
rect 3444 4870 3689 4912
rect 3793 4870 4054 4912
rect 3444 4846 4054 4870
rect 3444 4812 3489 4846
rect 3523 4812 3589 4846
rect 3623 4812 3689 4846
rect 3723 4812 3789 4846
rect 3823 4812 3889 4846
rect 3923 4812 3989 4846
rect 4023 4812 4054 4846
rect 3444 4746 4054 4812
rect 3444 4712 3489 4746
rect 3523 4712 3589 4746
rect 3623 4712 3689 4746
rect 3723 4712 3789 4746
rect 3823 4712 3889 4746
rect 3923 4712 3989 4746
rect 4023 4712 4054 4746
rect 3444 4681 4054 4712
rect 4152 4583 4236 5389
rect 2758 4505 2770 4577
rect 2842 4505 2854 4577
rect 2758 4441 2854 4505
rect 3093 4577 4405 4583
rect 3093 4505 3105 4577
rect 3204 4505 3268 4577
rect 3340 4505 4158 4577
rect 4230 4505 4294 4577
rect 4393 4505 4405 4577
rect 3093 4499 4405 4505
rect 4644 4577 4740 5395
rect 5310 5291 5442 6069
rect 4832 5246 5442 5291
rect 4832 5212 4877 5246
rect 4911 5212 4977 5246
rect 5011 5212 5077 5246
rect 5111 5212 5177 5246
rect 5211 5212 5277 5246
rect 5311 5212 5377 5246
rect 5411 5212 5442 5246
rect 4832 5146 5442 5212
rect 4832 5112 4877 5146
rect 4911 5112 4977 5146
rect 5011 5112 5077 5146
rect 5111 5112 5177 5146
rect 5211 5112 5277 5146
rect 5311 5112 5377 5146
rect 5411 5112 5442 5146
rect 4832 5046 5442 5112
rect 4832 5012 4877 5046
rect 4911 5012 4977 5046
rect 5011 5012 5077 5046
rect 5111 5012 5177 5046
rect 5211 5012 5277 5046
rect 5311 5012 5377 5046
rect 5411 5012 5442 5046
rect 4832 4946 5442 5012
rect 4832 4912 4877 4946
rect 4911 4912 4977 4946
rect 5011 4912 5077 4946
rect 5111 4912 5177 4946
rect 5211 4912 5277 4946
rect 5311 4912 5377 4946
rect 5411 4912 5442 4946
rect 4832 4846 5442 4912
rect 4832 4812 4877 4846
rect 4911 4812 4977 4846
rect 5011 4812 5077 4846
rect 5111 4812 5177 4846
rect 5211 4812 5277 4846
rect 5311 4812 5377 4846
rect 5411 4812 5442 4846
rect 4832 4746 5442 4812
rect 4832 4712 4877 4746
rect 4911 4712 4977 4746
rect 5011 4712 5077 4746
rect 5111 4712 5177 4746
rect 5211 4712 5277 4746
rect 5311 4712 5377 4746
rect 5411 4712 5442 4746
rect 4832 4681 5442 4712
rect 4644 4505 4656 4577
rect 4728 4505 4740 4577
rect 2758 4342 2770 4441
rect 2842 4342 2854 4441
rect 2758 4318 2854 4342
rect 3262 4441 3346 4499
rect 3262 4342 3268 4441
rect 3340 4435 3346 4441
rect 4152 4441 4236 4499
rect 3340 4342 3347 4435
rect 3262 4330 3347 4342
rect 2810 4266 2854 4318
rect 2758 4242 2854 4266
rect 2758 4143 2770 4242
rect 2842 4143 2854 4242
rect 2758 4091 2854 4143
rect 3263 4091 3347 4330
rect 4152 4342 4158 4441
rect 4230 4342 4236 4441
rect 4152 4091 4236 4342
rect 4644 4441 4740 4505
rect 4644 4342 4656 4441
rect 4728 4342 4740 4441
rect 4644 4318 4740 4342
rect 4644 4266 4688 4318
rect 4644 4242 4740 4266
rect 4644 4143 4656 4242
rect 4728 4143 4740 4242
rect 4644 4091 4740 4143
rect 2758 4079 4740 4091
rect 2758 4007 2770 4079
rect 2842 4007 2906 4079
rect 3005 4007 3105 4079
rect 3204 4007 3268 4079
rect 3340 4007 4158 4079
rect 4230 4007 4294 4079
rect 4393 4007 4493 4079
rect 4592 4007 4656 4079
rect 4728 4007 4740 4079
rect 2758 3995 4740 4007
rect 5310 3903 5442 4681
rect 2056 3858 2666 3903
rect 2056 3824 2101 3858
rect 2135 3824 2201 3858
rect 2235 3824 2301 3858
rect 2335 3824 2401 3858
rect 2435 3824 2501 3858
rect 2535 3824 2601 3858
rect 2635 3824 2666 3858
rect 2056 3758 2666 3824
rect 2056 3724 2101 3758
rect 2135 3724 2201 3758
rect 2235 3724 2301 3758
rect 2335 3724 2401 3758
rect 2435 3724 2501 3758
rect 2535 3724 2601 3758
rect 2635 3724 2666 3758
rect 2056 3658 2666 3724
rect 2056 3624 2101 3658
rect 2135 3624 2201 3658
rect 2235 3624 2301 3658
rect 2335 3624 2401 3658
rect 2435 3624 2501 3658
rect 2535 3624 2601 3658
rect 2635 3624 2666 3658
rect 2056 3558 2666 3624
rect 2056 3524 2101 3558
rect 2135 3524 2201 3558
rect 2235 3524 2301 3558
rect 2335 3524 2401 3558
rect 2435 3524 2501 3558
rect 2535 3524 2601 3558
rect 2635 3524 2666 3558
rect 2056 3458 2666 3524
rect 2056 3424 2101 3458
rect 2135 3424 2201 3458
rect 2235 3424 2301 3458
rect 2335 3424 2401 3458
rect 2435 3424 2501 3458
rect 2535 3424 2601 3458
rect 2635 3425 2666 3458
rect 3444 3858 4054 3903
rect 3444 3824 3489 3858
rect 3523 3824 3589 3858
rect 3623 3824 3689 3858
rect 3723 3824 3789 3858
rect 3823 3824 3889 3858
rect 3923 3824 3989 3858
rect 4023 3824 4054 3858
rect 3444 3758 4054 3824
rect 3444 3724 3489 3758
rect 3523 3724 3589 3758
rect 3623 3724 3689 3758
rect 3723 3724 3789 3758
rect 3823 3724 3889 3758
rect 3923 3724 3989 3758
rect 4023 3724 4054 3758
rect 3444 3658 4054 3724
rect 3444 3624 3489 3658
rect 3523 3624 3589 3658
rect 3623 3624 3689 3658
rect 3723 3624 3789 3658
rect 3823 3624 3889 3658
rect 3923 3624 3989 3658
rect 4023 3624 4054 3658
rect 3444 3558 4054 3624
rect 3444 3524 3489 3558
rect 3523 3524 3589 3558
rect 3623 3524 3689 3558
rect 3723 3524 3789 3558
rect 3823 3524 3889 3558
rect 3923 3524 3989 3558
rect 4023 3524 4054 3558
rect 3444 3458 4054 3524
rect 3444 3425 3489 3458
rect 2635 3424 3489 3425
rect 3523 3424 3589 3458
rect 3623 3424 3689 3458
rect 3723 3424 3789 3458
rect 3823 3424 3889 3458
rect 3923 3424 3989 3458
rect 4023 3425 4054 3458
rect 4832 3858 5442 3903
rect 4832 3824 4877 3858
rect 4911 3824 4977 3858
rect 5011 3824 5077 3858
rect 5111 3824 5177 3858
rect 5211 3824 5277 3858
rect 5311 3824 5377 3858
rect 5411 3824 5442 3858
rect 4832 3758 5442 3824
rect 4832 3724 4877 3758
rect 4911 3724 4977 3758
rect 5011 3724 5077 3758
rect 5111 3724 5177 3758
rect 5211 3724 5277 3758
rect 5311 3724 5377 3758
rect 5411 3724 5442 3758
rect 4832 3658 5442 3724
rect 4832 3624 4877 3658
rect 4911 3624 4977 3658
rect 5011 3624 5077 3658
rect 5111 3624 5177 3658
rect 5211 3624 5277 3658
rect 5311 3624 5377 3658
rect 5411 3624 5442 3658
rect 4832 3558 5442 3624
rect 4832 3524 4877 3558
rect 4911 3524 4977 3558
rect 5011 3524 5077 3558
rect 5111 3524 5177 3558
rect 5211 3524 5277 3558
rect 5311 3524 5377 3558
rect 5411 3524 5442 3558
rect 4832 3458 5442 3524
rect 4832 3425 4877 3458
rect 4023 3424 4877 3425
rect 4911 3424 4977 3458
rect 5011 3424 5077 3458
rect 5111 3424 5177 3458
rect 5211 3424 5277 3458
rect 5311 3424 5377 3458
rect 5411 3424 5442 3458
rect 2056 3358 5442 3424
rect 2056 3324 2101 3358
rect 2135 3324 2201 3358
rect 2235 3324 2301 3358
rect 2335 3324 2401 3358
rect 2435 3324 2501 3358
rect 2535 3324 2601 3358
rect 2635 3324 3489 3358
rect 3523 3324 3589 3358
rect 3623 3324 3689 3358
rect 3723 3324 3789 3358
rect 3823 3324 3889 3358
rect 3923 3324 3989 3358
rect 4023 3324 4877 3358
rect 4911 3324 4977 3358
rect 5011 3324 5077 3358
rect 5111 3324 5177 3358
rect 5211 3324 5277 3358
rect 5311 3324 5377 3358
rect 5411 3324 5442 3358
rect 2056 3293 5442 3324
rect 6030 5965 6128 6783
rect 6675 6679 6831 7044
rect 6220 6634 6831 6679
rect 6220 6600 6265 6634
rect 6299 6600 6365 6634
rect 6399 6600 6465 6634
rect 6499 6600 6565 6634
rect 6599 6600 6665 6634
rect 6699 6600 6765 6634
rect 6799 6600 6831 6634
rect 6220 6534 6831 6600
rect 6220 6500 6265 6534
rect 6299 6500 6365 6534
rect 6399 6500 6465 6534
rect 6499 6500 6565 6534
rect 6599 6500 6665 6534
rect 6699 6500 6765 6534
rect 6799 6500 6831 6534
rect 6220 6434 6831 6500
rect 6220 6400 6265 6434
rect 6299 6400 6365 6434
rect 6399 6400 6465 6434
rect 6499 6400 6565 6434
rect 6599 6400 6665 6434
rect 6699 6400 6765 6434
rect 6799 6400 6831 6434
rect 6220 6334 6831 6400
rect 6220 6300 6265 6334
rect 6299 6300 6365 6334
rect 6399 6300 6465 6334
rect 6499 6300 6565 6334
rect 6599 6300 6665 6334
rect 6699 6300 6765 6334
rect 6799 6300 6831 6334
rect 6220 6234 6831 6300
rect 6220 6200 6265 6234
rect 6299 6200 6365 6234
rect 6399 6200 6465 6234
rect 6499 6200 6565 6234
rect 6599 6200 6665 6234
rect 6699 6200 6765 6234
rect 6799 6200 6831 6234
rect 6220 6134 6831 6200
rect 6220 6100 6265 6134
rect 6299 6100 6365 6134
rect 6399 6100 6465 6134
rect 6499 6100 6565 6134
rect 6599 6100 6665 6134
rect 6699 6100 6765 6134
rect 6799 6100 6831 6134
rect 6220 6069 6831 6100
rect 6030 5893 6044 5965
rect 6116 5893 6128 5965
rect 6030 5829 6128 5893
rect 6030 5730 6044 5829
rect 6116 5730 6128 5829
rect 6030 5706 6128 5730
rect 6082 5704 6128 5706
rect 6675 5704 6831 6069
rect 6082 5656 6831 5704
rect 6082 5654 6128 5656
rect 6030 5630 6128 5654
rect 6030 5531 6044 5630
rect 6116 5531 6128 5630
rect 6030 5467 6128 5531
rect 6030 5395 6044 5467
rect 6116 5395 6128 5467
rect 6030 4577 6128 5395
rect 6675 5291 6831 5656
rect 6220 5246 6831 5291
rect 6220 5212 6265 5246
rect 6299 5212 6365 5246
rect 6399 5212 6465 5246
rect 6499 5212 6565 5246
rect 6599 5212 6665 5246
rect 6699 5212 6765 5246
rect 6799 5212 6831 5246
rect 6220 5146 6831 5212
rect 6220 5112 6265 5146
rect 6299 5112 6365 5146
rect 6399 5112 6465 5146
rect 6499 5112 6565 5146
rect 6599 5112 6665 5146
rect 6699 5112 6765 5146
rect 6799 5112 6831 5146
rect 6220 5046 6831 5112
rect 6220 5012 6265 5046
rect 6299 5012 6365 5046
rect 6399 5012 6465 5046
rect 6499 5012 6565 5046
rect 6599 5012 6665 5046
rect 6699 5012 6765 5046
rect 6799 5012 6831 5046
rect 6220 4946 6831 5012
rect 6220 4912 6265 4946
rect 6299 4912 6365 4946
rect 6399 4912 6465 4946
rect 6499 4912 6565 4946
rect 6599 4912 6665 4946
rect 6699 4912 6765 4946
rect 6799 4912 6831 4946
rect 6220 4846 6831 4912
rect 6220 4812 6265 4846
rect 6299 4812 6365 4846
rect 6399 4812 6465 4846
rect 6499 4812 6565 4846
rect 6599 4812 6665 4846
rect 6699 4812 6765 4846
rect 6799 4812 6831 4846
rect 6220 4746 6831 4812
rect 6220 4712 6265 4746
rect 6299 4712 6365 4746
rect 6399 4712 6465 4746
rect 6499 4712 6565 4746
rect 6599 4712 6665 4746
rect 6699 4712 6765 4746
rect 6799 4712 6831 4746
rect 6220 4681 6831 4712
rect 6030 4505 6044 4577
rect 6116 4505 6128 4577
rect 6030 4441 6128 4505
rect 6030 4342 6044 4441
rect 6116 4342 6128 4441
rect 6030 4318 6128 4342
rect 6082 4316 6128 4318
rect 6675 4316 6831 4681
rect 6082 4268 6831 4316
rect 6082 4266 6128 4268
rect 6030 4242 6128 4266
rect 6030 4143 6044 4242
rect 6116 4143 6128 4242
rect 6030 4079 6128 4143
rect 6030 4007 6044 4079
rect 6116 4007 6128 4079
rect 1369 3117 1382 3189
rect 1454 3117 1467 3189
rect 1369 3053 1467 3117
rect 1369 2954 1382 3053
rect 1454 2954 1467 3053
rect 1369 2928 1467 2954
rect 667 2880 1467 2928
rect 667 2515 823 2880
rect 1369 2854 1467 2880
rect 1369 2755 1382 2854
rect 1454 2755 1467 2854
rect 1369 2704 1467 2755
rect 6030 3189 6128 4007
rect 6675 3903 6831 4268
rect 6220 3858 6831 3903
rect 6220 3824 6265 3858
rect 6299 3824 6365 3858
rect 6399 3824 6465 3858
rect 6499 3824 6565 3858
rect 6599 3824 6665 3858
rect 6699 3824 6765 3858
rect 6799 3824 6831 3858
rect 6220 3758 6831 3824
rect 6220 3724 6265 3758
rect 6299 3724 6365 3758
rect 6399 3724 6465 3758
rect 6499 3724 6565 3758
rect 6599 3724 6665 3758
rect 6699 3724 6765 3758
rect 6799 3724 6831 3758
rect 6220 3658 6831 3724
rect 6220 3624 6265 3658
rect 6299 3624 6365 3658
rect 6399 3624 6465 3658
rect 6499 3624 6565 3658
rect 6599 3624 6665 3658
rect 6699 3624 6765 3658
rect 6799 3624 6831 3658
rect 6220 3558 6831 3624
rect 6220 3524 6265 3558
rect 6299 3524 6365 3558
rect 6399 3524 6465 3558
rect 6499 3524 6565 3558
rect 6599 3524 6665 3558
rect 6699 3524 6765 3558
rect 6799 3524 6831 3558
rect 6220 3458 6831 3524
rect 6220 3424 6265 3458
rect 6299 3424 6365 3458
rect 6399 3424 6465 3458
rect 6499 3424 6565 3458
rect 6599 3424 6665 3458
rect 6699 3424 6765 3458
rect 6799 3424 6831 3458
rect 6220 3358 6831 3424
rect 6220 3324 6265 3358
rect 6299 3324 6365 3358
rect 6399 3324 6465 3358
rect 6499 3324 6565 3358
rect 6599 3324 6665 3358
rect 6699 3324 6765 3358
rect 6799 3324 6831 3358
rect 6220 3293 6831 3324
rect 6030 3117 6044 3189
rect 6116 3117 6128 3189
rect 6030 3053 6128 3117
rect 6030 2954 6044 3053
rect 6116 2954 6128 3053
rect 6030 2928 6128 2954
rect 6675 2928 6831 3293
rect 6030 2880 6831 2928
rect 6030 2854 6128 2880
rect 6030 2755 6043 2854
rect 6115 2755 6128 2854
rect 6030 2704 6128 2755
rect 1369 2691 6128 2704
rect 1369 2619 1382 2691
rect 1454 2619 1518 2691
rect 1617 2619 1717 2691
rect 1816 2619 1880 2691
rect 1952 2619 2770 2691
rect 2842 2619 2906 2691
rect 3005 2619 3105 2691
rect 3204 2619 3268 2691
rect 3340 2619 4158 2691
rect 4230 2619 4294 2691
rect 4393 2619 4493 2691
rect 4592 2619 4656 2691
rect 4728 2619 5546 2691
rect 5618 2619 5682 2691
rect 5781 2619 5880 2691
rect 5979 2619 6043 2691
rect 6115 2619 6128 2691
rect 1369 2606 6128 2619
rect 658 1904 668 2515
rect 1278 2060 1288 2515
rect 1643 2060 1691 2606
rect 2056 2470 2666 2515
rect 2056 2436 2101 2470
rect 2135 2436 2201 2470
rect 2235 2436 2301 2470
rect 2335 2436 2401 2470
rect 2435 2436 2501 2470
rect 2535 2436 2601 2470
rect 2635 2436 2666 2470
rect 2056 2370 2666 2436
rect 2056 2336 2101 2370
rect 2135 2336 2201 2370
rect 2235 2336 2301 2370
rect 2335 2336 2401 2370
rect 2435 2336 2501 2370
rect 2535 2336 2601 2370
rect 2635 2336 2666 2370
rect 2056 2270 2666 2336
rect 2056 2236 2101 2270
rect 2135 2236 2201 2270
rect 2235 2236 2301 2270
rect 2335 2236 2401 2270
rect 2435 2236 2501 2270
rect 2535 2236 2601 2270
rect 2635 2236 2666 2270
rect 2056 2170 2666 2236
rect 2056 2136 2101 2170
rect 2135 2136 2201 2170
rect 2235 2136 2301 2170
rect 2335 2136 2401 2170
rect 2435 2136 2501 2170
rect 2535 2136 2601 2170
rect 2635 2136 2666 2170
rect 2056 2070 2666 2136
rect 2056 2060 2101 2070
rect 1278 2036 2101 2060
rect 2135 2036 2201 2070
rect 2235 2036 2301 2070
rect 2335 2036 2401 2070
rect 2435 2036 2501 2070
rect 2535 2036 2601 2070
rect 2635 2060 2666 2070
rect 3031 2060 3079 2606
rect 3444 2470 4054 2515
rect 3444 2436 3489 2470
rect 3523 2436 3589 2470
rect 3623 2436 3689 2470
rect 3723 2436 3789 2470
rect 3823 2436 3889 2470
rect 3923 2436 3989 2470
rect 4023 2436 4054 2470
rect 3444 2370 4054 2436
rect 3444 2336 3489 2370
rect 3523 2336 3589 2370
rect 3623 2336 3689 2370
rect 3723 2336 3789 2370
rect 3823 2336 3889 2370
rect 3923 2336 3989 2370
rect 4023 2336 4054 2370
rect 3444 2270 4054 2336
rect 3444 2236 3489 2270
rect 3523 2236 3589 2270
rect 3623 2236 3689 2270
rect 3723 2236 3789 2270
rect 3823 2236 3889 2270
rect 3923 2236 3989 2270
rect 4023 2236 4054 2270
rect 3444 2170 4054 2236
rect 3444 2136 3489 2170
rect 3523 2136 3589 2170
rect 3623 2136 3689 2170
rect 3723 2136 3789 2170
rect 3823 2136 3889 2170
rect 3923 2136 3989 2170
rect 4023 2136 4054 2170
rect 3444 2070 4054 2136
rect 3444 2060 3489 2070
rect 2635 2036 3489 2060
rect 3523 2036 3589 2070
rect 3623 2036 3689 2070
rect 3723 2036 3789 2070
rect 3823 2036 3889 2070
rect 3923 2036 3989 2070
rect 4023 2060 4054 2070
rect 4419 2060 4467 2606
rect 4832 2470 5442 2515
rect 4832 2436 4877 2470
rect 4911 2436 4977 2470
rect 5011 2436 5077 2470
rect 5111 2436 5177 2470
rect 5211 2436 5277 2470
rect 5311 2436 5377 2470
rect 5411 2436 5442 2470
rect 4832 2370 5442 2436
rect 4832 2336 4877 2370
rect 4911 2336 4977 2370
rect 5011 2336 5077 2370
rect 5111 2336 5177 2370
rect 5211 2336 5277 2370
rect 5311 2336 5377 2370
rect 5411 2336 5442 2370
rect 4832 2270 5442 2336
rect 4832 2236 4877 2270
rect 4911 2236 4977 2270
rect 5011 2236 5077 2270
rect 5111 2236 5177 2270
rect 5211 2236 5277 2270
rect 5311 2236 5377 2270
rect 5411 2236 5442 2270
rect 4832 2170 5442 2236
rect 4832 2136 4877 2170
rect 4911 2136 4977 2170
rect 5011 2136 5077 2170
rect 5111 2136 5177 2170
rect 5211 2136 5277 2170
rect 5311 2136 5377 2170
rect 5411 2136 5442 2170
rect 4832 2070 5442 2136
rect 4832 2060 4877 2070
rect 4023 2036 4877 2060
rect 4911 2036 4977 2070
rect 5011 2036 5077 2070
rect 5111 2036 5177 2070
rect 5211 2036 5277 2070
rect 5311 2036 5377 2070
rect 5411 2060 5442 2070
rect 5807 2060 5855 2606
rect 6675 2515 6831 2880
rect 6220 2470 6831 2515
rect 6220 2436 6265 2470
rect 6299 2436 6365 2470
rect 6399 2436 6465 2470
rect 6499 2436 6565 2470
rect 6599 2436 6665 2470
rect 6699 2436 6765 2470
rect 6799 2436 6831 2470
rect 6220 2417 6831 2436
rect 6220 2370 6830 2417
rect 6220 2336 6265 2370
rect 6299 2336 6365 2370
rect 6399 2336 6465 2370
rect 6499 2336 6565 2370
rect 6599 2336 6665 2370
rect 6699 2336 6765 2370
rect 6799 2336 6830 2370
rect 6220 2270 6830 2336
rect 6220 2236 6265 2270
rect 6299 2236 6365 2270
rect 6399 2236 6465 2270
rect 6499 2236 6565 2270
rect 6599 2236 6665 2270
rect 6699 2236 6765 2270
rect 6799 2236 6830 2270
rect 6220 2170 6830 2236
rect 6220 2136 6265 2170
rect 6299 2136 6365 2170
rect 6399 2136 6465 2170
rect 6499 2136 6565 2170
rect 6599 2136 6665 2170
rect 6699 2136 6765 2170
rect 6799 2136 6830 2170
rect 6220 2070 6830 2136
rect 6220 2060 6265 2070
rect 5411 2036 6265 2060
rect 6299 2036 6365 2070
rect 6399 2036 6465 2070
rect 6499 2036 6565 2070
rect 6599 2036 6665 2070
rect 6699 2036 6765 2070
rect 6799 2036 6830 2070
rect 1278 1970 6830 2036
rect 1278 1936 2101 1970
rect 2135 1936 2201 1970
rect 2235 1936 2301 1970
rect 2335 1936 2401 1970
rect 2435 1936 2501 1970
rect 2535 1936 2601 1970
rect 2635 1936 3489 1970
rect 3523 1936 3589 1970
rect 3623 1936 3689 1970
rect 3723 1936 3789 1970
rect 3823 1936 3889 1970
rect 3923 1936 3989 1970
rect 4023 1936 4877 1970
rect 4911 1936 4977 1970
rect 5011 1936 5077 1970
rect 5111 1936 5177 1970
rect 5211 1936 5277 1970
rect 5311 1936 5377 1970
rect 5411 1936 6265 1970
rect 6299 1936 6365 1970
rect 6399 1936 6465 1970
rect 6499 1936 6565 1970
rect 6599 1936 6665 1970
rect 6699 1936 6765 1970
rect 6799 1936 6830 1970
rect 1278 1905 6830 1936
rect 1278 1904 6566 1905
<< via1 >>
rect -17355 22379 -16923 22395
rect -17355 22341 -17337 22379
rect -17337 22341 -16940 22379
rect -16940 22341 -16923 22379
rect -17355 22325 -16923 22341
rect -13001 22379 -12949 22386
rect -13001 22341 -12949 22379
rect -17355 22213 -16923 22229
rect -17355 22175 -17337 22213
rect -17337 22175 -16940 22213
rect -16940 22175 -16923 22213
rect -17355 22159 -16923 22175
rect -13193 22213 -13141 22220
rect -13001 22334 -12949 22341
rect -8857 22379 -8805 22386
rect -8857 22341 -8805 22379
rect -8857 22334 -8805 22341
rect -4329 22379 -4277 22386
rect -4329 22341 -4277 22379
rect -13193 22175 -13141 22213
rect -13193 22168 -13141 22175
rect -8665 22213 -8613 22220
rect -8665 22175 -8613 22213
rect -8665 22168 -8613 22175
rect -4521 22213 -4469 22220
rect -4329 22334 -4277 22341
rect -185 22379 -133 22386
rect -185 22341 -133 22379
rect -185 22334 -133 22341
rect 4343 22379 4395 22386
rect 4343 22341 4395 22379
rect -4521 22175 -4469 22213
rect -4521 22168 -4469 22175
rect 7 22213 59 22220
rect 7 22175 59 22213
rect 7 22168 59 22175
rect 4151 22213 4203 22220
rect 4343 22334 4395 22341
rect 8487 22379 8539 22386
rect 8487 22341 8539 22379
rect 8487 22334 8539 22341
rect 4151 22175 4203 22213
rect 4151 22168 4203 22175
rect -13001 22047 -12949 22054
rect -13001 22009 -12949 22047
rect -13193 21881 -13141 21888
rect -13001 22002 -12949 22009
rect -8857 22047 -8805 22054
rect -8857 22009 -8805 22047
rect -8857 22002 -8805 22009
rect -4329 22047 -4277 22054
rect -4329 22009 -4277 22047
rect -4329 22002 -4277 22009
rect -185 22047 -133 22054
rect -185 22009 -133 22047
rect -185 22002 -133 22009
rect 352 22047 404 22054
rect 352 22009 404 22047
rect 352 22002 404 22009
rect 4343 22047 4395 22054
rect 4343 22009 4395 22047
rect -13193 21843 -13141 21881
rect -13193 21836 -13141 21843
rect -8665 21881 -8613 21888
rect -8665 21843 -8613 21881
rect -8665 21836 -8613 21843
rect -4521 21881 -4469 21888
rect -4521 21843 -4469 21881
rect -4521 21836 -4469 21843
rect -530 21881 -133 21888
rect -530 21843 -133 21881
rect -530 21836 -133 21843
rect 7 21881 59 21888
rect 7 21843 59 21881
rect 7 21836 59 21843
rect 4151 21881 4203 21888
rect 4343 22002 4395 22009
rect 8487 22047 8539 22054
rect 8487 22009 8539 22047
rect 8487 22002 8539 22009
rect 4151 21843 4203 21881
rect 4151 21836 4203 21843
rect 4688 21881 4740 21888
rect 4688 21843 4740 21881
rect 4688 21836 4740 21843
rect -13193 21715 -13141 21722
rect -13193 21677 -13141 21715
rect -13193 21670 -13141 21677
rect -8665 21715 -8613 21722
rect -8665 21677 -8613 21715
rect -13001 21549 -12949 21556
rect -13001 21511 -12949 21549
rect -13001 21504 -12949 21511
rect -8857 21549 -8805 21556
rect -8665 21670 -8613 21677
rect 7 21715 59 21722
rect 7 21677 59 21715
rect 7 21670 59 21677
rect 4151 21715 4203 21722
rect 4151 21677 4203 21715
rect 4151 21670 4203 21677
rect -8857 21511 -8805 21549
rect -8857 21504 -8805 21511
rect -4329 21549 -4277 21556
rect -4329 21511 -4277 21549
rect -4329 21504 -4277 21511
rect -185 21549 -133 21556
rect -185 21511 -133 21549
rect -185 21504 -133 21511
rect 4343 21549 4395 21556
rect 4343 21511 4395 21549
rect 4343 21504 4395 21511
rect 8487 21549 8539 21556
rect 8487 21511 8539 21549
rect 8487 21504 8539 21511
rect -17064 21383 -16940 21390
rect -17064 21345 -16940 21383
rect -17064 21338 -16940 21345
rect -13193 21383 -13141 21390
rect -13193 21345 -13141 21383
rect -13193 21338 -13141 21345
rect -8665 21383 -8613 21390
rect -8665 21345 -8613 21383
rect -17326 21217 -17254 21234
rect -17326 21179 -17254 21217
rect -17326 21162 -17254 21179
rect -13001 21217 -12949 21224
rect -13001 21179 -12949 21217
rect -13001 21172 -12949 21179
rect -8857 21217 -8805 21224
rect -8665 21338 -8613 21345
rect -4521 21383 -4469 21390
rect -4521 21345 -4469 21383
rect -4521 21338 -4469 21345
rect 7 21383 59 21390
rect 7 21345 59 21383
rect -8857 21179 -8805 21217
rect -8857 21172 -8805 21179
rect -4329 21217 -4277 21224
rect -4329 21179 -4277 21217
rect -4329 21172 -4277 21179
rect -185 21217 -133 21224
rect 7 21338 59 21345
rect 4151 21383 4203 21390
rect 4151 21345 4203 21383
rect 4151 21338 4203 21345
rect -185 21179 -133 21217
rect -185 21172 -133 21179
rect 4343 21217 4395 21224
rect 4343 21179 4395 21217
rect 4343 21172 4395 21179
rect 8487 21217 8539 21224
rect 8487 21179 8539 21217
rect 8487 21172 8539 21179
rect -17402 20077 -16759 20218
rect -13001 19653 -12604 19660
rect -13001 19615 -12604 19653
rect -13001 19608 -12604 19615
rect -1351 19123 257 19175
rect 1265 19123 2873 19175
rect -6844 18753 -6792 18760
rect -6844 18715 -6792 18753
rect -6844 18708 -6792 18715
rect -4765 18753 -4713 18760
rect -4765 18715 -4713 18753
rect -4765 18708 -4713 18715
rect -7017 18587 -6965 18594
rect -7017 18549 -6965 18587
rect -7017 18542 -6965 18549
rect -4593 18587 -4541 18594
rect -4401 18753 -4349 18760
rect -4401 18715 -4349 18753
rect -4401 18708 -4349 18715
rect -1977 18753 -1925 18760
rect -1977 18715 -1925 18753
rect -1977 18708 -1925 18715
rect 831 18753 883 18760
rect 831 18715 883 18753
rect -4593 18549 -4541 18587
rect -4593 18542 -4541 18549
rect -1785 18587 -1733 18594
rect -1785 18549 -1733 18587
rect -7734 18369 -7668 18435
rect -4401 18421 -4349 18428
rect -4401 18383 -4349 18421
rect -7017 18255 -6965 18262
rect -7017 18217 -6965 18255
rect -7017 18210 -6965 18217
rect -4593 18255 -4541 18262
rect -4401 18376 -4349 18383
rect -1977 18421 -1925 18428
rect -1785 18542 -1733 18549
rect 639 18587 691 18594
rect 831 18708 883 18715
rect 3255 18753 3307 18760
rect 3255 18715 3307 18753
rect 3255 18708 3307 18715
rect 6063 18753 6115 18760
rect 6063 18715 6115 18753
rect 639 18549 691 18587
rect 639 18542 691 18549
rect 3447 18587 3499 18594
rect 3447 18549 3499 18587
rect -1977 18383 -1925 18421
rect -1977 18376 -1925 18383
rect 831 18421 883 18428
rect 831 18383 883 18421
rect -4593 18217 -4541 18255
rect -4593 18210 -4541 18217
rect -1785 18255 -1733 18262
rect -1785 18217 -1733 18255
rect -1785 18210 -1733 18217
rect 639 18255 691 18262
rect 831 18376 883 18383
rect 3255 18421 3307 18428
rect 3447 18542 3499 18549
rect 5871 18587 5923 18594
rect 6063 18708 6115 18715
rect 8487 18753 8539 18760
rect 8487 18715 8539 18753
rect 8487 18708 8539 18715
rect 5871 18549 5923 18587
rect 5871 18542 5923 18549
rect 3255 18383 3307 18421
rect 3255 18376 3307 18383
rect 6063 18421 6115 18428
rect 6063 18383 6115 18421
rect 639 18217 691 18255
rect 639 18210 691 18217
rect 3447 18255 3499 18262
rect 3447 18217 3499 18255
rect 3447 18210 3499 18217
rect 5871 18255 5923 18262
rect 5871 18217 5923 18255
rect 5871 18210 5923 18217
rect 6063 18376 6115 18383
rect 8487 18421 8539 18428
rect 8487 18383 8539 18421
rect 8487 18376 8539 18383
rect 6236 18255 6288 18262
rect 6236 18217 6288 18255
rect 6236 18210 6288 18217
rect 8315 18255 8367 18262
rect 8315 18217 8367 18255
rect 8315 18210 8367 18217
rect -7017 17923 -6965 17930
rect -7017 17885 -6965 17923
rect -7017 17878 -6965 17885
rect -4593 17923 -4541 17930
rect -4593 17885 -4541 17923
rect -4593 17878 -4541 17885
rect -16438 17278 -16429 17454
rect -16429 17278 -16395 17454
rect -16395 17278 -16386 17454
rect -14380 17278 -14371 17454
rect -14371 17278 -14337 17454
rect -14337 17278 -14328 17454
rect -10264 17278 -10255 17454
rect -10255 17278 -10221 17454
rect -10221 17278 -10212 17454
rect -8206 17278 -8197 17454
rect -8197 17278 -8163 17454
rect -8163 17278 -8154 17454
rect -15875 17068 -14891 17077
rect -9701 17068 -8717 17077
rect -15875 17034 -14891 17068
rect -9701 17034 -8717 17068
rect -15875 17025 -14891 17034
rect -9701 17025 -8717 17034
rect -16517 16799 -16483 16975
rect -16483 16799 -16429 16975
rect -16429 16799 -16395 16975
rect -14380 16799 -14371 16975
rect -14371 16799 -14337 16975
rect -14337 16799 -14328 16975
rect -12322 16799 -12313 16975
rect -12313 16799 -12279 16975
rect -12279 16799 -12270 16975
rect -10264 16799 -10255 16975
rect -10255 16799 -10221 16975
rect -10221 16799 -10212 16975
rect -16614 16725 -16562 16777
rect -16438 16626 -16386 16678
rect -8030 16725 -7978 16777
rect -16614 16527 -16562 16579
rect -8206 16626 -8154 16678
rect -14380 16329 -14371 16505
rect -14371 16329 -14337 16505
rect -14337 16329 -14328 16505
rect -12322 16329 -12313 16505
rect -12313 16329 -12279 16505
rect -12279 16329 -12270 16505
rect -10264 16329 -10255 16505
rect -10255 16329 -10221 16505
rect -10221 16329 -10212 16505
rect -8030 16527 -7978 16579
rect -8030 16339 -7978 16391
rect -15875 16270 -14891 16279
rect -9701 16270 -8717 16279
rect -15875 16236 -14891 16270
rect -9701 16236 -8717 16270
rect -15875 16227 -14891 16236
rect -9701 16227 -8717 16236
rect -16438 15850 -16429 16026
rect -16429 15850 -16395 16026
rect -16395 15850 -16386 16026
rect -14380 15850 -14371 16026
rect -14371 15850 -14337 16026
rect -14337 15850 -14328 16026
rect -10264 15850 -10255 16026
rect -10255 15850 -10221 16026
rect -10221 15850 -10212 16026
rect -8206 15850 -8197 16026
rect -8197 15850 -8163 16026
rect -8163 15850 -8154 16026
rect -7417 17184 -7408 17360
rect -7408 17184 -7374 17360
rect -7374 17184 -7365 17360
rect -5359 17184 -5350 17360
rect -5350 17184 -5316 17360
rect -5316 17184 -5307 17360
rect -5359 16752 -5350 16928
rect -5350 16752 -5316 16928
rect -5316 16752 -5307 16928
rect -3301 16752 -3292 16928
rect -3292 16752 -3258 16928
rect -3258 16752 -3249 16928
rect -7592 16668 -7540 16720
rect -3126 16668 -3074 16720
rect -7592 16490 -7540 16542
rect -3126 16490 -3074 16542
rect -7417 16282 -7408 16458
rect -7408 16282 -7374 16458
rect -7374 16282 -7365 16458
rect -5359 16282 -5350 16458
rect -5350 16282 -5316 16458
rect -5316 16282 -5307 16458
rect -3292 16282 -3258 16458
rect -3258 16282 -3240 16458
rect -5359 15850 -5350 16026
rect -5350 15850 -5316 16026
rect -5316 15850 -5307 16026
rect -3301 15850 -3292 16026
rect -3292 15850 -3258 16026
rect -3258 15850 -3249 16026
rect -2178 17275 -2044 17409
rect -1091 17171 -1039 17223
rect -575 17171 -523 17223
rect -978 16904 -894 16913
rect -978 16870 -894 16904
rect -978 16861 -894 16870
rect 43 17276 95 17452
rect 4151 17276 4166 17452
rect 4166 17276 4200 17452
rect 4200 17276 4215 17452
rect 43 16882 95 17058
rect 8383 16882 8435 17058
rect 43 16488 95 16664
rect 8383 16488 8435 16664
rect -92 16094 -58 16270
rect -58 16094 -40 16270
rect 4263 16094 4278 16270
rect 4278 16094 4312 16270
rect 4312 16094 4327 16270
rect 8383 16094 8435 16270
rect -11726 15505 -10742 15514
rect -11726 15471 -10742 15505
rect -11726 15462 -10742 15471
rect -9668 15505 -8684 15514
rect -9668 15471 -8684 15505
rect -9668 15462 -8684 15471
rect -10231 15236 -10222 15412
rect -10222 15236 -10188 15412
rect -10188 15236 -10179 15412
rect -12377 15144 -12325 15153
rect -12377 15110 -12368 15144
rect -12368 15110 -12334 15144
rect -12334 15110 -12325 15144
rect -12377 15101 -12325 15110
rect -10231 14842 -10222 15018
rect -10222 14842 -10188 15018
rect -10188 14842 -10179 15018
rect -7462 15301 -7428 15477
rect -7428 15301 -7410 15477
rect -5325 15301 -5316 15465
rect -5316 15301 -5282 15465
rect -5282 15301 -5273 15465
rect -5325 15289 -5273 15301
rect -3179 15351 -3170 15423
rect -3170 15351 -3136 15423
rect -3136 15351 -3127 15423
rect -5325 14825 -5316 15001
rect -5316 14825 -5282 15001
rect -5282 14825 -5273 15001
rect -3180 14882 -3170 14942
rect -3170 14882 -3136 14942
rect -3136 14882 -3128 14942
rect -1062 15551 -1010 15558
rect -1062 15513 -1010 15551
rect -1062 15506 -1010 15513
rect 774 15551 826 15558
rect 774 15513 826 15551
rect 582 15385 634 15392
rect 774 15506 826 15513
rect 2420 15551 2472 15558
rect 2420 15513 2470 15551
rect 2470 15513 2472 15551
rect 2420 15506 2472 15513
rect 582 15347 634 15385
rect 582 15340 634 15347
rect 2073 15385 2193 15392
rect 2073 15347 2193 15385
rect 582 15219 634 15226
rect 2073 15340 2193 15347
rect 582 15181 634 15219
rect 582 15174 634 15181
rect 2073 15219 2193 15226
rect 2073 15181 2193 15219
rect -1062 15053 -1010 15060
rect 2073 15174 2193 15181
rect -1062 15015 -1010 15053
rect -1062 15008 -1010 15015
rect 774 15053 826 15060
rect 774 15015 826 15053
rect 774 15008 826 15015
rect 2418 15053 2470 15060
rect 2418 15015 2470 15053
rect 2418 15008 2470 15015
rect 4264 15821 4328 15885
rect 2709 15246 2773 15310
rect 3805 15618 5089 15627
rect 3805 15584 5089 15618
rect 3805 15575 5089 15584
rect 3092 15378 3101 15534
rect 3101 15378 3135 15534
rect 3135 15378 3144 15534
rect 8379 15650 8439 15710
rect 6463 15618 7747 15629
rect 6463 15584 7747 15618
rect 6463 15573 7747 15584
rect 8408 15378 8417 15534
rect 8417 15378 8451 15534
rect 8451 15378 8460 15534
rect 6463 15328 7747 15337
rect 6463 15294 7747 15328
rect 6463 15285 7747 15294
rect 3805 15186 5089 15195
rect 3805 15152 5089 15186
rect 3805 15143 5089 15152
rect 3092 14946 3101 15102
rect 3101 14946 3135 15102
rect 3135 14946 3144 15102
rect 8408 14946 8417 15102
rect 8417 14946 8451 15102
rect 8451 14946 8460 15102
rect 783 11390 792 12166
rect 792 11390 826 12166
rect 826 11390 835 12166
rect 1041 11390 1050 12166
rect 1050 11390 1084 12166
rect 1084 11390 1093 12166
rect 1041 10396 1050 11172
rect 1050 10396 1084 11172
rect 1084 10396 1093 11172
rect 1933 11390 1942 12166
rect 1942 11390 1976 12166
rect 1976 11390 1985 12166
rect 1596 11298 1718 11307
rect 1596 11264 1630 11298
rect 1630 11264 1718 11298
rect 1596 11255 1718 11264
rect 1933 10396 1942 11172
rect 1942 10396 1976 11172
rect 1976 10396 1985 11172
rect 2825 11390 2834 12166
rect 2834 11390 2868 12166
rect 2868 11390 2877 12166
rect 2488 11298 2610 11307
rect 2488 11264 2522 11298
rect 2522 11264 2610 11298
rect 2488 11255 2610 11264
rect 2825 10396 2834 11172
rect 2834 10396 2868 11172
rect 2868 10396 2877 11172
rect 3717 11390 3726 12166
rect 3726 11390 3760 12166
rect 3760 11390 3769 12166
rect 4428 11855 4604 11864
rect 4428 11821 4604 11855
rect 4428 11812 4604 11821
rect 4428 11509 4604 11518
rect 4428 11475 4604 11509
rect 4428 11466 4604 11475
rect 3380 11298 3502 11307
rect 3380 11264 3414 11298
rect 3414 11264 3502 11298
rect 3380 11255 3502 11264
rect 4645 11255 4697 11307
rect 3717 10396 3726 11172
rect 3726 10396 3760 11172
rect 3760 10396 3769 11172
rect 5001 11266 5377 11275
rect 5001 11232 5377 11266
rect 5001 11223 5377 11232
rect 5595 11266 5971 11275
rect 5595 11232 5971 11266
rect 5595 11223 5971 11232
rect 4428 10741 4604 10750
rect 4428 10707 4604 10741
rect 4428 10698 4604 10707
rect 4428 10395 4604 10404
rect 4428 10361 4604 10395
rect 4428 10352 4604 10361
rect 1415 5654 1467 5706
rect 1415 4266 1467 4318
rect 2235 6434 2501 6500
rect 2235 6400 2301 6434
rect 2301 6400 2335 6434
rect 2335 6400 2401 6434
rect 2401 6400 2435 6434
rect 2435 6400 2501 6434
rect 2235 6334 2501 6400
rect 2235 6300 2301 6334
rect 2301 6300 2335 6334
rect 2335 6300 2401 6334
rect 2401 6300 2435 6334
rect 2435 6300 2501 6334
rect 2235 6234 2501 6300
rect 2758 5654 2810 5706
rect 4688 5654 4740 5706
rect 3689 5112 3723 5118
rect 3723 5112 3789 5118
rect 3789 5112 3793 5118
rect 3689 5046 3793 5112
rect 3689 5012 3723 5046
rect 3723 5012 3789 5046
rect 3789 5012 3793 5046
rect 3689 4946 3793 5012
rect 3689 4912 3723 4946
rect 3723 4912 3789 4946
rect 3789 4912 3793 4946
rect 3689 4870 3793 4912
rect 2758 4266 2810 4318
rect 4688 4266 4740 4318
rect 6030 5654 6082 5706
rect 6030 4266 6082 4318
rect 668 2470 1278 2515
rect 668 2436 713 2470
rect 713 2436 747 2470
rect 747 2436 813 2470
rect 813 2436 847 2470
rect 847 2436 913 2470
rect 913 2436 947 2470
rect 947 2436 1013 2470
rect 1013 2436 1047 2470
rect 1047 2436 1113 2470
rect 1113 2436 1147 2470
rect 1147 2436 1213 2470
rect 1213 2436 1247 2470
rect 1247 2436 1278 2470
rect 668 2370 1278 2436
rect 668 2336 713 2370
rect 713 2336 747 2370
rect 747 2336 813 2370
rect 813 2336 847 2370
rect 847 2336 913 2370
rect 913 2336 947 2370
rect 947 2336 1013 2370
rect 1013 2336 1047 2370
rect 1047 2336 1113 2370
rect 1113 2336 1147 2370
rect 1147 2336 1213 2370
rect 1213 2336 1247 2370
rect 1247 2336 1278 2370
rect 668 2270 1278 2336
rect 668 2236 713 2270
rect 713 2236 747 2270
rect 747 2236 813 2270
rect 813 2236 847 2270
rect 847 2236 913 2270
rect 913 2236 947 2270
rect 947 2236 1013 2270
rect 1013 2236 1047 2270
rect 1047 2236 1113 2270
rect 1113 2236 1147 2270
rect 1147 2236 1213 2270
rect 1213 2236 1247 2270
rect 1247 2236 1278 2270
rect 668 2170 1278 2236
rect 668 2136 713 2170
rect 713 2136 747 2170
rect 747 2136 813 2170
rect 813 2136 847 2170
rect 847 2136 913 2170
rect 913 2136 947 2170
rect 947 2136 1013 2170
rect 1013 2136 1047 2170
rect 1047 2136 1113 2170
rect 1113 2136 1147 2170
rect 1147 2136 1213 2170
rect 1213 2136 1247 2170
rect 1247 2136 1278 2170
rect 668 2070 1278 2136
rect 668 2036 713 2070
rect 713 2036 747 2070
rect 747 2036 813 2070
rect 813 2036 847 2070
rect 847 2036 913 2070
rect 913 2036 947 2070
rect 947 2036 1013 2070
rect 1013 2036 1047 2070
rect 1047 2036 1113 2070
rect 1113 2036 1147 2070
rect 1147 2036 1213 2070
rect 1213 2036 1247 2070
rect 1247 2036 1278 2070
rect 668 1970 1278 2036
rect 668 1936 713 1970
rect 713 1936 747 1970
rect 747 1936 813 1970
rect 813 1936 847 1970
rect 847 1936 913 1970
rect 913 1936 947 1970
rect 947 1936 1013 1970
rect 1013 1936 1047 1970
rect 1047 1936 1113 1970
rect 1113 1936 1147 1970
rect 1147 1936 1213 1970
rect 1213 1936 1247 1970
rect 1247 1936 1278 1970
rect 668 1904 1278 1936
<< metal2 >>
rect -17355 22404 -16923 22405
rect -17610 22395 -16923 22404
rect -17610 22394 -17355 22395
rect -17611 22325 -17355 22394
rect -17611 22315 -16923 22325
rect -13097 22334 -13001 22386
rect -12949 22334 -12939 22386
rect -8867 22334 -8857 22386
rect -8805 22334 -8709 22386
rect -17611 22314 -17268 22315
rect -17611 20658 -17487 22314
rect -17355 22229 -16923 22239
rect -13097 22220 -13045 22334
rect -13203 22168 -13193 22220
rect -13141 22168 -13045 22220
rect -8761 22220 -8709 22334
rect -4425 22334 -4329 22386
rect -4277 22334 -4267 22386
rect -195 22334 -185 22386
rect -133 22334 -37 22386
rect -4425 22220 -4373 22334
rect -8761 22168 -8665 22220
rect -8613 22168 -8603 22220
rect -4531 22168 -4521 22220
rect -4469 22168 -4373 22220
rect -89 22220 -37 22334
rect 4247 22334 4343 22386
rect 4395 22334 4405 22386
rect 8477 22334 8487 22386
rect 8539 22334 8635 22386
rect 4247 22220 4299 22334
rect -89 22168 7 22220
rect 59 22168 69 22220
rect 4141 22168 4151 22220
rect 4203 22168 4299 22220
rect -17355 22149 -16923 22159
rect 352 22054 404 22064
rect 8583 22054 8635 22334
rect -13097 22002 -13001 22054
rect -12949 22002 -12939 22054
rect -8867 22002 -8857 22054
rect -8805 22002 -8709 22054
rect -13097 21888 -13045 22002
rect -13203 21836 -13193 21888
rect -13141 21836 -13045 21888
rect -8761 21971 -8709 22002
rect -4425 22002 -4329 22054
rect -4277 22002 -4267 22054
rect -195 22002 -185 22054
rect -133 22002 -37 22054
rect -4425 21971 -4373 22002
rect -8761 21919 -4373 21971
rect -8761 21888 -8709 21919
rect -4425 21888 -4373 21919
rect -8761 21836 -8665 21888
rect -8613 21836 -8603 21888
rect -4531 21836 -4521 21888
rect -4469 21836 -4373 21888
rect -530 21888 -133 21898
rect -89 21888 -37 22002
rect -89 21836 7 21888
rect 59 21836 69 21888
rect -530 21826 -133 21836
rect -8684 21733 -8675 21805
rect -8603 21733 -8594 21805
rect -8675 21722 -8603 21733
rect -13203 21670 -13193 21722
rect -13141 21670 -13045 21722
rect -8675 21670 -8665 21722
rect -8613 21670 -8603 21722
rect -13097 21556 -13045 21670
rect -8761 21587 -4373 21639
rect -8761 21556 -8709 21587
rect -13097 21504 -13001 21556
rect -12949 21504 -12939 21556
rect -8867 21504 -8857 21556
rect -8805 21504 -8709 21556
rect -4425 21556 -4373 21587
rect -4425 21504 -4329 21556
rect -4277 21504 -4267 21556
rect -17064 21390 -16940 21400
rect -13203 21338 -13193 21390
rect -13141 21338 -13045 21390
rect -17326 21234 -17254 21244
rect -17326 21152 -17254 21162
rect -17064 20811 -16940 21338
rect -13097 21224 -13045 21338
rect -8761 21338 -8665 21390
rect -8613 21338 -8603 21390
rect -4531 21338 -4521 21390
rect -4469 21338 -4373 21390
rect -8761 21224 -8709 21338
rect -13097 21172 -13001 21224
rect -12949 21172 -12939 21224
rect -8867 21172 -8857 21224
rect -8805 21172 -8709 21224
rect -4425 21224 -4373 21338
rect -4425 21172 -4329 21224
rect -4277 21172 -4267 21224
rect -17064 20697 -17059 20811
rect -16945 20697 -16940 20811
rect -364 20808 -298 21826
rect -89 21670 7 21722
rect 59 21670 69 21722
rect -89 21556 -37 21670
rect -195 21504 -185 21556
rect -133 21504 -37 21556
rect -89 21338 7 21390
rect 59 21338 69 21390
rect -89 21224 -37 21338
rect -195 21172 -185 21224
rect -133 21172 -37 21224
rect 352 21154 404 22002
rect 4247 22002 4343 22054
rect 4395 22002 4405 22054
rect 8477 22002 8487 22054
rect 8539 22002 8635 22054
rect 4247 21888 4299 22002
rect 4141 21836 4151 21888
rect 4203 21836 4299 21888
rect 4688 21888 4740 21898
rect 4141 21670 4151 21722
rect 4203 21670 4299 21722
rect 4247 21556 4299 21670
rect 4247 21504 4343 21556
rect 4395 21504 4405 21556
rect 4141 21338 4151 21390
rect 4203 21338 4299 21390
rect 4247 21224 4299 21338
rect 4247 21172 4343 21224
rect 4395 21172 4405 21224
rect 348 21145 408 21154
rect 348 21076 408 21085
rect 4688 20938 4740 21836
rect 8477 21504 8487 21556
rect 8539 21504 8635 21556
rect 8583 21224 8635 21504
rect 8477 21172 8487 21224
rect 8539 21172 8635 21224
rect 4675 20878 4684 20938
rect 4744 20878 4753 20938
rect -364 20752 -359 20808
rect -303 20752 -298 20808
rect -364 20747 -298 20752
rect -359 20743 -303 20747
rect -17064 20692 -16940 20697
rect -17059 20688 -16945 20692
rect -17611 20534 -16542 20658
rect -17402 20218 -16759 20228
rect -17402 20067 -16759 20077
rect -16666 17149 -16542 20534
rect -13001 19660 -12604 19670
rect -13001 19598 -12604 19608
rect -12694 18926 -12634 19598
rect -8763 19438 -8703 19447
rect -8763 19260 -8703 19378
rect -8763 19200 -7242 19260
rect -7626 19128 -7502 19138
rect -7378 19004 -7369 19128
rect -7626 18994 -7502 19004
rect -7878 18926 -7822 18933
rect -12694 18924 -7820 18926
rect -12694 18868 -7878 18924
rect -7822 18868 -7820 18924
rect -12694 18866 -7820 18868
rect -7878 18859 -7822 18866
rect -7734 18435 -7668 18445
rect -7734 18359 -7668 18369
rect -7502 17594 -7378 18880
rect -7302 17711 -7242 19200
rect -4497 19123 -1351 19175
rect 257 19123 1265 19175
rect 2873 19123 6019 19175
rect -6856 18706 -6846 18762
rect -6790 18706 -6780 18762
rect -4777 18706 -4767 18762
rect -4711 18706 -4701 18762
rect -7029 18540 -7019 18596
rect -6963 18540 -6953 18596
rect -4605 18540 -4595 18596
rect -4539 18540 -4529 18596
rect -4497 18428 -4445 19123
rect -4413 18706 -4403 18762
rect -4347 18706 -4337 18762
rect -1989 18706 -1979 18762
rect -1923 18706 -1913 18762
rect 735 18760 787 19123
rect 5967 18760 6019 19123
rect 735 18708 831 18760
rect 883 18708 893 18760
rect 3245 18708 3255 18760
rect 3307 18708 3403 18760
rect 735 18594 787 18708
rect -1881 18542 -1785 18594
rect -1733 18542 -1723 18594
rect 629 18542 639 18594
rect 691 18542 787 18594
rect -1881 18428 -1829 18542
rect -4497 18376 -4401 18428
rect -4349 18376 -4339 18428
rect -1987 18376 -1977 18428
rect -1925 18376 -1829 18428
rect -4497 18262 -4445 18376
rect -7109 18210 -7017 18262
rect -6965 18210 -6955 18262
rect -4603 18210 -4593 18262
rect -4541 18210 -4445 18262
rect -1881 18262 -1829 18376
rect 735 18428 787 18542
rect 3351 18594 3403 18708
rect 5967 18708 6063 18760
rect 6115 18708 6125 18760
rect 8477 18708 8487 18760
rect 8539 18708 8635 18760
rect 5967 18594 6019 18708
rect 3351 18542 3447 18594
rect 3499 18542 3509 18594
rect 5861 18542 5871 18594
rect 5923 18542 6019 18594
rect 3351 18428 3403 18542
rect 735 18376 831 18428
rect 883 18376 893 18428
rect 3245 18376 3255 18428
rect 3307 18376 3403 18428
rect 735 18262 787 18376
rect -1881 18210 -1785 18262
rect -1733 18210 -1723 18262
rect 629 18210 639 18262
rect 691 18210 787 18262
rect -7109 17847 -7057 18210
rect -7027 17878 -7017 17930
rect -6965 17878 -6955 17930
rect -7027 17847 -6955 17878
rect -4603 17878 -4593 17930
rect -4541 17878 -4531 17930
rect -4603 17847 -4531 17878
rect -1881 17847 -1829 18210
rect -1361 17847 -1351 17854
rect -7109 17795 -1351 17847
rect -1361 17788 -1351 17795
rect 257 17847 267 17854
rect 1255 17847 1265 17854
rect 257 17795 1265 17847
rect 257 17788 267 17795
rect 1255 17788 1265 17795
rect 2873 17847 2883 17854
rect 3351 17847 3403 18376
rect 6051 18374 6061 18430
rect 6117 18374 6127 18430
rect 8475 18374 8485 18430
rect 8541 18374 8551 18430
rect 3435 18208 3445 18264
rect 3501 18208 3511 18264
rect 5859 18208 5869 18264
rect 5925 18208 5935 18264
rect 6224 18208 6234 18264
rect 6290 18208 6300 18264
rect 8303 18208 8313 18264
rect 8369 18208 8379 18264
rect 8583 17847 8635 18708
rect 2873 17795 8635 17847
rect 2873 17788 2883 17795
rect -159 17711 -103 17719
rect -7302 17709 -101 17711
rect -7302 17653 -159 17709
rect -103 17653 -94 17709
rect -7302 17651 -101 17653
rect -159 17643 -103 17651
rect -1777 17594 -1549 17599
rect -7502 17589 -1544 17594
rect -16438 17504 -8154 17556
rect -16438 17464 -16386 17504
rect -8206 17464 -8154 17504
rect -7502 17475 -1777 17589
rect -1549 17475 -1540 17589
rect -7502 17470 -1663 17475
rect -1777 17465 -1663 17470
rect -16440 17454 -16384 17464
rect -16440 17268 -16384 17278
rect -14380 17454 -14328 17464
rect -16666 17025 -16394 17149
rect -16518 16975 -16394 17025
rect -15875 17079 -14891 17089
rect -15875 17013 -14891 17023
rect -16518 16800 -16517 16975
rect -16395 16800 -16394 16975
rect -14380 16975 -14328 17278
rect -10264 17454 -10212 17464
rect -16517 16789 -16395 16799
rect -16620 16777 -16556 16783
rect -16620 16725 -16614 16777
rect -16562 16725 -16556 16777
rect -16620 16719 -16556 16725
rect -16611 16585 -16565 16719
rect -16440 16680 -16384 16690
rect -16440 16614 -16384 16624
rect -16620 16579 -16556 16585
rect -16620 16527 -16614 16579
rect -16562 16527 -16556 16579
rect -16620 16521 -16556 16527
rect -14380 16505 -14328 16799
rect -12324 16975 -12268 16985
rect -12324 16974 -12322 16975
rect -12270 16974 -12268 16975
rect -12324 16789 -12268 16799
rect -10264 16975 -10212 17278
rect -8208 17454 -8152 17464
rect -2178 17409 -2044 17419
rect -8208 17268 -8152 17278
rect -7419 17360 -7363 17370
rect -7419 17174 -7363 17184
rect -5359 17360 -5307 17370
rect -2182 17280 -2178 17404
rect -2044 17280 -2040 17404
rect -1549 17470 -1544 17475
rect -1663 17351 -1549 17361
rect 43 17452 95 17462
rect -2178 17265 -2044 17275
rect -2842 17233 -2770 17242
rect -5307 17184 -5305 17224
rect -9701 17079 -8717 17089
rect -9701 17013 -8717 17023
rect -5359 16938 -5305 17184
rect -2770 17223 -523 17233
rect -2770 17171 -1091 17223
rect -1039 17171 -575 17223
rect 43 17193 95 17276
rect 4151 17452 4215 17462
rect 4151 17266 4215 17276
rect -2770 17161 -523 17171
rect -2842 17152 -2770 17161
rect -170 17141 8648 17193
rect -15875 16281 -14891 16291
rect -15875 16215 -14891 16225
rect -16440 16026 -16384 16036
rect -16440 15840 -16384 15850
rect -14380 16026 -14328 16329
rect -12322 16505 -12270 16789
rect -12322 16319 -12270 16329
rect -10264 16505 -10212 16799
rect -5361 16928 -5305 16938
rect -8036 16777 -7972 16783
rect -8036 16725 -8030 16777
rect -7978 16725 -7972 16777
rect -5361 16742 -5305 16752
rect -3301 16928 -3249 16938
rect -1120 16857 -1111 16917
rect -1051 16913 -1042 16917
rect -978 16913 -894 16923
rect -1051 16861 -978 16913
rect -1051 16857 -1042 16861
rect -3249 16855 -1364 16857
rect -3249 16799 -1422 16855
rect -1366 16799 -1357 16855
rect -978 16851 -894 16861
rect -1281 16803 -1221 16812
rect -3249 16797 -1364 16799
rect -8036 16719 -7972 16725
rect -7598 16720 -7534 16726
rect -8208 16680 -8152 16690
rect -8208 16614 -8152 16624
rect -8027 16585 -7981 16719
rect -7598 16668 -7592 16720
rect -7540 16668 -7534 16720
rect -7598 16662 -7534 16668
rect -8036 16579 -7972 16585
rect -8036 16527 -8030 16579
rect -7978 16527 -7972 16579
rect -7589 16548 -7543 16662
rect -3301 16631 -3249 16752
rect -1281 16734 -1221 16743
rect -3132 16720 -3068 16726
rect -3132 16668 -3126 16720
rect -3074 16668 -3068 16720
rect -3132 16662 -3068 16668
rect -7417 16579 -3249 16631
rect -3123 16628 -3077 16662
rect -170 16628 -118 17141
rect 41 17058 97 17068
rect 41 16872 97 16882
rect 8383 17058 8435 17068
rect 8383 16799 8435 16882
rect 43 16747 8435 16799
rect 43 16674 95 16747
rect -3123 16582 -118 16628
rect -8036 16521 -7972 16527
rect -7598 16542 -7534 16548
rect -7598 16490 -7592 16542
rect -7540 16490 -7534 16542
rect -7598 16484 -7534 16490
rect -7417 16458 -7365 16579
rect -3123 16548 -3077 16582
rect -3132 16542 -3068 16548
rect -3132 16490 -3126 16542
rect -3074 16490 -3068 16542
rect -3132 16484 -3068 16490
rect -8036 16339 -8030 16391
rect -7978 16339 -7417 16391
rect -14380 15840 -14328 15850
rect -10264 16026 -10212 16329
rect -9701 16281 -8717 16291
rect -7417 16272 -7365 16282
rect -5361 16458 -5305 16468
rect -5361 16272 -5305 16282
rect -3292 16458 -3240 16468
rect -2426 16453 -2366 16462
rect -1668 16453 -1544 16463
rect -1109 16453 -1053 16460
rect -2366 16393 -1668 16453
rect -1544 16451 -1051 16453
rect -1544 16395 -1109 16451
rect -1053 16395 -1051 16451
rect -1544 16393 -1051 16395
rect -170 16405 -118 16582
rect 41 16664 97 16674
rect 41 16478 97 16488
rect 8381 16664 8437 16674
rect 8381 16478 8437 16488
rect 8596 16405 8648 17141
rect -2426 16384 -2366 16393
rect -1668 16383 -1544 16393
rect -1109 16386 -1053 16393
rect -170 16353 8648 16405
rect -3128 16312 -3072 16319
rect -9701 16215 -8717 16225
rect -10264 15840 -10212 15850
rect -8208 16026 -8152 16036
rect -5361 16026 -5307 16272
rect -3292 16173 -3240 16282
rect -3130 16310 -40 16312
rect -3130 16254 -3128 16310
rect -3072 16270 -40 16310
rect -3072 16254 -92 16270
rect -3130 16252 -92 16254
rect -3128 16245 -3072 16252
rect -3292 16121 -236 16173
rect -5361 16008 -5359 16026
rect -8208 15840 -8152 15850
rect -5359 15840 -5307 15850
rect -3303 16026 -3247 16036
rect -288 15929 -236 16121
rect -92 16084 -40 16094
rect 4263 16270 4327 16280
rect 4263 16084 4327 16094
rect 8383 16270 8435 16353
rect 8383 16084 8435 16094
rect -161 16034 -101 16044
rect 6458 16030 6467 16034
rect -101 15978 6467 16030
rect 6458 15974 6467 15978
rect 6527 15974 6536 16034
rect -161 15964 -101 15974
rect 3079 15929 3088 15933
rect -1971 15916 -1875 15926
rect -375 15916 -319 15917
rect -3303 15840 -3247 15850
rect -2977 15856 -2968 15916
rect -2908 15856 -1971 15916
rect -2977 15849 -1971 15856
rect -1875 15914 -318 15916
rect -1875 15858 -1279 15914
rect -1223 15909 -318 15914
rect -1223 15907 -317 15909
rect -1223 15858 -375 15907
rect -1875 15851 -375 15858
rect -319 15851 -317 15907
rect -288 15877 3088 15929
rect 3079 15873 3088 15877
rect 3148 15873 3157 15933
rect 4264 15885 4328 15895
rect -1875 15849 -317 15851
rect -16438 15800 -16386 15840
rect -8206 15800 -8154 15840
rect -1971 15839 -1875 15849
rect -375 15841 -319 15849
rect 4259 15825 4264 15881
rect 4328 15825 4333 15881
rect 4264 15811 4328 15821
rect -16438 15748 -8154 15800
rect -1668 15791 -1544 15801
rect -10820 15658 -10742 15748
rect -9668 15658 -9590 15748
rect -1544 15737 3857 15789
rect -1668 15725 -1544 15735
rect -10820 15656 -2908 15658
rect -10820 15600 -2966 15656
rect -2910 15600 -2901 15656
rect -1424 15653 -1364 15663
rect 2888 15653 2944 15661
rect -10820 15598 -2908 15600
rect -10820 15524 -10742 15598
rect -11726 15514 -10742 15524
rect -11726 15452 -10742 15462
rect -9668 15524 -9590 15598
rect 2879 15651 2944 15653
rect 2879 15649 2888 15651
rect -1364 15597 2888 15649
rect -1424 15583 -1364 15593
rect -1152 15558 -1000 15568
rect -9668 15514 -8684 15524
rect -1152 15506 -1062 15558
rect -1010 15506 -1000 15558
rect -1152 15496 -1000 15506
rect 678 15506 774 15558
rect 826 15506 836 15558
rect -9668 15452 -8684 15462
rect -7889 15431 -7880 15491
rect -7820 15487 -7811 15491
rect -7820 15477 -7410 15487
rect -7820 15435 -7462 15477
rect -7820 15431 -7811 15435
rect -10231 15412 -10179 15422
rect -7462 15291 -7410 15301
rect -5325 15465 -5273 15475
rect -12377 15153 -12325 15163
rect -17788 15101 -12377 15153
rect -12377 15091 -12325 15101
rect -10231 15018 -10179 15236
rect -10231 14832 -10179 14842
rect -3179 15423 -3127 15433
rect -3127 15418 -2770 15423
rect -3127 15356 -2837 15418
rect -2775 15356 -2766 15418
rect -2675 15413 -1322 15418
rect -2679 15357 -2670 15413
rect -2614 15357 -1322 15413
rect -3127 15351 -2770 15356
rect -2675 15352 -1322 15357
rect -1256 15352 -1247 15418
rect -3179 15341 -3127 15351
rect -5325 15001 -5273 15289
rect -1152 15088 -1100 15496
rect 678 15392 730 15506
rect 572 15340 582 15392
rect 634 15340 730 15392
rect 678 15226 730 15340
rect 572 15174 582 15226
rect 634 15174 730 15226
rect -1155 15079 -1065 15088
rect 678 15070 730 15174
rect 2073 15392 2193 15597
rect 2879 15595 2888 15597
rect 2944 15595 2953 15651
rect 3805 15637 3857 15737
rect 8379 15710 8439 15720
rect 8372 15652 8379 15708
rect 8439 15652 8446 15708
rect 6463 15639 6532 15649
rect 8379 15640 8439 15650
rect 3805 15627 5089 15637
rect 2888 15585 2944 15595
rect 3805 15565 5089 15575
rect 6532 15629 7747 15639
rect 6532 15563 7747 15573
rect 2410 15506 2420 15558
rect 2472 15506 2560 15558
rect 6463 15553 6532 15563
rect 2073 15226 2193 15340
rect 2073 15164 2193 15174
rect 2508 15310 2560 15506
rect 3090 15534 3146 15544
rect 3090 15368 3146 15378
rect 8406 15534 8462 15544
rect 8406 15368 8462 15378
rect 5905 15337 7747 15347
rect 2508 15246 2709 15310
rect 2773 15246 2779 15310
rect 5905 15285 6463 15337
rect 5905 15276 7747 15285
rect 5575 15275 7747 15276
rect 2508 15070 2560 15246
rect 5575 15205 5977 15275
rect 3805 15204 5977 15205
rect 3805 15195 5647 15204
rect 5089 15143 5647 15195
rect 3805 15133 5647 15143
rect 2886 15115 2946 15125
rect -1065 15060 -1000 15070
rect 678 15060 826 15070
rect -1065 15008 -1062 15060
rect -1010 15008 -898 15060
rect 678 15008 774 15060
rect -1065 14998 -1000 15008
rect 678 14998 826 15008
rect 2418 15060 2560 15070
rect 2470 15008 2560 15060
rect 2877 15055 2886 15115
rect 2946 15111 2955 15115
rect 3090 15111 3146 15112
rect 2946 15102 3147 15111
rect 2946 15059 3090 15102
rect 2946 15055 2955 15059
rect 2886 15045 2946 15055
rect 2418 14998 2560 15008
rect -1155 14980 -1065 14989
rect -3180 14942 -3128 14952
rect -3128 14940 -2366 14942
rect -3128 14884 -2424 14940
rect -2368 14884 -2359 14940
rect -3128 14882 -2366 14884
rect -3180 14872 -3128 14882
rect -5325 14815 -5273 14825
rect -2187 14813 -2178 14947
rect -2044 14942 -582 14947
rect 3146 15059 3147 15102
rect 8406 15102 8462 15112
rect -2044 14818 -711 14942
rect -587 14818 -578 14942
rect 3090 14936 3146 14946
rect 8406 14936 8462 14946
rect -2044 14813 -582 14818
rect -1668 14715 -1544 14725
rect -7743 14573 -7734 14639
rect -7668 14573 -1739 14639
rect -1805 14306 -1739 14573
rect -1544 14591 -1420 14601
rect -913 14591 -799 14596
rect -1420 14586 -794 14591
rect -1420 14467 -913 14586
rect -1668 14457 -1420 14467
rect -799 14467 -794 14586
rect 776 14582 842 14587
rect 772 14526 781 14582
rect 837 14526 846 14582
rect -913 14348 -799 14358
rect -266 14306 -210 14310
rect -1805 14301 -205 14306
rect -1805 14245 -266 14301
rect -210 14245 -205 14301
rect -1805 14240 -205 14245
rect -266 14236 -210 14240
rect -1322 14020 -415 14025
rect -1326 13964 -1317 14020
rect -1261 13964 -415 14020
rect -1322 13959 -415 13964
rect -349 13959 -340 14025
rect 776 12166 842 14526
rect 4724 14430 4784 14439
rect 4724 14361 4784 14370
rect 2817 14306 2884 14316
rect 4326 14275 4382 14282
rect 2817 14230 2884 14240
rect 4324 14273 4384 14275
rect 1926 14175 1992 14184
rect 1034 14020 1100 14025
rect 1030 13964 1039 14020
rect 1095 13964 1104 14020
rect 776 11390 783 12166
rect 835 11390 842 12166
rect 776 11380 842 11390
rect 1034 12166 1100 13964
rect 1034 11390 1041 12166
rect 1093 11390 1100 12166
rect 1034 11307 1100 11390
rect 1926 12166 1992 14109
rect 1926 11390 1933 12166
rect 1985 11390 1992 12166
rect 1926 11307 1992 11390
rect 2817 12166 2883 14230
rect 4324 14217 4326 14273
rect 4382 14217 4384 14273
rect 2817 11390 2825 12166
rect 2877 11390 2883 12166
rect 2817 11307 2883 11390
rect 3717 12166 3769 12176
rect 1034 11255 1596 11307
rect 1718 11255 1728 11307
rect 1926 11255 2488 11307
rect 2610 11255 2620 11307
rect 2817 11255 3380 11307
rect 3502 11255 3512 11307
rect 1034 11172 1100 11255
rect 1034 10396 1041 11172
rect 1093 10396 1100 11172
rect 1034 10386 1100 10396
rect 1926 11172 1992 11255
rect 1926 10396 1933 11172
rect 1985 10396 1992 11172
rect 1926 10388 1992 10396
rect 2817 11172 2883 11255
rect 2817 10396 2825 11172
rect 2877 10396 2883 11172
rect 1933 10386 1985 10388
rect 2817 10386 2883 10396
rect 3717 11172 3769 11390
rect 4324 10750 4384 14217
rect 4428 11864 4604 11874
rect 4728 11864 4780 14361
rect 4604 11812 4780 11864
rect 4428 11802 4604 11812
rect 4428 11518 4604 11528
rect 4604 11466 4863 11518
rect 4428 11456 4604 11466
rect 4645 11307 4697 11317
rect 4697 11255 4783 11307
rect 4645 11245 4697 11255
rect 4428 10750 4604 10760
rect 4324 10698 4428 10750
rect 4428 10688 4604 10698
rect 4731 10495 4783 11255
rect 4811 10589 4863 11466
rect 4991 11275 9119 11296
rect 4991 11223 5001 11275
rect 5377 11223 5595 11275
rect 5971 11223 9119 11275
rect 4991 11202 9119 11223
rect 4811 10537 9119 10589
rect 4731 10443 9119 10495
rect -1158 9162 -1062 9171
rect -1715 9068 -1629 9072
rect -1720 9066 -1158 9068
rect 3717 9123 3769 10396
rect 4428 10404 4604 10414
rect 4604 10352 9119 10404
rect 4428 10342 4604 10352
rect -1720 9063 -1062 9066
rect -1720 8977 -1715 9063
rect -1629 8977 -1062 9063
rect -1720 8972 -1062 8977
rect -918 8988 -794 8998
rect -725 8989 -716 9123
rect -582 9118 3769 9123
rect -582 8994 2291 9118
rect 2415 8994 3769 9118
rect -582 8989 3769 8994
rect -1715 8968 -1629 8972
rect -794 8864 -670 8874
rect -927 8740 -918 8864
rect -670 8740 3803 8864
rect -918 8730 -670 8740
rect 2235 6500 2501 6510
rect 2235 6224 2501 6234
rect 1405 5654 1415 5706
rect 1467 5654 2758 5706
rect 2810 5654 2820 5706
rect 3679 5118 3803 8740
rect 4678 5654 4688 5706
rect 4740 5654 6030 5706
rect 6082 5654 6092 5706
rect 3679 4870 3689 5118
rect 3793 4870 3803 5118
rect 1405 4266 1415 4318
rect 1467 4266 2758 4318
rect 2810 4266 2820 4318
rect 4678 4266 4688 4318
rect 4740 4266 6030 4318
rect 6082 4266 6092 4318
rect 668 2515 1278 2525
rect 668 1894 1278 1904
<< via2 >>
rect -17355 22159 -16923 22229
rect -8675 21733 -8603 21805
rect -17321 21167 -17259 21229
rect -17059 20697 -16945 20811
rect 348 21085 408 21145
rect 4684 20878 4744 20938
rect -359 20752 -303 20808
rect -17402 20077 -16759 20218
rect -8763 19378 -8703 19438
rect -7626 19004 -7378 19128
rect -7878 18868 -7822 18924
rect -7502 18880 -7378 19004
rect -7734 18369 -7668 18435
rect -6846 18760 -6790 18762
rect -6846 18708 -6844 18760
rect -6844 18708 -6792 18760
rect -6792 18708 -6790 18760
rect -6846 18706 -6790 18708
rect -4767 18760 -4711 18762
rect -4767 18708 -4765 18760
rect -4765 18708 -4713 18760
rect -4713 18708 -4711 18760
rect -4767 18706 -4711 18708
rect -7019 18594 -6963 18596
rect -7019 18542 -7017 18594
rect -7017 18542 -6965 18594
rect -6965 18542 -6963 18594
rect -7019 18540 -6963 18542
rect -4595 18594 -4539 18596
rect -4595 18542 -4593 18594
rect -4593 18542 -4541 18594
rect -4541 18542 -4539 18594
rect -4595 18540 -4539 18542
rect -4403 18760 -4347 18762
rect -4403 18708 -4401 18760
rect -4401 18708 -4349 18760
rect -4349 18708 -4347 18760
rect -4403 18706 -4347 18708
rect -1979 18760 -1923 18762
rect -1979 18708 -1977 18760
rect -1977 18708 -1925 18760
rect -1925 18708 -1923 18760
rect -1979 18706 -1923 18708
rect -1351 17788 257 17854
rect 1265 17788 2873 17854
rect 6061 18428 6117 18430
rect 6061 18376 6063 18428
rect 6063 18376 6115 18428
rect 6115 18376 6117 18428
rect 6061 18374 6117 18376
rect 8485 18428 8541 18430
rect 8485 18376 8487 18428
rect 8487 18376 8539 18428
rect 8539 18376 8541 18428
rect 8485 18374 8541 18376
rect 3445 18262 3501 18264
rect 3445 18210 3447 18262
rect 3447 18210 3499 18262
rect 3499 18210 3501 18262
rect 3445 18208 3501 18210
rect 5869 18262 5925 18264
rect 5869 18210 5871 18262
rect 5871 18210 5923 18262
rect 5923 18210 5925 18262
rect 5869 18208 5925 18210
rect 6234 18262 6290 18264
rect 6234 18210 6236 18262
rect 6236 18210 6288 18262
rect 6288 18210 6290 18262
rect 6234 18208 6290 18210
rect 8313 18262 8369 18264
rect 8313 18210 8315 18262
rect 8315 18210 8367 18262
rect 8367 18210 8369 18262
rect 8313 18208 8369 18210
rect -159 17653 -103 17709
rect -1777 17475 -1549 17589
rect -16440 17278 -16438 17454
rect -16438 17278 -16386 17454
rect -16386 17278 -16384 17454
rect -15875 17077 -14891 17079
rect -15875 17025 -14891 17077
rect -15875 17023 -14891 17025
rect -16440 16678 -16384 16680
rect -16440 16626 -16438 16678
rect -16438 16626 -16386 16678
rect -16386 16626 -16384 16678
rect -16440 16624 -16384 16626
rect -12324 16799 -12322 16974
rect -12322 16799 -12270 16974
rect -12270 16799 -12268 16974
rect -8208 17278 -8206 17454
rect -8206 17278 -8154 17454
rect -8154 17278 -8152 17454
rect -7419 17184 -7417 17360
rect -7417 17184 -7365 17360
rect -7365 17184 -7363 17360
rect -2173 17280 -2049 17404
rect -1663 17361 -1549 17475
rect -9701 17077 -8717 17079
rect -9701 17025 -8717 17077
rect -9701 17023 -8717 17025
rect -2842 17161 -2770 17233
rect 4151 17276 4215 17452
rect -15875 16279 -14891 16281
rect -15875 16227 -14891 16279
rect -15875 16225 -14891 16227
rect -16440 15850 -16438 16026
rect -16438 15850 -16386 16026
rect -16386 15850 -16384 16026
rect -5361 16752 -5359 16928
rect -5359 16752 -5307 16928
rect -5307 16752 -5305 16928
rect -1111 16857 -1051 16917
rect -1422 16799 -1366 16855
rect -8208 16678 -8152 16680
rect -8208 16626 -8206 16678
rect -8206 16626 -8154 16678
rect -8154 16626 -8152 16678
rect -8208 16624 -8152 16626
rect -1281 16743 -1221 16803
rect 41 16882 43 17058
rect 43 16882 95 17058
rect 95 16882 97 17058
rect -9701 16279 -8717 16281
rect -9701 16227 -8717 16279
rect -5361 16282 -5359 16458
rect -5359 16282 -5307 16458
rect -5307 16282 -5305 16458
rect -2426 16393 -2366 16453
rect -1668 16393 -1544 16453
rect -1109 16395 -1053 16451
rect 41 16488 43 16664
rect 43 16488 95 16664
rect 95 16488 97 16664
rect 8381 16488 8383 16664
rect 8383 16488 8435 16664
rect 8435 16488 8437 16664
rect -9701 16225 -8717 16227
rect -8208 15850 -8206 16026
rect -8206 15850 -8154 16026
rect -8154 15850 -8152 16026
rect -3128 16254 -3072 16310
rect -3303 15850 -3301 16026
rect -3301 15850 -3249 16026
rect -3249 15850 -3247 16026
rect 4263 16094 4327 16270
rect -161 15974 -101 16034
rect 6467 15974 6527 16034
rect -2968 15856 -2908 15916
rect -1971 15849 -1875 15916
rect -1279 15858 -1223 15914
rect -375 15851 -319 15907
rect 3088 15873 3148 15933
rect 4264 15821 4328 15885
rect -1668 15735 -1544 15791
rect -2966 15600 -2910 15656
rect -1424 15593 -1364 15653
rect -7880 15431 -7820 15491
rect -2837 15356 -2775 15418
rect -2670 15357 -2614 15413
rect -1322 15352 -1256 15418
rect -1155 14989 -1065 15079
rect 2888 15595 2944 15651
rect 8381 15652 8437 15708
rect 6463 15629 6532 15639
rect 6463 15573 6532 15629
rect 6463 15563 6532 15573
rect 3090 15378 3092 15534
rect 3092 15378 3144 15534
rect 3144 15378 3146 15534
rect 8406 15378 8408 15534
rect 8408 15378 8460 15534
rect 8460 15378 8462 15534
rect 2886 15055 2946 15115
rect -2424 14884 -2368 14940
rect -2178 14813 -2044 14947
rect 3090 14946 3092 15102
rect 3092 14946 3144 15102
rect 3144 14946 3146 15102
rect -711 14818 -587 14942
rect 8406 14946 8408 15102
rect 8408 14946 8460 15102
rect 8460 14946 8462 15102
rect -7734 14573 -7668 14639
rect -1668 14591 -1544 14715
rect -1668 14467 -1420 14591
rect -913 14358 -799 14586
rect 781 14526 837 14582
rect -266 14245 -210 14301
rect -1317 13964 -1261 14020
rect -415 13959 -349 14025
rect 4724 14370 4784 14430
rect 2817 14240 2884 14306
rect 1926 14109 1992 14175
rect 1039 13964 1095 14020
rect 4326 14217 4382 14273
rect -1158 9066 -1062 9162
rect -1715 8977 -1629 9063
rect -716 8989 -582 9123
rect 2291 8994 2415 9118
rect -918 8864 -794 8988
rect -918 8740 -670 8864
rect 2235 6234 2501 6500
rect 668 1904 1278 2515
<< metal3 >>
rect -17365 22232 -16913 22234
rect -17617 22229 -16913 22232
rect -17617 22159 -17355 22229
rect -16923 22159 -16913 22229
rect -17617 22156 -16913 22159
rect -17617 20629 -17541 22156
rect -17365 22154 -16913 22156
rect -8680 21805 -8598 21810
rect -17481 21733 -8675 21805
rect -8603 21733 -8598 21805
rect -17481 21234 -17409 21733
rect -8763 21668 -8598 21733
rect -17481 21229 -17254 21234
rect -17481 21167 -17321 21229
rect -17259 21167 -17254 21229
rect -17481 21162 -17254 21167
rect -17064 20811 -13191 20816
rect -17064 20697 -17059 20811
rect -16945 20697 -13191 20811
rect -17064 20692 -13191 20697
rect -17617 20553 -13377 20629
rect -17412 20218 -16749 20223
rect -17412 20077 -17402 20218
rect -16759 20077 -16749 20218
rect -17412 20072 -16749 20077
rect -13453 18920 -13377 20553
rect -13315 19128 -13191 20692
rect -8763 19443 -8703 21668
rect 343 21145 413 21150
rect 8570 21147 8634 21153
rect 343 21085 348 21145
rect 408 21085 8570 21145
rect 343 21080 413 21085
rect 8570 21077 8634 21083
rect 4679 20938 4749 20943
rect 8427 20938 8433 20940
rect 4679 20878 4684 20938
rect 4744 20878 8433 20938
rect 4679 20873 4749 20878
rect 8427 20876 8433 20878
rect 8497 20876 8503 20940
rect 8309 20813 8373 20818
rect -364 20812 8374 20813
rect -364 20808 8309 20812
rect -364 20752 -359 20808
rect -303 20752 8309 20808
rect -364 20748 8309 20752
rect 8373 20748 8374 20812
rect -364 20747 8374 20748
rect 8309 20742 8373 20747
rect -8768 19438 -8698 19443
rect -8768 19378 -8763 19438
rect -8703 19378 -8698 19438
rect -8768 19373 -8698 19378
rect -1351 19182 257 19192
rect 1265 19182 2873 19192
rect -7636 19128 -7368 19133
rect -13315 19004 -7626 19128
rect -7636 18999 -7502 19004
rect -7883 18924 -7817 18929
rect -13453 18844 -12258 18920
rect -7883 18868 -7878 18924
rect -7822 18868 -7817 18924
rect -7512 18880 -7502 18999
rect -7378 18880 -7368 19128
rect -7512 18875 -7368 18880
rect -7121 19116 -1351 19182
rect 257 19116 1265 19182
rect 2873 19116 8643 19182
rect -7883 18863 -7817 18868
rect -16450 17454 -16374 17459
rect -16450 17278 -16440 17454
rect -16384 17278 -16374 17454
rect -16450 17273 -16374 17278
rect -16442 17164 -16382 17273
rect -16617 17104 -15825 17164
rect -16617 16200 -16557 17104
rect -15885 17084 -15825 17104
rect -15885 17079 -14881 17084
rect -15885 17023 -15875 17079
rect -14891 17023 -14881 17079
rect -15885 17018 -14881 17023
rect -12334 16974 -12258 18844
rect -8218 17454 -8142 17459
rect -8218 17278 -8208 17454
rect -8152 17278 -8142 17454
rect -8218 17273 -8142 17278
rect -8210 17164 -8150 17273
rect -8767 17104 -7975 17164
rect -8767 17084 -8707 17104
rect -9711 17079 -8707 17084
rect -9711 17023 -9701 17079
rect -8717 17023 -8707 17079
rect -9711 17018 -8707 17023
rect -12334 16799 -12324 16974
rect -12268 16799 -12258 16974
rect -12334 16794 -12258 16799
rect -16450 16682 -16374 16685
rect -8218 16682 -8142 16685
rect -16450 16680 -8142 16682
rect -16450 16624 -16440 16680
rect -16384 16624 -8208 16680
rect -8152 16624 -8142 16680
rect -16450 16622 -8142 16624
rect -16450 16619 -16374 16622
rect -8218 16619 -8142 16622
rect -15885 16281 -14881 16286
rect -15885 16225 -15875 16281
rect -14891 16225 -14881 16281
rect -15885 16220 -14881 16225
rect -9711 16281 -8707 16286
rect -9711 16225 -9701 16281
rect -8717 16225 -8707 16281
rect -9711 16220 -8707 16225
rect -15885 16200 -15825 16220
rect -16617 16140 -15825 16200
rect -8767 16200 -8707 16220
rect -8035 16200 -7975 17104
rect -8767 16140 -7975 16200
rect -16442 16031 -16382 16140
rect -8210 16031 -8150 16140
rect -16450 16026 -16374 16031
rect -16450 15850 -16440 16026
rect -16384 15850 -16374 16026
rect -16450 15845 -16374 15850
rect -8218 16026 -8142 16031
rect -8218 15850 -8208 16026
rect -8152 15850 -8142 16026
rect -8218 15845 -8142 15850
rect -7880 15496 -7820 18863
rect -7121 18606 -7045 19116
rect -6850 18772 -6786 18776
rect -4771 18772 -4707 18776
rect -1893 18772 -1817 19116
rect -1351 19106 257 19116
rect 1265 19106 2873 19116
rect -6895 18766 -6741 18772
rect -6895 18702 -6850 18766
rect -6786 18702 -6741 18766
rect -6895 18696 -6741 18702
rect -4816 18766 -4662 18772
rect -4816 18702 -4771 18766
rect -4707 18702 -4662 18766
rect -4816 18696 -4662 18702
rect -4504 18762 -4342 18772
rect -4504 18706 -4403 18762
rect -4347 18706 -4342 18762
rect -6850 18692 -6786 18696
rect -4771 18692 -4707 18696
rect -4504 18684 -4342 18706
rect -1984 18762 -1817 18772
rect -1984 18706 -1979 18762
rect -1923 18706 -1817 18762
rect -1984 18696 -1817 18706
rect -4600 18618 -4342 18684
rect -7121 18596 -6958 18606
rect -7121 18540 -7019 18596
rect -6963 18540 -6958 18596
rect -7121 18530 -6958 18540
rect -4600 18596 -4438 18618
rect -4600 18540 -4595 18596
rect -4539 18540 -4438 18596
rect -4600 18530 -4438 18540
rect -7744 18435 -7658 18440
rect -7744 18369 -7734 18435
rect -7668 18369 -7658 18435
rect -7744 18364 -7658 18369
rect -7885 15491 -7815 15496
rect -7885 15431 -7880 15491
rect -7820 15431 -7815 15491
rect -7885 15426 -7815 15431
rect -7734 14644 -7668 18364
rect -4504 17854 -4438 18530
rect 3339 18274 3415 19116
rect 8567 18440 8643 19116
rect 5960 18430 6122 18440
rect 5960 18374 6061 18430
rect 6117 18374 6122 18430
rect 5960 18352 6122 18374
rect 8480 18430 8643 18440
rect 8480 18374 8485 18430
rect 8541 18374 8643 18430
rect 8480 18364 8643 18374
rect 5864 18286 6122 18352
rect 3339 18264 3506 18274
rect 3339 18208 3445 18264
rect 3501 18208 3506 18264
rect 3339 18198 3506 18208
rect 5864 18264 6026 18286
rect 6230 18274 6294 18278
rect 8309 18274 8373 18278
rect 5864 18208 5869 18264
rect 5925 18208 6026 18264
rect 5864 18198 6026 18208
rect 6185 18268 6339 18274
rect 6185 18204 6230 18268
rect 6294 18204 6339 18268
rect 6185 18198 6339 18204
rect 8265 18268 8418 18274
rect 8265 18204 8309 18268
rect 8373 18204 8418 18268
rect 8265 18198 8418 18204
rect -1356 17854 262 17864
rect 1260 17854 2878 17864
rect 5960 17854 6026 18198
rect 6230 18194 6294 18198
rect 8309 18194 8373 18198
rect -4504 17788 -1351 17854
rect 257 17788 1265 17854
rect 2873 17788 6026 17854
rect -1356 17778 262 17788
rect 1260 17778 2878 17788
rect -2674 17640 -2610 17645
rect -2675 17639 -2609 17640
rect -2675 17575 -2674 17639
rect -2610 17575 -2609 17639
rect -7429 17360 -7353 17365
rect -7429 17184 -7419 17360
rect -7363 17184 -7353 17360
rect -7429 17179 -7353 17184
rect -2847 17233 -2765 17238
rect -7421 17098 -7361 17179
rect -2847 17161 -2842 17233
rect -2770 17161 -2765 17233
rect -2847 17156 -2765 17161
rect -7596 17038 -7361 17098
rect -7596 16635 -7536 17038
rect -5371 16928 -5295 16933
rect -5375 16752 -5365 16928
rect -5301 16752 -5291 16928
rect -5371 16747 -5295 16752
rect -7596 16575 -3070 16635
rect -5371 16458 -5295 16463
rect -5375 16282 -5365 16458
rect -5301 16282 -5291 16458
rect -3130 16315 -3070 16575
rect -3133 16310 -3067 16315
rect -5371 16277 -5295 16282
rect -3133 16254 -3128 16310
rect -3072 16254 -3067 16310
rect -3133 16249 -3067 16254
rect -3130 16172 -3070 16249
rect -3305 16112 -3070 16172
rect -3305 16031 -3245 16112
rect -3313 16026 -3237 16031
rect -3313 15850 -3303 16026
rect -3247 15850 -3237 16026
rect -2973 15916 -2903 15921
rect -2973 15856 -2968 15916
rect -2908 15856 -2903 15916
rect -2973 15851 -2903 15856
rect -3313 15845 -3237 15850
rect -2968 15661 -2908 15851
rect -2971 15656 -2905 15661
rect -2971 15600 -2966 15656
rect -2910 15600 -2905 15656
rect -2971 15595 -2905 15600
rect -2842 15418 -2770 17156
rect -2842 15356 -2837 15418
rect -2775 15356 -2770 15418
rect -2842 15351 -2770 15356
rect -2675 15413 -2609 17575
rect -1787 17589 -1539 17594
rect -1787 17475 -1777 17589
rect -1787 17470 -1663 17475
rect -2178 17404 -2044 17409
rect -2178 17280 -2173 17404
rect -2049 17280 -2044 17404
rect -1673 17361 -1663 17470
rect -1549 17361 -1539 17589
rect -1673 17356 -1539 17361
rect -2431 16453 -2361 16458
rect -2431 16393 -2426 16453
rect -2366 16393 -2361 16453
rect -2431 16388 -2361 16393
rect -2675 15357 -2670 15413
rect -2614 15357 -2609 15413
rect -2675 15352 -2609 15357
rect -2426 14945 -2366 16388
rect -2178 14952 -2044 17280
rect -1668 16458 -1544 17356
rect -1116 16917 -1046 16922
rect -1427 16855 -1361 16860
rect -1427 16799 -1422 16855
rect -1366 16799 -1361 16855
rect -1116 16857 -1111 16917
rect -1051 16857 -1046 16917
rect -1116 16852 -1046 16857
rect -1427 16794 -1361 16799
rect -1286 16803 -1216 16808
rect -1678 16453 -1534 16458
rect -1678 16393 -1668 16453
rect -1544 16393 -1534 16453
rect -1678 16388 -1534 16393
rect -1981 15916 -1865 15921
rect -1981 15849 -1971 15916
rect -1875 15849 -1865 15916
rect -1981 15844 -1865 15849
rect -1971 15205 -1875 15844
rect -1668 15796 -1544 16388
rect -1678 15791 -1534 15796
rect -1678 15735 -1668 15791
rect -1544 15735 -1534 15791
rect -1678 15730 -1534 15735
rect -1980 15111 -1970 15205
rect -1876 15111 -1866 15205
rect -1971 15110 -1875 15111
rect -2183 14947 -2039 14952
rect -2429 14940 -2363 14945
rect -2429 14884 -2424 14940
rect -2368 14884 -2363 14940
rect -2429 14879 -2363 14884
rect -2183 14813 -2178 14947
rect -2044 14813 -2039 14947
rect -2183 14808 -2039 14813
rect -1668 14720 -1544 15730
rect -1424 15658 -1364 16794
rect -1286 16743 -1281 16803
rect -1221 16743 -1216 16803
rect -1286 16738 -1216 16743
rect -1281 15919 -1221 16738
rect -1111 16456 -1051 16852
rect -1114 16451 -1048 16456
rect -1114 16395 -1109 16451
rect -1053 16395 -1048 16451
rect -1114 16390 -1048 16395
rect -1284 15914 -1218 15919
rect -1284 15858 -1279 15914
rect -1223 15858 -1218 15914
rect -1284 15853 -1218 15858
rect -1434 15653 -1354 15658
rect -1434 15593 -1424 15653
rect -1364 15593 -1354 15653
rect -1434 15588 -1354 15593
rect -1327 15418 -1251 15423
rect -1327 15352 -1322 15418
rect -1256 15352 -1251 15418
rect -1327 15347 -1251 15352
rect -1678 14715 -1534 14720
rect -7739 14639 -7663 14644
rect -7739 14573 -7734 14639
rect -7668 14573 -7663 14639
rect -7739 14568 -7663 14573
rect -17654 14454 -13882 14482
rect -17654 11030 -13966 14454
rect -13902 11030 -13882 14454
rect -17654 11002 -13882 11030
rect -13642 14454 -9870 14482
rect -13642 11030 -9954 14454
rect -9890 11030 -9870 14454
rect -13642 11002 -9870 11030
rect -9630 14454 -5858 14482
rect -9630 11030 -5942 14454
rect -5878 11030 -5858 14454
rect -9630 11002 -5858 11030
rect -5618 14454 -1846 14482
rect -1678 14467 -1668 14715
rect -1544 14596 -1534 14715
rect -1544 14591 -1410 14596
rect -1420 14467 -1410 14591
rect -1678 14462 -1410 14467
rect -5618 11030 -1930 14454
rect -1866 11030 -1846 14454
rect -1322 14020 -1256 15347
rect -1160 15079 -1060 15084
rect -1160 14989 -1155 15079
rect -1065 14989 -1060 15079
rect -1160 14984 -1060 14989
rect -1322 13964 -1317 14020
rect -1261 13964 -1256 14020
rect -1322 13959 -1256 13964
rect -5618 11002 -1846 11030
rect -17654 10734 -13882 10762
rect -17654 7310 -13966 10734
rect -13902 7310 -13882 10734
rect -17654 7282 -13882 7310
rect -13642 10734 -9870 10762
rect -13642 7310 -9954 10734
rect -9890 9070 -9870 10734
rect -9630 10734 -5858 10762
rect -9630 9070 -5942 10734
rect -9890 8974 -5942 9070
rect -9890 7310 -9870 8974
rect -13642 7282 -9870 7310
rect -9630 7310 -5942 8974
rect -5878 7310 -5858 10734
rect -9630 7282 -5858 7310
rect -5618 10734 -1846 10762
rect -5618 7310 -1930 10734
rect -1866 7310 -1846 10734
rect -1158 9167 -1062 14984
rect -716 14942 -582 14947
rect -716 14818 -711 14942
rect -587 14818 -582 14942
rect -923 14586 -789 14591
rect -923 14358 -913 14586
rect -799 14358 -789 14586
rect -923 14353 -789 14358
rect -1163 9162 -1057 9167
rect -1719 9068 -1625 9073
rect -1720 9067 -1624 9068
rect -1720 8973 -1719 9067
rect -1625 8973 -1624 9067
rect -1163 9066 -1158 9162
rect -1062 9066 -1057 9162
rect -1163 9061 -1057 9066
rect -918 8993 -794 14353
rect -716 9128 -582 14818
rect -511 14175 -445 17778
rect -169 17709 -93 17714
rect -169 17653 -159 17709
rect -103 17653 -93 17709
rect -169 17648 -93 17653
rect -161 16039 -101 17648
rect 4141 17452 4225 17457
rect 4141 17276 4151 17452
rect 4215 17276 4225 17452
rect 4141 17271 4225 17276
rect 31 17058 107 17063
rect 31 16882 41 17058
rect 97 16882 107 17058
rect 31 16877 107 16882
rect 39 16803 99 16877
rect 39 16743 8439 16803
rect 8379 16669 8439 16743
rect 31 16664 107 16669
rect 31 16488 41 16664
rect 97 16488 107 16664
rect 31 16483 107 16488
rect 8371 16664 8447 16669
rect 8371 16488 8381 16664
rect 8437 16488 8447 16664
rect 8371 16483 8447 16488
rect -171 16034 -91 16039
rect -171 15974 -161 16034
rect -101 15974 -91 16034
rect -171 15969 -91 15974
rect -385 15909 -309 15912
rect 39 15909 99 16483
rect 4253 16270 4337 16275
rect 4253 16094 4263 16270
rect 4327 16094 4337 16270
rect 4253 16089 4337 16094
rect -385 15907 99 15909
rect -385 15851 -375 15907
rect -319 15851 99 15907
rect 3083 15933 3153 15938
rect 3083 15873 3088 15933
rect 3148 15873 3153 15933
rect 4264 15890 4328 16089
rect 6462 16034 6532 16039
rect 6462 15974 6467 16034
rect 6527 15974 6532 16034
rect 3083 15868 3153 15873
rect 4254 15885 4338 15890
rect -385 15849 99 15851
rect -385 15846 -309 15849
rect 2878 15651 2954 15656
rect 2878 15595 2888 15651
rect 2944 15595 2954 15651
rect 2878 15590 2954 15595
rect 2886 15120 2946 15590
rect 3088 15539 3148 15868
rect 4254 15821 4264 15885
rect 4328 15821 4338 15885
rect 4254 15816 4338 15821
rect 6462 15644 6532 15974
rect 8379 15713 8439 16483
rect 8376 15708 8442 15713
rect 8376 15652 8381 15708
rect 8437 15652 8442 15708
rect 8376 15647 8442 15652
rect 6453 15639 6542 15644
rect 6453 15563 6463 15639
rect 6532 15563 6542 15639
rect 6453 15558 6542 15563
rect 3080 15534 3156 15539
rect 8396 15534 8472 15539
rect 3076 15378 3086 15534
rect 3150 15378 3160 15534
rect 8396 15378 8406 15534
rect 8462 15378 8472 15534
rect 3080 15373 3156 15378
rect 8396 15373 8472 15378
rect 8404 15270 8464 15373
rect 3088 15210 8464 15270
rect 2876 15115 2956 15120
rect 2876 15055 2886 15115
rect 2946 15055 2956 15115
rect 3088 15107 3148 15210
rect 2876 15050 2956 15055
rect 3080 15102 3156 15107
rect 8396 15102 8472 15107
rect 3080 14946 3090 15102
rect 3146 14946 3156 15102
rect 8392 14946 8402 15102
rect 8466 14946 8476 15102
rect 3080 14941 3156 14946
rect 8396 14941 8472 14946
rect 776 14586 8593 14587
rect 776 14582 8528 14586
rect 776 14526 781 14582
rect 837 14526 8528 14582
rect 776 14522 8528 14526
rect 8592 14522 8598 14586
rect 776 14521 8593 14522
rect 4719 14430 4789 14435
rect 8646 14430 8652 14432
rect 4719 14370 4724 14430
rect 4784 14370 8652 14430
rect 4719 14365 4789 14370
rect 8646 14368 8652 14370
rect 8716 14368 8722 14432
rect 2807 14306 2894 14311
rect -271 14301 2817 14306
rect -271 14245 -266 14301
rect -210 14245 2817 14301
rect -271 14240 2817 14245
rect 2884 14240 2894 14306
rect 2807 14235 2894 14240
rect 4321 14275 4387 14278
rect 8769 14275 8775 14277
rect 4321 14273 8775 14275
rect 4321 14217 4326 14273
rect 4382 14217 8775 14273
rect 4321 14215 8775 14217
rect 4321 14212 4387 14215
rect 8769 14213 8775 14215
rect 8839 14213 8845 14277
rect 1921 14175 1997 14180
rect -511 14109 1926 14175
rect 1992 14109 1997 14175
rect 1921 14104 1997 14109
rect -420 14025 -344 14030
rect -420 13959 -415 14025
rect -349 14020 1100 14025
rect -349 13964 1039 14020
rect 1095 13964 1100 14020
rect -349 13959 1100 13964
rect -420 13954 -344 13959
rect -721 9123 -577 9128
rect -1720 8972 -1624 8973
rect -928 8988 -784 8993
rect -1719 8967 -1625 8972
rect -928 8740 -918 8988
rect -794 8869 -784 8988
rect -721 8989 -716 9123
rect -582 8989 -577 9123
rect -721 8984 -577 8989
rect 2286 9118 2420 9123
rect 2286 8994 2291 9118
rect 2415 8994 2420 9118
rect -794 8864 -660 8869
rect -670 8740 -660 8864
rect -928 8735 -660 8740
rect 2286 7516 2420 8994
rect -5618 7282 -1846 7310
rect -11971 7042 -11875 7282
rect -7938 7042 -7842 7282
rect -17654 7014 -13882 7042
rect -17654 3590 -13966 7014
rect -13902 3590 -13882 7014
rect -17654 3562 -13882 3590
rect -13642 7014 -9870 7042
rect -13642 3590 -9954 7014
rect -9890 5350 -9870 7014
rect -9630 7014 -5858 7042
rect -9630 5350 -5942 7014
rect -9890 5254 -5942 5350
rect -9890 3590 -9870 5254
rect -13642 3562 -9870 3590
rect -9630 3590 -5942 5254
rect -5878 3590 -5858 7014
rect -9630 3562 -5858 3590
rect -5618 7014 -1846 7042
rect -5618 3590 -1930 7014
rect -1866 3590 -1846 7014
rect 2300 6505 2406 7516
rect 2225 6500 2511 6505
rect 2225 6234 2235 6500
rect 2501 6234 2511 6500
rect 2225 6229 2511 6234
rect -5618 3562 -1846 3590
rect -17654 3294 -13882 3322
rect -17654 -130 -13966 3294
rect -13902 -130 -13882 3294
rect -17654 -158 -13882 -130
rect -13642 3294 -9870 3322
rect -13642 -130 -9954 3294
rect -9890 -130 -9870 3294
rect -13642 -158 -9870 -130
rect -9630 3294 -5858 3322
rect -9630 -130 -5942 3294
rect -5878 -130 -5858 3294
rect -9630 -158 -5858 -130
rect -5618 3294 -1846 3322
rect -5618 -130 -1930 3294
rect -1866 -130 -1846 3294
rect 658 2515 1288 2520
rect 658 1904 668 2515
rect 1278 1904 1288 2515
rect 658 1899 1288 1904
rect -5618 -158 -1846 -130
<< via3 >>
rect -17402 20077 -16759 20218
rect 8570 21083 8634 21147
rect 8433 20876 8497 20940
rect 8309 20748 8373 20812
rect -1351 19116 257 19182
rect 1265 19116 2873 19182
rect -6850 18762 -6786 18766
rect -6850 18706 -6846 18762
rect -6846 18706 -6790 18762
rect -6790 18706 -6786 18762
rect -6850 18702 -6786 18706
rect -4771 18762 -4707 18766
rect -4771 18706 -4767 18762
rect -4767 18706 -4711 18762
rect -4711 18706 -4707 18762
rect -4771 18702 -4707 18706
rect 6230 18264 6294 18268
rect 6230 18208 6234 18264
rect 6234 18208 6290 18264
rect 6290 18208 6294 18264
rect 6230 18204 6294 18208
rect 8309 18264 8373 18268
rect 8309 18208 8313 18264
rect 8313 18208 8369 18264
rect 8369 18208 8373 18264
rect 8309 18204 8373 18208
rect -2674 17575 -2610 17639
rect -5365 16752 -5361 16928
rect -5361 16752 -5305 16928
rect -5305 16752 -5301 16928
rect -5365 16282 -5361 16458
rect -5361 16282 -5305 16458
rect -5305 16282 -5301 16458
rect -1970 15111 -1876 15205
rect -13966 11030 -13902 14454
rect -9954 11030 -9890 14454
rect -5942 11030 -5878 14454
rect -1930 11030 -1866 14454
rect -13966 7310 -13902 10734
rect -9954 7310 -9890 10734
rect -5942 7310 -5878 10734
rect -1930 7310 -1866 10734
rect -1719 9063 -1625 9067
rect -1719 8977 -1715 9063
rect -1715 8977 -1629 9063
rect -1629 8977 -1625 9063
rect -1719 8973 -1625 8977
rect 4151 17276 4215 17452
rect 4263 16094 4327 16270
rect 3086 15378 3090 15534
rect 3090 15378 3146 15534
rect 3146 15378 3150 15534
rect 8402 14946 8406 15102
rect 8406 14946 8462 15102
rect 8462 14946 8466 15102
rect 8528 14522 8592 14586
rect 8652 14368 8716 14432
rect 8775 14213 8839 14277
rect -13966 3590 -13902 7014
rect -9954 3590 -9890 7014
rect -5942 3590 -5878 7014
rect -1930 3590 -1866 7014
rect -13966 -130 -13902 3294
rect -9954 -130 -9890 3294
rect -5942 -130 -5878 3294
rect -1930 -130 -1866 3294
rect 668 1904 1278 2515
<< mimcap >>
rect -17614 14402 -14214 14442
rect -17614 11082 -17574 14402
rect -14254 11082 -14214 14402
rect -17614 11042 -14214 11082
rect -13602 14402 -10202 14442
rect -13602 11082 -13562 14402
rect -10242 11082 -10202 14402
rect -13602 11042 -10202 11082
rect -9590 14402 -6190 14442
rect -9590 11082 -9550 14402
rect -6230 11082 -6190 14402
rect -9590 11042 -6190 11082
rect -5578 14402 -2178 14442
rect -5578 11082 -5538 14402
rect -2218 11082 -2178 14402
rect -5578 11042 -2178 11082
rect -17614 10682 -14214 10722
rect -17614 7362 -17574 10682
rect -14254 7362 -14214 10682
rect -17614 7322 -14214 7362
rect -13602 10682 -10202 10722
rect -13602 7362 -13562 10682
rect -10242 7362 -10202 10682
rect -13602 7322 -10202 7362
rect -9590 10682 -6190 10722
rect -9590 7362 -9550 10682
rect -6230 7362 -6190 10682
rect -9590 7322 -6190 7362
rect -5578 10682 -2178 10722
rect -5578 7362 -5538 10682
rect -2218 7362 -2178 10682
rect -5578 7322 -2178 7362
rect -17614 6962 -14214 7002
rect -17614 3642 -17574 6962
rect -14254 3642 -14214 6962
rect -17614 3602 -14214 3642
rect -13602 6962 -10202 7002
rect -13602 3642 -13562 6962
rect -10242 3642 -10202 6962
rect -13602 3602 -10202 3642
rect -9590 6962 -6190 7002
rect -9590 3642 -9550 6962
rect -6230 3642 -6190 6962
rect -9590 3602 -6190 3642
rect -5578 6962 -2178 7002
rect -5578 3642 -5538 6962
rect -2218 3642 -2178 6962
rect -5578 3602 -2178 3642
rect -17614 3242 -14214 3282
rect -17614 -78 -17574 3242
rect -14254 -78 -14214 3242
rect -17614 -118 -14214 -78
rect -13602 3242 -10202 3282
rect -13602 -78 -13562 3242
rect -10242 -78 -10202 3242
rect -13602 -118 -10202 -78
rect -9590 3242 -6190 3282
rect -9590 -78 -9550 3242
rect -6230 -78 -6190 3242
rect -9590 -118 -6190 -78
rect -5578 3242 -2178 3282
rect -5578 -78 -5538 3242
rect -2218 -78 -2178 3242
rect -5578 -118 -2178 -78
<< mimcapcontact >>
rect -17574 11082 -14254 14402
rect -13562 11082 -10242 14402
rect -9550 11082 -6230 14402
rect -5538 11082 -2218 14402
rect -17574 7362 -14254 10682
rect -13562 7362 -10242 10682
rect -9550 7362 -6230 10682
rect -5538 7362 -2218 10682
rect -17574 3642 -14254 6962
rect -13562 3642 -10242 6962
rect -9550 3642 -6230 6962
rect -5538 3642 -2218 6962
rect -17574 -78 -14254 3242
rect -13562 -78 -10242 3242
rect -9550 -78 -6230 3242
rect -5538 -78 -2218 3242
<< metal4 >>
rect 8569 21147 8635 21148
rect 8569 21083 8570 21147
rect 8634 21083 8635 21147
rect 8569 21082 8635 21083
rect 8432 20940 8498 20941
rect 8432 20876 8433 20940
rect 8497 20876 8498 20940
rect 8432 20875 8498 20876
rect 8308 20812 8374 20813
rect 8308 20748 8309 20812
rect 8373 20748 8374 20812
rect -17403 20218 -16758 20219
rect -17403 20077 -17402 20218
rect -16759 20077 -16758 20218
rect -17403 20076 -16758 20077
rect -17402 14403 -16759 20076
rect -1352 19182 258 19183
rect 1264 19182 2874 19183
rect -6977 19116 -1351 19182
rect 257 19116 1265 19182
rect 2873 19116 6295 19182
rect -6977 17640 -6911 19116
rect -6851 18766 -6785 18767
rect -6851 18702 -6850 18766
rect -6786 18702 -6785 18766
rect -6851 17854 -6785 18702
rect -4772 18766 -4706 19116
rect -1352 19115 258 19116
rect 1264 19115 2874 19116
rect -4772 18702 -4771 18766
rect -4707 18702 -4706 18766
rect -4772 18701 -4706 18702
rect 6229 18268 6295 19116
rect 6229 18204 6230 18268
rect 6294 18204 6295 18268
rect 6229 18203 6295 18204
rect 8308 18268 8374 20748
rect 8308 18204 8309 18268
rect 8373 18204 8374 18268
rect 8308 17854 8374 18204
rect -6851 17788 8374 17854
rect 8308 17675 8374 17788
rect 8435 17808 8495 20875
rect 8572 17957 8632 21082
rect 8572 17897 8837 17957
rect 8435 17748 8714 17808
rect -6977 17639 -2609 17640
rect -6977 17575 -2674 17639
rect -2610 17575 -2609 17639
rect 8308 17609 8593 17675
rect -6977 17574 -2609 17575
rect 4150 17452 4272 17453
rect 4150 17276 4151 17452
rect 4215 17276 4272 17452
rect 4150 17275 4272 17276
rect -5366 16928 -5300 16929
rect -5366 16752 -5365 16928
rect -5301 16752 -5300 16928
rect -5366 16751 -5300 16752
rect -5365 16459 -5301 16751
rect -5366 16458 -5300 16459
rect -5366 16282 -5365 16458
rect -5301 16282 -5300 16458
rect -5366 16281 -5300 16282
rect 4206 16271 4272 17275
rect 4206 16270 4328 16271
rect 4206 16094 4263 16270
rect 4327 16094 4328 16270
rect 4206 16093 4328 16094
rect 3085 15534 3151 15535
rect 3085 15378 3086 15534
rect 3150 15378 3151 15534
rect 3085 15377 3151 15378
rect 3088 15270 3148 15377
rect 3088 15210 8464 15270
rect -1971 15205 -1410 15206
rect -1971 15111 -1970 15205
rect -1876 15111 -1410 15205
rect -1971 15110 -1410 15111
rect -13982 14454 -13886 14470
rect -17575 14402 -14253 14403
rect -17575 11082 -17574 14402
rect -14254 12790 -14253 14402
rect -13982 12790 -13966 14454
rect -14254 12694 -13966 12790
rect -14254 11082 -14253 12694
rect -17575 11081 -14253 11082
rect -16227 10683 -15584 11081
rect -13982 11030 -13966 12694
rect -13902 12790 -13886 14454
rect -9970 14454 -9874 14470
rect -13563 14402 -10241 14403
rect -13563 12790 -13562 14402
rect -13902 12694 -13562 12790
rect -13902 11620 -13886 12694
rect -13902 11030 -13884 11620
rect -13563 11082 -13562 12694
rect -10242 12790 -10241 14402
rect -9970 12790 -9954 14454
rect -10242 12694 -9954 12790
rect -10242 11082 -10241 12694
rect -13563 11081 -10241 11082
rect -13982 10734 -13884 11030
rect -9970 11030 -9954 12694
rect -9890 12790 -9874 14454
rect -5958 14454 -5862 14470
rect -9551 14402 -6229 14403
rect -9551 12790 -9550 14402
rect -9890 12694 -9550 12790
rect -9890 11030 -9874 12694
rect -9551 11082 -9550 12694
rect -6230 12790 -6229 14402
rect -5958 12790 -5942 14454
rect -6230 12694 -5942 12790
rect -6230 11082 -6229 12694
rect -9551 11081 -6229 11082
rect -9970 11014 -9874 11030
rect -5958 11030 -5942 12694
rect -5878 12790 -5862 14454
rect -1946 14454 -1850 14470
rect -5539 14402 -2217 14403
rect -5539 12790 -5538 14402
rect -5878 12694 -5538 12790
rect -5878 11030 -5862 12694
rect -5623 12692 -5538 12694
rect -5539 11082 -5538 12692
rect -2218 12790 -2217 14402
rect -1946 12790 -1930 14454
rect -2218 12692 -1930 12790
rect -2218 11082 -2217 12692
rect -5539 11081 -2217 11082
rect -5958 11014 -5862 11030
rect -1946 11030 -1930 12692
rect -1866 11030 -1850 14454
rect -1946 11014 -1850 11030
rect -17575 10682 -14253 10683
rect -17575 7362 -17574 10682
rect -14254 7362 -14253 10682
rect -17575 7361 -14253 7362
rect -16227 6963 -15584 7361
rect -13982 7310 -13966 10734
rect -13902 7310 -13884 10734
rect -9970 10734 -9874 10750
rect -13563 10682 -10241 10683
rect -13563 7362 -13562 10682
rect -10242 7362 -10241 10682
rect -13563 7361 -10241 7362
rect -13982 7014 -13884 7310
rect -17575 6962 -14253 6963
rect -17575 3642 -17574 6962
rect -14254 3642 -14253 6962
rect -17575 3641 -14253 3642
rect -16227 3243 -15584 3641
rect -13982 3590 -13966 7014
rect -13902 3590 -13884 7014
rect -11971 7210 -11875 7361
rect -9970 7310 -9954 10734
rect -9890 7310 -9874 10734
rect -5958 10734 -5862 10750
rect -9551 10682 -6229 10683
rect -9551 7362 -9550 10682
rect -6230 7362 -6229 10682
rect -9551 7361 -6229 7362
rect -9970 7294 -9874 7310
rect -7938 7210 -7842 7361
rect -5958 7310 -5942 10734
rect -5878 9068 -5862 10734
rect -1946 10734 -1850 10750
rect -5539 10682 -2217 10683
rect -5539 9068 -5538 10682
rect -5878 8972 -5538 9068
rect -5878 7310 -5862 8972
rect -5539 7362 -5538 8972
rect -2218 9068 -2217 10682
rect -1946 9068 -1930 10734
rect -2218 8972 -1930 9068
rect -2218 7362 -2217 8972
rect -5539 7361 -2217 7362
rect -5958 7294 -5862 7310
rect -1946 7310 -1930 8972
rect -1866 9068 -1850 10734
rect -1866 9067 -1624 9068
rect -1866 8973 -1719 9067
rect -1625 8973 -1624 9067
rect -1866 8972 -1624 8973
rect -1866 7310 -1850 8972
rect -1946 7294 -1850 7310
rect -1506 7210 -1410 15110
rect 8404 15103 8464 15210
rect 8401 15102 8467 15103
rect 8401 14946 8402 15102
rect 8466 14946 8467 15102
rect 8401 14945 8467 14946
rect 8527 14586 8593 17609
rect 8527 14522 8528 14586
rect 8592 14522 8593 14586
rect 8527 14521 8593 14522
rect 8654 14433 8714 17748
rect 8651 14432 8717 14433
rect 8651 14368 8652 14432
rect 8716 14368 8717 14432
rect 8651 14367 8717 14368
rect 8777 14278 8837 17897
rect 8774 14277 8840 14278
rect 8774 14213 8775 14277
rect 8839 14213 8840 14277
rect 8774 14212 8840 14213
rect -11971 7114 -1410 7210
rect -11971 6963 -11875 7114
rect -9970 7014 -9874 7030
rect -13563 6962 -10241 6963
rect -13563 3642 -13562 6962
rect -10242 3642 -10241 6962
rect -13563 3641 -10241 3642
rect -13982 3294 -13884 3590
rect -9970 3590 -9954 7014
rect -9890 3590 -9874 7014
rect -7938 6963 -7842 7114
rect -5958 7014 -5862 7030
rect -9551 6962 -6229 6963
rect -9551 3642 -9550 6962
rect -6230 3642 -6229 6962
rect -9551 3641 -6229 3642
rect -9970 3574 -9874 3590
rect -5958 3590 -5942 7014
rect -5878 3590 -5862 7014
rect -1946 7014 -1850 7030
rect -1946 7006 -1930 7014
rect -3926 6963 -3830 7006
rect -5539 6962 -2217 6963
rect -5539 3642 -5538 6962
rect -2218 3642 -2217 6962
rect -5539 3641 -2217 3642
rect -5958 3574 -5862 3590
rect -17575 3242 -14253 3243
rect -17575 -78 -17574 3242
rect -14254 1904 -14253 3242
rect -13982 1904 -13966 3294
rect -14254 1261 -13966 1904
rect -14254 -78 -14253 1261
rect -17575 -79 -14253 -78
rect -13982 -130 -13966 1261
rect -13902 2987 -13884 3294
rect -9970 3294 -9874 3310
rect -13563 3242 -10241 3243
rect -13902 1904 -13886 2987
rect -13563 1904 -13562 3242
rect -13902 1261 -13562 1904
rect -13902 -130 -13886 1261
rect -13563 -78 -13562 1261
rect -10242 1904 -10241 3242
rect -9970 1904 -9954 3294
rect -10242 1261 -9954 1904
rect -10242 -78 -10241 1261
rect -13563 -79 -10241 -78
rect -13982 -146 -13886 -130
rect -9970 -130 -9954 1261
rect -9890 1904 -9874 3294
rect -5958 3294 -5862 3310
rect -9551 3242 -6229 3243
rect -9551 1904 -9550 3242
rect -9890 1261 -9550 1904
rect -9890 -130 -9874 1261
rect -9551 -78 -9550 1261
rect -6230 1904 -6229 3242
rect -5958 1904 -5942 3294
rect -6230 1261 -5942 1904
rect -6230 -78 -6229 1261
rect -9551 -79 -6229 -78
rect -9970 -146 -9874 -130
rect -5958 -130 -5942 1261
rect -5878 1904 -5862 3294
rect -3926 3243 -3830 3641
rect -1947 3590 -1930 7006
rect -1866 7006 -1850 7014
rect -1866 3590 -1849 7006
rect -1947 3294 -1849 3590
rect -5539 3242 -2217 3243
rect -5539 1904 -5538 3242
rect -5878 1261 -5538 1904
rect -5878 -130 -5862 1261
rect -5539 -78 -5538 1261
rect -2218 2487 -2217 3242
rect -1947 3174 -1930 3294
rect -1946 2487 -1930 3174
rect -2218 1261 -1930 2487
rect -2218 -78 -2217 1261
rect -5539 -79 -2217 -78
rect -5958 -146 -5862 -130
rect -1946 -130 -1930 1261
rect -1866 3174 -1849 3294
rect -1866 2487 -1850 3174
rect 667 2515 1279 2516
rect 667 2487 668 2515
rect -1866 1904 668 2487
rect 1278 1904 1279 2515
rect -1866 1903 1279 1904
rect -1866 1873 1208 1903
rect -1866 1846 668 1873
rect -1866 -130 -1850 1846
rect -1946 -146 -1850 -130
<< labels >>
flabel metal4 -17203 19230 -17203 19230 0 FreeSans 1600 0 0 0 AVSS
port 2 nsew
flabel metal2 -16596 19440 -16596 19440 0 FreeSans 1600 0 0 0 VREF
port 3 nsew
flabel metal1 9111 9954 9111 9954 0 FreeSans 160 0 0 0 TRIM3
port 4 nsew
flabel metal1 9111 10033 9111 10033 0 FreeSans 160 0 0 0 TRIM2
port 5 nsew
flabel metal1 9111 10113 9111 10113 0 FreeSans 160 0 0 0 TRIM1
port 6 nsew
flabel metal1 9111 10193 9111 10193 0 FreeSans 160 0 0 0 TRIM0
port 7 nsew
flabel metal2 9111 10379 9111 10379 0 FreeSans 160 0 0 0 VBGSC
port 8 nsew
flabel metal2 9111 10471 9111 10471 0 FreeSans 160 0 0 0 VENA
port 9 nsew
flabel metal2 9111 10564 9111 10564 0 FreeSans 160 0 0 0 VBGTC
port 10 nsew
flabel metal1 9111 10941 9111 10941 0 FreeSans 160 0 0 0 ENA
port 11 nsew
flabel metal2 9111 11252 9111 11252 0 FreeSans 160 0 0 0 AVDD
port 12 nsew
flabel metal1 9110 9871 9110 9871 0 FreeSans 160 0 0 0 DVDD
port 13 nsew
flabel metal1 9110 9790 9110 9790 0 FreeSans 160 0 0 0 DVSS
port 14 nsew
flabel metal2 -17769 15128 -17769 15128 0 FreeSans 160 0 0 0 IPTAT
port 15 nsew
flabel metal2 3772 8637 3772 8637 0 FreeSans 1600 0 0 0 bjt_0.A
flabel metal1 3059 6604 3059 6604 0 FreeSans 1600 0 0 0 bjt_0.B
flabel metal1 4440 7325 4440 7325 0 FreeSans 1600 0 0 0 bjt_0.AVSS
flabel locali 6465 2094 6569 2342 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[0,0].Emitter
flabel locali 5894 2153 5943 2254 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[0,0].Collector
flabel locali 6053 2130 6093 2248 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[0,0].Base
flabel locali 6465 3482 6569 3730 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[0,1].Emitter
flabel locali 5894 3541 5943 3642 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[0,1].Collector
flabel locali 6053 3518 6093 3636 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[0,1].Base
flabel locali 6465 4870 6569 5118 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[0,2].Emitter
flabel locali 5894 4929 5943 5030 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[0,2].Collector
flabel locali 6053 4906 6093 5024 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[0,2].Base
flabel locali 6465 6258 6569 6506 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[0,3].Emitter
flabel locali 5894 6317 5943 6418 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[0,3].Collector
flabel locali 6053 6294 6093 6412 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[0,3].Base
flabel locali 6465 7646 6569 7894 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[0,4].Emitter
flabel locali 5894 7705 5943 7806 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[0,4].Collector
flabel locali 6053 7682 6093 7800 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[0,4].Base
flabel locali 5077 2094 5181 2342 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[1,0].Emitter
flabel locali 4506 2153 4555 2254 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[1,0].Collector
flabel locali 4665 2130 4705 2248 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[1,0].Base
flabel locali 5077 3482 5181 3730 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[1,1].Emitter
flabel locali 4506 3541 4555 3642 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[1,1].Collector
flabel locali 4665 3518 4705 3636 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[1,1].Base
flabel locali 5077 4870 5181 5118 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[1,2].Emitter
flabel locali 4506 4929 4555 5030 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[1,2].Collector
flabel locali 4665 4906 4705 5024 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[1,2].Base
flabel locali 5077 6258 5181 6506 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[1,3].Emitter
flabel locali 4506 6317 4555 6418 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[1,3].Collector
flabel locali 4665 6294 4705 6412 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[1,3].Base
flabel locali 5077 7646 5181 7894 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[1,4].Emitter
flabel locali 4506 7705 4555 7806 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[1,4].Collector
flabel locali 4665 7682 4705 7800 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[1,4].Base
flabel locali 3689 2094 3793 2342 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[2,0].Emitter
flabel locali 3118 2153 3167 2254 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[2,0].Collector
flabel locali 3277 2130 3317 2248 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[2,0].Base
flabel locali 3689 3482 3793 3730 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[2,1].Emitter
flabel locali 3118 3541 3167 3642 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[2,1].Collector
flabel locali 3277 3518 3317 3636 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[2,1].Base
flabel locali 3689 4870 3793 5118 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[2,2].Emitter
flabel locali 3118 4929 3167 5030 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[2,2].Collector
flabel locali 3277 4906 3317 5024 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[2,2].Base
flabel locali 3689 6258 3793 6506 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[2,3].Emitter
flabel locali 3118 6317 3167 6418 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[2,3].Collector
flabel locali 3277 6294 3317 6412 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[2,3].Base
flabel locali 3689 7646 3793 7894 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[2,4].Emitter
flabel locali 3118 7705 3167 7806 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[2,4].Collector
flabel locali 3277 7682 3317 7800 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[2,4].Base
flabel locali 2301 2094 2405 2342 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3,0].Emitter
flabel locali 1730 2153 1779 2254 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3,0].Collector
flabel locali 1889 2130 1929 2248 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3,0].Base
flabel locali 2301 3482 2405 3730 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3,1].Emitter
flabel locali 1730 3541 1779 3642 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3,1].Collector
flabel locali 1889 3518 1929 3636 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3,1].Base
flabel locali 2301 4870 2405 5118 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3,2].Emitter
flabel locali 1730 4929 1779 5030 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3,2].Collector
flabel locali 1889 4906 1929 5024 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3,2].Base
flabel locali 2301 6258 2405 6506 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3,3].Emitter
flabel locali 1730 6317 1779 6418 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3,3].Collector
flabel locali 1889 6294 1929 6412 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3,3].Base
flabel locali 2301 7646 2405 7894 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3,4].Emitter
flabel locali 1730 7705 1779 7806 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3,4].Collector
flabel locali 1889 7682 1929 7800 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3,4].Base
flabel locali 913 2094 1017 2342 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4,0].Emitter
flabel locali 342 2153 391 2254 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4,0].Collector
flabel locali 501 2130 541 2248 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4,0].Base
flabel locali 913 3482 1017 3730 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4,1].Emitter
flabel locali 342 3541 391 3642 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4,1].Collector
flabel locali 501 3518 541 3636 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4,1].Base
flabel locali 913 4870 1017 5118 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4,2].Emitter
flabel locali 342 4929 391 5030 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4,2].Collector
flabel locali 501 4906 541 5024 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4,2].Base
flabel locali 913 6258 1017 6506 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4,3].Emitter
flabel locali 342 6317 391 6418 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4,3].Collector
flabel locali 501 6294 541 6412 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4,3].Base
flabel locali 913 7646 1017 7894 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4,4].Emitter
flabel locali 342 7705 391 7806 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4,4].Collector
flabel locali 501 7682 541 7800 0 FreeSans 400 0 0 0 bjt_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4,4].Base
flabel metal2 1065 12159 1065 12159 0 FreeSans 160 0 0 0 digital_0.S3
flabel metal1 813 12168 813 12168 0 FreeSans 160 0 0 0 digital_0.D3
flabel metal1 1050 12245 1050 12245 0 FreeSans 160 0 0 0 digital_0.trim3
flabel metal2 1947 12161 1947 12161 0 FreeSans 160 0 0 0 digital_0.S2
flabel metal1 1921 12243 1921 12243 0 FreeSans 160 0 0 0 digital_0.trim2
flabel metal1 2810 12248 2810 12248 0 FreeSans 160 0 0 0 digital_0.trim1
flabel metal1 3705 12241 3705 12241 0 FreeSans 160 0 0 0 digital_0.trim0
flabel metal2 2856 12169 2856 12169 0 FreeSans 160 0 0 0 digital_0.S1
flabel metal2 3742 12164 3742 12164 0 FreeSans 160 0 0 0 digital_0.S0
flabel metal1 4669 11294 4669 11294 0 FreeSans 160 0 0 0 digital_0.VENA
flabel metal1 4356 11006 4356 11006 0 FreeSans 160 0 0 0 digital_0.VBGSC
flabel metal1 4356 11622 4356 11622 0 FreeSans 160 0 0 0 digital_0.VBGTC
flabel metal1 4423 10726 4423 10726 0 FreeSans 160 0 0 0 digital_0.SVBGSC
flabel metal1 4424 11842 4424 11842 0 FreeSans 160 0 0 0 digital_0.SVBGTC
flabel metal2 4998 11252 4998 11252 0 FreeSans 160 0 0 0 digital_0.AVDD
flabel metal1 4919 11262 4919 11262 0 FreeSans 160 0 0 0 digital_0.ENA
flabel metal1 5478 10789 5478 10789 0 FreeSans 160 0 0 0 digital_0.VDDE
flabel dnwell 4932 10612 4932 10612 0 FreeSans 160 0 0 0 digital_0.DVDD
flabel pwell 4754 10369 4754 10369 0 FreeSans 160 0 0 0 digital_0.DVSS
flabel metal1 4682 10721 4682 10721 0 FreeSans 160 0 0 0 digital_0.vena_1.G
flabel metal1 4360 10719 4360 10719 0 FreeSans 160 0 0 0 digital_0.vena_1.D
flabel metal1 4608 10725 4608 10725 0 FreeSans 160 0 0 0 digital_0.vena_1.S
flabel psubdiffcont 4419 11163 4419 11163 0 FreeSans 160 0 0 0 digital_0.vena_1.DVSS
flabel metal1 4682 11841 4682 11841 0 FreeSans 160 0 0 0 digital_0.vena_0.G
flabel metal1 4360 11843 4360 11843 0 FreeSans 160 0 0 0 digital_0.vena_0.D
flabel metal1 4608 11837 4608 11837 0 FreeSans 160 0 0 0 digital_0.vena_0.S
flabel psubdiffcont 4419 11399 4419 11399 0 FreeSans 160 0 0 0 digital_0.vena_0.DVSS
flabel metal2 3744 11196 3744 11196 0 FreeSans 160 0 0 0 digital_0.trim_3.S
flabel metal1 3748 12236 3748 12236 0 FreeSans 160 0 0 0 digital_0.trim_3.G
flabel metal1 3483 11361 3483 11361 0 FreeSans 160 0 0 0 digital_0.trim_3.D
flabel psubdiffcont 4195 11278 4195 11278 0 FreeSans 160 0 0 0 digital_0.trim_3.DVSS
flabel metal2 2852 11196 2852 11196 0 FreeSans 160 0 0 0 digital_0.trim_2.S
flabel metal1 2856 12236 2856 12236 0 FreeSans 160 0 0 0 digital_0.trim_2.G
flabel metal1 2591 11361 2591 11361 0 FreeSans 160 0 0 0 digital_0.trim_2.D
flabel psubdiffcont 3303 11278 3303 11278 0 FreeSans 160 0 0 0 digital_0.trim_2.DVSS
flabel metal2 1960 11196 1960 11196 0 FreeSans 160 0 0 0 digital_0.trim_1.S
flabel metal1 1964 12236 1964 12236 0 FreeSans 160 0 0 0 digital_0.trim_1.G
flabel metal1 1699 11361 1699 11361 0 FreeSans 160 0 0 0 digital_0.trim_1.D
flabel psubdiffcont 2411 11278 2411 11278 0 FreeSans 160 0 0 0 digital_0.trim_1.DVSS
flabel metal2 1068 11196 1068 11196 0 FreeSans 160 0 0 0 digital_0.trim_0.S
flabel metal1 1072 12236 1072 12236 0 FreeSans 160 0 0 0 digital_0.trim_0.G
flabel metal1 807 11361 807 11361 0 FreeSans 160 0 0 0 digital_0.trim_0.D
flabel psubdiffcont 1519 11278 1519 11278 0 FreeSans 160 0 0 0 digital_0.trim_0.DVSS
flabel metal1 5477 10790 5477 10790 0 FreeSans 160 0 0 0 digital_0.pmos_ena_0.VDDE
flabel metal2 5578 11244 5578 11244 0 FreeSans 160 0 0 0 digital_0.pmos_ena_0.AVDD
flabel metal1 6051 10924 6051 10924 0 FreeSans 160 0 0 0 digital_0.pmos_ena_0.G
flabel nsubdiffcont 6008 10614 6008 10614 0 FreeSans 160 0 0 0 digital_0.pmos_ena_0.DVDD
flabel metal2 2536 15426 2536 15426 0 FreeSans 160 0 0 0 resistor_op_tt_0.A
flabel metal1 2500 15360 2500 15360 0 FreeSans 160 0 0 0 resistor_op_tt_0.C
flabel metal1 -1089 15365 -1089 15365 0 FreeSans 160 0 0 0 resistor_op_tt_0.B
flabel metal2 -1123 15435 -1123 15435 0 FreeSans 160 0 0 0 resistor_op_tt_0.D
flabel metal1 2556 14863 2556 14863 0 FreeSans 160 0 0 0 resistor_op_tt_0.AVSS
flabel metal1 -3238 15213 -3238 15213 0 FreeSans 1600 0 0 0 pmos_startup_0.D3
flabel metal1 -7360 15238 -7360 15238 0 FreeSans 1600 0 0 0 pmos_startup_0.D2
flabel metal1 -3193 14916 -3193 14916 0 FreeSans 1600 0 0 0 pmos_startup_0.D4
flabel metal1 -5295 14775 -5295 14775 0 FreeSans 1600 0 0 0 pmos_startup_0.VDDE
flabel metal1 -10210 14729 -10210 14729 0 FreeSans 1600 0 0 0 pmos_iptat_0.VDDE
flabel metal1 -8145 15133 -8145 15133 0 FreeSans 1600 0 0 0 pmos_iptat_0.D
flabel metal1 -8678 15483 -8678 15483 0 FreeSans 1600 0 0 0 pmos_iptat_0.G
flabel metal1 8690 15751 8690 15751 0 FreeSans 160 0 0 0 differential_pair_0.AVSS
flabel metal1 5775 14888 5775 14888 0 FreeSans 160 0 0 0 differential_pair_0.S
flabel metal2 6072 15299 6072 15299 0 FreeSans 160 0 0 0 differential_pair_0.PLUS
flabel metal1 6015 15183 6015 15183 0 FreeSans 160 0 0 0 differential_pair_0.MINUS
flabel metal3 8432 15304 8432 15304 0 FreeSans 160 0 0 0 differential_pair_0.D3
flabel metal4 8443 15191 8443 15191 0 FreeSans 160 0 0 0 differential_pair_0.D4
flabel metal1 -5329 17495 -5329 17495 1 FreeSans 160 0 0 0 pmos_current_bgr_2_0.vdde
flabel metal3 -7386 17145 -7386 17145 1 FreeSans 160 0 0 0 pmos_current_bgr_2_0.D3
flabel metal1 -7400 16647 -7400 16647 1 FreeSans 160 0 0 0 pmos_current_bgr_2_0.D9
flabel metal2 -7392 16512 -7392 16512 1 FreeSans 160 0 0 0 pmos_current_bgr_2_0.D8
flabel metal1 -3001 15654 -3001 15654 0 FreeSans 1600 0 0 0 pmos_current_bgr_2_0.VDDE
flabel metal1 -7268 17097 -7268 17097 1 FreeSans 160 0 0 0 pmos_current_bgr_2_0.D4
flabel metal3 -8189 17195 -8189 17195 0 FreeSans 800 0 0 0 pmos_current_bgr_0.D10
flabel metal1 -8186 16732 -8186 16732 0 FreeSans 800 0 0 0 pmos_current_bgr_0.D2
flabel metal2 -12297 16747 -12297 16747 0 FreeSans 800 0 0 0 pmos_current_bgr_0.D1
flabel metal1 -9018 17150 -9018 17150 0 FreeSans 800 0 0 0 pmos_current_bgr_0.G10
flabel metal1 -10241 15714 -10241 15714 0 FreeSans 800 0 0 0 pmos_current_bgr_0.vdde
flabel metal2 76 16706 76 16706 0 FreeSans 160 0 0 0 nmos_tail_current_0.D3
flabel metal3 68 16838 68 16838 0 FreeSans 160 0 0 0 nmos_tail_current_0.D4
flabel metal2 72 17214 72 17214 0 FreeSans 160 0 0 0 nmos_tail_current_0.D1
flabel metal4 4242 16134 4242 16134 0 FreeSans 160 0 0 0 nmos_tail_current_0.S2
flabel metal1 -184 15918 -184 15918 0 FreeSans 160 0 0 0 nmos_tail_current_0.AVSS
flabel metal1 68 16188 68 16188 0 FreeSans 160 0 0 0 nmos_tail_current_0.D2
flabel metal1 -807 17533 -807 17533 0 FreeSans 800 0 0 0 nmos_startup_0.AVSS
flabel metal1 -986 17176 -986 17176 0 FreeSans 800 0 0 0 nmos_startup_0.G1
flabel via1 -544 17206 -544 17206 0 FreeSans 800 0 0 0 nmos_startup_0.D1
flabel metal1 -13008 20464 -13008 20464 0 FreeSans 1600 0 0 0 resistorstart_0.B
flabel metal1 -13007 19641 -13007 19641 0 FreeSans 1600 0 0 0 resistorstart_0.A
flabel metal1 8522 19390 8522 19390 0 FreeSans 1600 0 0 0 resistorstart_0.AVSS
flabel pwell 8699 17764 8699 17764 0 FreeSans 160 0 0 0 res_trim_0.AVSS
flabel metal2 398 19152 398 19152 0 FreeSans 1600 0 0 0 res_trim_0.3
flabel metal3 602 17852 602 17852 0 FreeSans 1600 0 0 0 res_trim_0.2
flabel metal4 726 19154 726 19154 0 FreeSans 1600 0 0 0 res_trim_0.1
flabel metal1 764 17958 764 17958 0 FreeSans 1600 0 0 0 res_trim_0.B
flabel metal4 1358 17814 1358 17814 0 FreeSans 1600 0 0 0 res_trim_0.A
flabel metal1 -17334 21176 -17334 21176 0 FreeSans 800 0 0 0 resist_const_0.B
flabel metal1 -17328 21342 -17328 21342 0 FreeSans 800 0 0 0 resist_const_0.D
flabel metal1 -792 21941 -792 21941 0 FreeSans 800 0 0 0 resist_const_0.VBGSC
flabel metal1 4312 21864 4312 21864 0 FreeSans 800 0 0 0 resist_const_0.VBGTC
flabel metal1 -17327 22172 -17327 22172 0 FreeSans 800 0 0 0 resist_const_0.C
flabel metal1 -17318 22338 -17318 22338 0 FreeSans 800 0 0 0 resist_const_0.A
flabel metal1 -17488 20848 -17488 20848 0 FreeSans 800 0 0 0 resist_const_0.AVSS
flabel metal1 -8658 21724 -8658 21724 0 FreeSans 800 0 0 0 resist_const_0.E
flabel metal1 -143 21872 -143 21872 0 FreeSans 1600 0 0 0 resist_const_0.F
flabel metal4 -9125 7162 -9125 7162 0 FreeSans 1600 0 0 0 cap_op_0.A
flabel metal3 -9780 9016 -9780 9016 0 FreeSans 1600 0 0 0 cap_op_0.B
flabel metal4 -3883 3396 -3883 3396 0 FreeSans 1600 0 0 0 cap_op_0.AVSS
<< end >>
