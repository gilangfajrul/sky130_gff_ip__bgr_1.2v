** sch_path: /foss/designs/sky130_gff_ip__bgr_1.2v/xschem/op_tb-ac.sch
**.subckt op_tb-ac
Vdd v_dd GND 1.8
Vinn v_inn v_ss 0.9
x1 v_out v_dd v_ss v_inp v_inn v_ss v_dd op
Vgnd v_ss GND 0
C1 v_out v_ss 1p m=1
Vinp v_inp v_ss ac 1 sin(0.9 1 1) dc 0.9
**** begin user architecture code
.lib /foss/pdks/sky130A/libs.tech/combined/sky130.lib.spice tt


.temp 27
.option savecurrents
.control
option sparse
save all
op
write op_tb-ac.raw
set appendwrite

ac dec 101 1 100MEG
write op_tb-ac.raw
meas ac phase_margin find vp(v_out) when vdb(v_out)=0
let phase_marginconv = 'phase_margin/pi*180+180'
print phase_marginconv
let phase='vp(v_out)/pi*180+180'
plot vdb(v_out) phase

meas ac dcgain MAX vmag(v_out) FROM=10 TO=10k
let f3db = dcgain/sqrt(2)
meas ac fbw WHEN vmag(v_out)=f3db FALL=1
let gainerror=(dcgain-1)/1
print dcgain
print fbw
print gainerror

noise v(v_out) Vin dec 101 1k 100MEG
print onoise_total

.endc


 .include ./op_tb-ac.save

**** end user architecture code
**.ends

* expanding   symbol:  op.sym # of pins=7
** sym_path: /foss/designs/sky130_gff_ip__bgr_1.2v/xschem/op.sym
** sch_path: /foss/designs/sky130_gff_ip__bgr_1.2v/xschem/op.sch
.subckt op vo_out vdd vss vi_p vi_n psubs nwell
*.iopin vss
*.iopin vdd
*.opin vo_out
*.ipin vi_p
*.ipin vi_n
*.iopin psubs
*.iopin nwell
XM1 net3 vi_n net1 psubs sky130_fd_pr__nfet_01v8 L=5 W=1.35 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
**** begin user architecture code


.include ./sizing_opamp.spice


**** end user architecture code
XM3 net3 net3 vdd nwell sky130_fd_pr__pfet_01v8 L=5 W=1.25 nf=1 ad=0.3625 as=0.3625 pd=3.08 ps=3.08 nrd=0.232 nrs=0.232 sa=0 sb=0
+ sd=0 mult=1 m=1
XM6 net4 net4 vss psubs sky130_fd_pr__nfet_01v8 L=5 W=4 nf=1 ad=1.16 as=1.16 pd=8.58 ps=8.58 nrd=0.0725 nrs=0.0725 sa=0 sb=0 sd=0
+ mult=1 m=1
I0 vdd net4 20e-6
XM5 net1 net4 vss psubs sky130_fd_pr__nfet_01v8 L=5 W=0.75 nf=1 ad=0.2175 as=0.2175 pd=2.08 ps=2.08 nrd=0.386666666666667
+ nrs=0.386666666666667 sa=0 sb=0 sd=0 mult=1 m=1
XM7 vo_out net2 vdd nwell sky130_fd_pr__pfet_01v8 L=5 W=8.5 nf=1 ad=2.465 as=2.465 pd=17.58 ps=17.58 nrd=0.0341176470588235
+ nrs=0.0341176470588235 sa=0 sb=0 sd=0 mult=1 m=1
XM8 vo_out net4 vss psubs sky130_fd_pr__nfet_01v8 L=5 W=0.55 nf=1 ad=0.1595 as=0.1595 pd=1.68 ps=1.68 nrd=0.527272727272727
+ nrs=0.527272727272727 sa=0 sb=0 sd=0 mult=1 m=1
XM2 net2 vi_p net1 psubs sky130_fd_pr__nfet_01v8 L=5 W=1.35 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 net2 net3 vdd nwell sky130_fd_pr__pfet_01v8 L=5 W=1.25 nf=1 ad=0.3625 as=0.3625 pd=3.08 ps=3.08 nrd=0.232 nrs=0.232 sa=0 sb=0
+ sd=0 mult=1 m=1
XR1 net5 net2 vss sky130_fd_pr__res_high_po_0p35 L=10 mult=1 m=1
XC1 vo_out net5 sky130_fd_pr__cap_mim_m3_1 W=128 L=128 MF=1 m=1
.ends

.GLOBAL GND
.end
