magic
tech sky130A
magscale 1 2
timestamp 1716290715
<< nwell >>
rect 524 297 9160 1257
<< pdiff >>
rect 8852 1062 8910 1074
rect 8852 886 8864 1062
rect 8898 886 8910 1062
rect 8852 874 8910 886
<< pdiffc >>
rect 8864 886 8898 1062
<< nsubdiff >>
rect 560 1187 620 1221
rect 9026 1187 9086 1221
rect 560 1161 594 1187
rect 9052 1161 9086 1187
rect 560 367 594 393
rect 9052 367 9086 393
rect 560 333 620 367
rect 9026 333 9086 367
<< nsubdiffcont >>
rect 620 1187 9026 1221
rect 560 393 594 1161
rect 9052 393 9086 1161
rect 620 333 9026 367
<< poly >>
rect 665 1111 736 1154
rect 706 1074 736 1111
rect 8910 1111 8981 1154
rect 8910 1074 8940 1111
rect 1381 807 2207 854
rect 3381 807 4207 854
rect 5439 807 6265 854
rect 7439 807 8265 854
rect 1381 700 2207 747
rect 3381 700 4207 747
rect 5439 700 6265 747
rect 7439 706 8265 747
rect 706 443 736 461
rect 665 400 736 443
rect 8910 443 8940 480
rect 8910 400 8981 443
<< locali >>
rect 560 1187 620 1221
rect 9026 1187 9086 1221
rect 560 1161 594 1187
rect 9052 1161 9086 1187
rect 660 1074 694 1078
rect 8864 1062 8898 1078
rect 8952 1074 8986 1078
rect 8864 870 8898 886
rect 8952 476 8986 480
rect 560 367 594 393
rect 9052 367 9086 393
rect 560 333 620 367
rect 9026 333 9086 367
<< viali >>
rect 4800 1187 4846 1221
rect 560 1112 594 1153
rect 666 1112 735 1153
rect 8911 1112 8980 1153
rect 9052 1112 9086 1153
rect 8864 886 8898 1062
rect 1394 814 2194 848
rect 3394 814 4194 848
rect 5452 814 6252 848
rect 7452 814 8252 848
rect 1394 706 2194 740
rect 3394 706 4194 740
rect 5452 706 6252 740
rect 7452 706 8252 740
rect 560 401 594 442
rect 666 401 735 442
rect 8911 401 8980 442
rect 9052 401 9086 442
rect 4798 333 4844 367
<< metal1 >>
rect 4788 1221 4858 1227
rect 4788 1187 4800 1221
rect 4846 1187 4858 1221
rect 4788 1181 4858 1187
rect 554 1153 600 1165
rect 654 1153 747 1165
rect 554 1112 560 1153
rect 594 1112 666 1153
rect 735 1112 747 1153
rect 554 1100 600 1112
rect 654 1106 747 1112
rect 654 1074 700 1106
rect 4800 1070 4846 1181
rect 8899 1153 8992 1165
rect 9046 1153 9092 1165
rect 8899 1112 8911 1153
rect 8980 1112 9052 1153
rect 9086 1112 9092 1153
rect 8899 1106 8992 1112
rect 8946 1074 8992 1106
rect 9046 1100 9092 1112
rect 8858 1062 8904 1074
rect 742 808 788 882
rect 1382 848 2206 854
rect 1382 814 1394 848
rect 2194 814 2206 848
rect 1382 809 2206 814
rect 3382 848 4206 854
rect 3382 814 3394 848
rect 4194 814 4206 848
rect 1382 808 2207 809
rect 3382 808 4206 814
rect 742 807 4206 808
rect 742 747 4094 807
rect 4194 747 4206 807
rect 742 746 4206 747
rect 1382 740 2206 746
rect 1382 706 1394 740
rect 2194 706 2206 740
rect 1382 700 2206 706
rect 3382 740 4206 746
rect 3382 706 3394 740
rect 4194 706 4206 740
rect 3382 700 4206 706
rect 4798 672 4844 906
rect 8845 886 8855 1062
rect 8907 886 8917 1062
rect 8858 874 8904 886
rect 5440 848 6264 854
rect 5440 814 5452 848
rect 6252 814 6264 848
rect 5440 808 6264 814
rect 7440 848 8264 854
rect 7440 814 7452 848
rect 8252 814 8264 848
rect 7440 808 8264 814
rect 5440 807 8904 808
rect 5440 747 5452 807
rect 5552 747 8904 807
rect 5440 746 8904 747
rect 5440 740 6264 746
rect 5440 706 5452 740
rect 6252 706 6264 740
rect 5440 700 6264 706
rect 7440 740 8264 746
rect 7440 706 7452 740
rect 8252 706 8264 740
rect 7440 700 8264 706
rect 8858 676 8904 746
rect 729 492 739 668
rect 791 492 801 668
rect 554 442 600 454
rect 654 448 700 485
rect 654 442 747 448
rect 554 401 560 442
rect 594 401 666 442
rect 735 401 747 442
rect 554 389 600 401
rect 654 389 747 401
rect 4798 373 4844 480
rect 8946 448 8992 480
rect 8899 442 8992 448
rect 9046 442 9092 454
rect 8899 401 8911 442
rect 8980 401 9052 442
rect 9086 401 9092 442
rect 8899 389 8992 401
rect 9046 389 9092 401
rect 4786 367 4856 373
rect 4786 333 4798 367
rect 4844 333 4856 367
rect 4786 327 4856 333
<< via1 >>
rect 4094 747 4194 807
rect 8855 886 8864 1062
rect 8864 886 8898 1062
rect 8898 886 8907 1062
rect 5452 747 5552 807
rect 739 492 791 668
<< metal2 >>
rect 8855 1062 8907 1072
rect 8855 828 8907 886
rect 710 812 819 822
rect 8826 818 8935 828
rect 4094 807 4194 817
rect 5452 807 5552 817
rect 4194 747 5452 807
rect 4094 737 4194 747
rect 5452 737 5552 747
rect 710 726 819 736
rect 8826 732 8935 742
rect 739 668 791 726
rect 739 482 791 492
<< via2 >>
rect 710 736 819 812
rect 8826 742 8935 818
<< metal3 >>
rect 8816 818 8945 823
rect 8816 817 8826 818
rect 700 812 8826 817
rect 700 736 710 812
rect 819 742 8826 812
rect 8935 742 8945 818
rect 819 737 8945 742
rect 819 736 829 737
rect 700 731 829 736
use sky130_fd_pr__pfet_01v8_2XU96L  sky130_fd_pr__pfet_01v8_2XU96L_0 ~/chipalooza/sky130_gff_ip__bgr_1.2v/magic
timestamp 1716189928
transform 1 0 8925 0 1 580
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XU96L  sky130_fd_pr__pfet_01v8_2XU96L_1
timestamp 1716189928
transform 1 0 721 0 1 580
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XU96L  sky130_fd_pr__pfet_01v8_2XU96L_2
timestamp 1716189928
transform 1 0 721 0 1 974
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XU96L  sky130_fd_pr__pfet_01v8_2XU96L_3
timestamp 1716189928
transform 1 0 8925 0 1 974
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_H288V5  sky130_fd_pr__pfet_01v8_H288V5_0
timestamp 1716133296
transform 1 0 4823 0 1 974
box -4123 -162 4123 162
use sky130_fd_pr__pfet_01v8_H288V5  sky130_fd_pr__pfet_01v8_H288V5_1
timestamp 1716133296
transform 1 0 4823 0 1 580
box -4123 -162 4123 162
<< end >>
