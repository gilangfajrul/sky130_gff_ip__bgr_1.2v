magic
tech sky130A
magscale 1 2
timestamp 1716353109
<< nmos >>
rect -15 -70 15 70
<< ndiff >>
rect -73 58 -15 70
rect -73 -58 -61 58
rect -27 -58 -15 58
rect -73 -70 -15 -58
rect 15 58 73 70
rect 15 -58 27 58
rect 61 -58 73 58
rect 15 -70 73 -58
<< ndiffc >>
rect -61 -58 -27 58
rect 27 -58 61 58
<< poly >>
rect -15 70 15 96
rect -15 -96 15 -70
<< locali >>
rect -61 58 -27 74
rect -61 -74 -27 -58
rect 27 58 61 74
rect 27 -74 61 -58
<< viali >>
rect -61 -58 -27 58
rect 27 -58 61 58
<< metal1 >>
rect -67 58 -21 70
rect -67 -58 -61 58
rect -27 -58 -21 58
rect -67 -70 -21 -58
rect 21 58 67 70
rect 21 -58 27 58
rect 61 -58 67 58
rect 21 -70 67 -58
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.7 l 0.150 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
