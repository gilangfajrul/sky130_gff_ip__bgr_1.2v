magic
tech sky130A
magscale 1 2
timestamp 1716392830
<< nwell >>
rect -677 -3995 677 3995
<< nsubdiff >>
rect -641 3925 -545 3959
rect 545 3925 641 3959
rect -641 3863 -607 3925
rect 607 3863 641 3925
rect -641 -3925 -607 -3863
rect 607 -3925 641 -3863
rect -641 -3959 -545 -3925
rect 545 -3959 641 -3925
<< nsubdiffcont >>
rect -545 3925 545 3959
rect -641 -3863 -607 3863
rect 607 -3863 641 3863
rect -545 -3959 545 -3925
<< xpolycontact >>
rect -450 3388 -380 3820
rect -450 1988 -380 2420
rect -284 3388 -214 3820
rect -284 1988 -214 2420
rect -118 3388 -48 3820
rect -118 1988 -48 2420
rect 48 3388 118 3820
rect 48 1988 118 2420
rect 214 3388 284 3820
rect 214 1988 284 2420
rect 380 3388 450 3820
rect 380 1988 450 2420
rect -450 1452 -380 1884
rect -450 52 -380 484
rect -284 1452 -214 1884
rect -284 52 -214 484
rect -118 1452 -48 1884
rect -118 52 -48 484
rect 48 1452 118 1884
rect 48 52 118 484
rect 214 1452 284 1884
rect 214 52 284 484
rect 380 1452 450 1884
rect 380 52 450 484
rect -450 -484 -380 -52
rect -450 -1884 -380 -1452
rect -284 -484 -214 -52
rect -284 -1884 -214 -1452
rect -118 -484 -48 -52
rect -118 -1884 -48 -1452
rect 48 -484 118 -52
rect 48 -1884 118 -1452
rect 214 -484 284 -52
rect 214 -1884 284 -1452
rect 380 -484 450 -52
rect 380 -1884 450 -1452
rect -450 -2420 -380 -1988
rect -450 -3820 -380 -3388
rect -284 -2420 -214 -1988
rect -284 -3820 -214 -3388
rect -118 -2420 -48 -1988
rect -118 -3820 -48 -3388
rect 48 -2420 118 -1988
rect 48 -3820 118 -3388
rect 214 -2420 284 -1988
rect 214 -3820 284 -3388
rect 380 -2420 450 -1988
rect 380 -3820 450 -3388
<< ppolyres >>
rect -450 2420 -380 3388
rect -284 2420 -214 3388
rect -118 2420 -48 3388
rect 48 2420 118 3388
rect 214 2420 284 3388
rect 380 2420 450 3388
rect -450 484 -380 1452
rect -284 484 -214 1452
rect -118 484 -48 1452
rect 48 484 118 1452
rect 214 484 284 1452
rect 380 484 450 1452
rect -450 -1452 -380 -484
rect -284 -1452 -214 -484
rect -118 -1452 -48 -484
rect 48 -1452 118 -484
rect 214 -1452 284 -484
rect 380 -1452 450 -484
rect -450 -3388 -380 -2420
rect -284 -3388 -214 -2420
rect -118 -3388 -48 -2420
rect 48 -3388 118 -2420
rect 214 -3388 284 -2420
rect 380 -3388 450 -2420
<< locali >>
rect -641 3925 -545 3959
rect 545 3925 641 3959
rect -641 3863 -607 3925
rect 607 3863 641 3925
rect -641 -3925 -607 -3863
rect 607 -3925 641 -3863
rect -641 -3959 -545 -3925
rect 545 -3959 641 -3925
<< viali >>
rect -434 3405 -396 3802
rect -268 3405 -230 3802
rect -102 3405 -64 3802
rect 64 3405 102 3802
rect 230 3405 268 3802
rect 396 3405 434 3802
rect -434 2006 -396 2403
rect -268 2006 -230 2403
rect -102 2006 -64 2403
rect 64 2006 102 2403
rect 230 2006 268 2403
rect 396 2006 434 2403
rect -434 1469 -396 1866
rect -268 1469 -230 1866
rect -102 1469 -64 1866
rect 64 1469 102 1866
rect 230 1469 268 1866
rect 396 1469 434 1866
rect -434 70 -396 467
rect -268 70 -230 467
rect -102 70 -64 467
rect 64 70 102 467
rect 230 70 268 467
rect 396 70 434 467
rect -434 -467 -396 -70
rect -268 -467 -230 -70
rect -102 -467 -64 -70
rect 64 -467 102 -70
rect 230 -467 268 -70
rect 396 -467 434 -70
rect -434 -1866 -396 -1469
rect -268 -1866 -230 -1469
rect -102 -1866 -64 -1469
rect 64 -1866 102 -1469
rect 230 -1866 268 -1469
rect 396 -1866 434 -1469
rect -434 -2403 -396 -2006
rect -268 -2403 -230 -2006
rect -102 -2403 -64 -2006
rect 64 -2403 102 -2006
rect 230 -2403 268 -2006
rect 396 -2403 434 -2006
rect -434 -3802 -396 -3405
rect -268 -3802 -230 -3405
rect -102 -3802 -64 -3405
rect 64 -3802 102 -3405
rect 230 -3802 268 -3405
rect 396 -3802 434 -3405
<< metal1 >>
rect -440 3802 -390 3814
rect -440 3405 -434 3802
rect -396 3405 -390 3802
rect -440 3393 -390 3405
rect -274 3802 -224 3814
rect -274 3405 -268 3802
rect -230 3405 -224 3802
rect -274 3393 -224 3405
rect -108 3802 -58 3814
rect -108 3405 -102 3802
rect -64 3405 -58 3802
rect -108 3393 -58 3405
rect 58 3802 108 3814
rect 58 3405 64 3802
rect 102 3405 108 3802
rect 58 3393 108 3405
rect 224 3802 274 3814
rect 224 3405 230 3802
rect 268 3405 274 3802
rect 224 3393 274 3405
rect 390 3802 440 3814
rect 390 3405 396 3802
rect 434 3405 440 3802
rect 390 3393 440 3405
rect -440 2403 -390 2415
rect -440 2006 -434 2403
rect -396 2006 -390 2403
rect -440 1994 -390 2006
rect -274 2403 -224 2415
rect -274 2006 -268 2403
rect -230 2006 -224 2403
rect -274 1994 -224 2006
rect -108 2403 -58 2415
rect -108 2006 -102 2403
rect -64 2006 -58 2403
rect -108 1994 -58 2006
rect 58 2403 108 2415
rect 58 2006 64 2403
rect 102 2006 108 2403
rect 58 1994 108 2006
rect 224 2403 274 2415
rect 224 2006 230 2403
rect 268 2006 274 2403
rect 224 1994 274 2006
rect 390 2403 440 2415
rect 390 2006 396 2403
rect 434 2006 440 2403
rect 390 1994 440 2006
rect -440 1866 -390 1878
rect -440 1469 -434 1866
rect -396 1469 -390 1866
rect -440 1457 -390 1469
rect -274 1866 -224 1878
rect -274 1469 -268 1866
rect -230 1469 -224 1866
rect -274 1457 -224 1469
rect -108 1866 -58 1878
rect -108 1469 -102 1866
rect -64 1469 -58 1866
rect -108 1457 -58 1469
rect 58 1866 108 1878
rect 58 1469 64 1866
rect 102 1469 108 1866
rect 58 1457 108 1469
rect 224 1866 274 1878
rect 224 1469 230 1866
rect 268 1469 274 1866
rect 224 1457 274 1469
rect 390 1866 440 1878
rect 390 1469 396 1866
rect 434 1469 440 1866
rect 390 1457 440 1469
rect -440 467 -390 479
rect -440 70 -434 467
rect -396 70 -390 467
rect -440 58 -390 70
rect -274 467 -224 479
rect -274 70 -268 467
rect -230 70 -224 467
rect -274 58 -224 70
rect -108 467 -58 479
rect -108 70 -102 467
rect -64 70 -58 467
rect -108 58 -58 70
rect 58 467 108 479
rect 58 70 64 467
rect 102 70 108 467
rect 58 58 108 70
rect 224 467 274 479
rect 224 70 230 467
rect 268 70 274 467
rect 224 58 274 70
rect 390 467 440 479
rect 390 70 396 467
rect 434 70 440 467
rect 390 58 440 70
rect -440 -70 -390 -58
rect -440 -467 -434 -70
rect -396 -467 -390 -70
rect -440 -479 -390 -467
rect -274 -70 -224 -58
rect -274 -467 -268 -70
rect -230 -467 -224 -70
rect -274 -479 -224 -467
rect -108 -70 -58 -58
rect -108 -467 -102 -70
rect -64 -467 -58 -70
rect -108 -479 -58 -467
rect 58 -70 108 -58
rect 58 -467 64 -70
rect 102 -467 108 -70
rect 58 -479 108 -467
rect 224 -70 274 -58
rect 224 -467 230 -70
rect 268 -467 274 -70
rect 224 -479 274 -467
rect 390 -70 440 -58
rect 390 -467 396 -70
rect 434 -467 440 -70
rect 390 -479 440 -467
rect -440 -1469 -390 -1457
rect -440 -1866 -434 -1469
rect -396 -1866 -390 -1469
rect -440 -1878 -390 -1866
rect -274 -1469 -224 -1457
rect -274 -1866 -268 -1469
rect -230 -1866 -224 -1469
rect -274 -1878 -224 -1866
rect -108 -1469 -58 -1457
rect -108 -1866 -102 -1469
rect -64 -1866 -58 -1469
rect -108 -1878 -58 -1866
rect 58 -1469 108 -1457
rect 58 -1866 64 -1469
rect 102 -1866 108 -1469
rect 58 -1878 108 -1866
rect 224 -1469 274 -1457
rect 224 -1866 230 -1469
rect 268 -1866 274 -1469
rect 224 -1878 274 -1866
rect 390 -1469 440 -1457
rect 390 -1866 396 -1469
rect 434 -1866 440 -1469
rect 390 -1878 440 -1866
rect -440 -2006 -390 -1994
rect -440 -2403 -434 -2006
rect -396 -2403 -390 -2006
rect -440 -2415 -390 -2403
rect -274 -2006 -224 -1994
rect -274 -2403 -268 -2006
rect -230 -2403 -224 -2006
rect -274 -2415 -224 -2403
rect -108 -2006 -58 -1994
rect -108 -2403 -102 -2006
rect -64 -2403 -58 -2006
rect -108 -2415 -58 -2403
rect 58 -2006 108 -1994
rect 58 -2403 64 -2006
rect 102 -2403 108 -2006
rect 58 -2415 108 -2403
rect 224 -2006 274 -1994
rect 224 -2403 230 -2006
rect 268 -2403 274 -2006
rect 224 -2415 274 -2403
rect 390 -2006 440 -1994
rect 390 -2403 396 -2006
rect 434 -2403 440 -2006
rect 390 -2415 440 -2403
rect -440 -3405 -390 -3393
rect -440 -3802 -434 -3405
rect -396 -3802 -390 -3405
rect -440 -3814 -390 -3802
rect -274 -3405 -224 -3393
rect -274 -3802 -268 -3405
rect -230 -3802 -224 -3405
rect -274 -3814 -224 -3802
rect -108 -3405 -58 -3393
rect -108 -3802 -102 -3405
rect -64 -3802 -58 -3405
rect -108 -3814 -58 -3802
rect 58 -3405 108 -3393
rect 58 -3802 64 -3405
rect 102 -3802 108 -3405
rect 58 -3814 108 -3802
rect 224 -3405 274 -3393
rect 224 -3802 230 -3405
rect 268 -3802 274 -3405
rect 224 -3814 274 -3802
rect 390 -3405 440 -3393
rect 390 -3802 396 -3405
rect 434 -3802 440 -3405
rect 390 -3814 440 -3802
<< properties >>
string FIXED_BBOX -624 -3942 624 3942
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.350 l 5 m 4 nx 6 wmin 0.350 lmin 0.50 rho 319.8 val 5.681k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.350 vias 1 n_guard 1 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
