magic
tech sky130A
magscale 1 2
timestamp 1720030824
<< xpolycontact >>
rect -450 1252 -380 1684
rect -450 52 -380 484
rect -284 1252 -214 1684
rect -284 52 -214 484
rect -118 1252 -48 1684
rect -118 52 -48 484
rect 48 1252 118 1684
rect 48 52 118 484
rect 214 1252 284 1684
rect 214 52 284 484
rect 380 1252 450 1684
rect 380 52 450 484
rect -450 -484 -380 -52
rect -450 -1684 -380 -1252
rect -284 -484 -214 -52
rect -284 -1684 -214 -1252
rect -118 -484 -48 -52
rect -118 -1684 -48 -1252
rect 48 -484 118 -52
rect 48 -1684 118 -1252
rect 214 -484 284 -52
rect 214 -1684 284 -1252
rect 380 -484 450 -52
rect 380 -1684 450 -1252
<< ppolyres >>
rect -450 484 -380 1252
rect -284 484 -214 1252
rect -118 484 -48 1252
rect 48 484 118 1252
rect 214 484 284 1252
rect 380 484 450 1252
rect -450 -1252 -380 -484
rect -284 -1252 -214 -484
rect -118 -1252 -48 -484
rect 48 -1252 118 -484
rect 214 -1252 284 -484
rect 380 -1252 450 -484
<< viali >>
rect -434 1269 -396 1666
rect -268 1269 -230 1666
rect -102 1269 -64 1666
rect 64 1269 102 1666
rect 230 1269 268 1666
rect 396 1269 434 1666
rect -434 70 -396 467
rect -268 70 -230 467
rect -102 70 -64 467
rect 64 70 102 467
rect 230 70 268 467
rect 396 70 434 467
rect -434 -467 -396 -70
rect -268 -467 -230 -70
rect -102 -467 -64 -70
rect 64 -467 102 -70
rect 230 -467 268 -70
rect 396 -467 434 -70
rect -434 -1666 -396 -1269
rect -268 -1666 -230 -1269
rect -102 -1666 -64 -1269
rect 64 -1666 102 -1269
rect 230 -1666 268 -1269
rect 396 -1666 434 -1269
<< metal1 >>
rect -440 1666 -390 1678
rect -440 1269 -434 1666
rect -396 1269 -390 1666
rect -440 1257 -390 1269
rect -274 1666 -224 1678
rect -274 1269 -268 1666
rect -230 1269 -224 1666
rect -274 1257 -224 1269
rect -108 1666 -58 1678
rect -108 1269 -102 1666
rect -64 1269 -58 1666
rect -108 1257 -58 1269
rect 58 1666 108 1678
rect 58 1269 64 1666
rect 102 1269 108 1666
rect 58 1257 108 1269
rect 224 1666 274 1678
rect 224 1269 230 1666
rect 268 1269 274 1666
rect 224 1257 274 1269
rect 390 1666 440 1678
rect 390 1269 396 1666
rect 434 1269 440 1666
rect 390 1257 440 1269
rect -440 467 -390 479
rect -440 70 -434 467
rect -396 70 -390 467
rect -440 58 -390 70
rect -274 467 -224 479
rect -274 70 -268 467
rect -230 70 -224 467
rect -274 58 -224 70
rect -108 467 -58 479
rect -108 70 -102 467
rect -64 70 -58 467
rect -108 58 -58 70
rect 58 467 108 479
rect 58 70 64 467
rect 102 70 108 467
rect 58 58 108 70
rect 224 467 274 479
rect 224 70 230 467
rect 268 70 274 467
rect 224 58 274 70
rect 390 467 440 479
rect 390 70 396 467
rect 434 70 440 467
rect 390 58 440 70
rect -440 -70 -390 -58
rect -440 -467 -434 -70
rect -396 -467 -390 -70
rect -440 -479 -390 -467
rect -274 -70 -224 -58
rect -274 -467 -268 -70
rect -230 -467 -224 -70
rect -274 -479 -224 -467
rect -108 -70 -58 -58
rect -108 -467 -102 -70
rect -64 -467 -58 -70
rect -108 -479 -58 -467
rect 58 -70 108 -58
rect 58 -467 64 -70
rect 102 -467 108 -70
rect 58 -479 108 -467
rect 224 -70 274 -58
rect 224 -467 230 -70
rect 268 -467 274 -70
rect 224 -479 274 -467
rect 390 -70 440 -58
rect 390 -467 396 -70
rect 434 -467 440 -70
rect 390 -479 440 -467
rect -440 -1269 -390 -1257
rect -440 -1666 -434 -1269
rect -396 -1666 -390 -1269
rect -440 -1678 -390 -1666
rect -274 -1269 -224 -1257
rect -274 -1666 -268 -1269
rect -230 -1666 -224 -1269
rect -274 -1678 -224 -1666
rect -108 -1269 -58 -1257
rect -108 -1666 -102 -1269
rect -64 -1666 -58 -1269
rect -108 -1678 -58 -1666
rect 58 -1269 108 -1257
rect 58 -1666 64 -1269
rect 102 -1666 108 -1269
rect 58 -1678 108 -1666
rect 224 -1269 274 -1257
rect 224 -1666 230 -1269
rect 268 -1666 274 -1269
rect 224 -1678 274 -1666
rect 390 -1269 440 -1257
rect 390 -1666 396 -1269
rect 434 -1666 440 -1269
rect 390 -1678 440 -1666
<< properties >>
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.350 l 4 m 2 nx 6 wmin 0.350 lmin 0.50 rho 319.8 val 4.768k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
