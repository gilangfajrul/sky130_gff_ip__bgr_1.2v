magic
tech sky130A
magscale 1 2
timestamp 1717432846
<< psubdiff >>
rect -561 824 -501 858
rect 3935 824 3995 858
rect -561 798 -527 824
rect 3961 798 3995 824
rect -561 -55 -527 -29
rect 3961 -55 3995 -29
rect -561 -89 -501 -55
rect 3935 -89 3995 -55
<< psubdiffcont >>
rect -501 824 3935 858
rect -561 -29 -527 798
rect 3961 -29 3995 798
rect -501 -89 3935 -55
<< poly >>
rect -400 375 -370 454
rect -462 359 -370 375
rect -462 325 -446 359
rect -412 325 -370 359
rect -462 309 -370 325
rect -400 228 -370 309
rect 3804 375 3834 453
rect 3804 359 3896 375
rect 3804 325 3846 359
rect 3880 325 3896 359
rect 3804 309 3896 325
rect 3804 238 3834 309
<< polycont >>
rect -446 325 -412 359
rect 3846 325 3880 359
<< locali >>
rect -561 824 -501 858
rect 3935 824 3995 858
rect -561 798 -527 824
rect 3961 798 3995 824
rect -446 359 -412 375
rect -446 309 -412 325
rect 3846 359 3880 375
rect 3846 309 3880 325
rect -561 -55 -527 -29
rect 3961 -55 3995 -29
rect -561 -89 -501 -55
rect 3935 -89 3995 -55
<< viali >>
rect -561 325 -527 359
rect -446 325 -412 359
rect 3846 325 3880 359
rect 3961 325 3995 359
<< metal1 >>
rect -520 747 -510 799
rect -458 796 -448 799
rect 3882 796 3892 799
rect -458 750 3892 796
rect -458 747 -448 750
rect 1694 616 1740 750
rect 3882 747 3892 750
rect 3944 747 3954 799
rect -452 371 -406 485
rect -377 480 -367 616
rect -315 480 -305 616
rect 3739 480 3749 616
rect 3801 480 3811 616
rect 1192 390 1578 436
rect -567 359 -406 371
rect -567 325 -561 359
rect -527 325 -446 359
rect -412 325 -406 359
rect -567 313 -406 325
rect 1532 365 1578 390
rect 2244 387 2254 439
rect 3238 387 3248 439
rect 3840 371 3886 475
rect 1532 319 1902 365
rect -452 213 -406 313
rect 186 245 196 297
rect 1180 245 1190 297
rect 1856 294 1902 319
rect 3840 359 4001 371
rect 3840 325 3846 359
rect 3880 325 3961 359
rect 3995 325 4001 359
rect 3840 313 4001 325
rect 1856 248 2242 294
rect 3840 211 3886 313
rect -377 68 -367 204
rect -315 68 -305 204
rect 3739 68 3749 204
rect 3801 68 3811 204
rect -520 -43 -510 9
rect -458 6 -448 9
rect 1694 6 1740 56
rect 3882 6 3892 9
rect -458 -40 3892 6
rect -458 -43 -448 -40
rect 3882 -43 3892 -40
rect 3944 -43 3954 9
<< via1 >>
rect -510 747 -458 799
rect 3892 747 3944 799
rect -367 480 -315 616
rect 3749 480 3801 616
rect 2254 387 3238 439
rect 196 245 1180 297
rect -367 68 -315 204
rect 3749 68 3801 204
rect -510 -43 -458 9
rect 3892 -43 3944 9
<< metal2 >>
rect -510 799 -458 809
rect -510 9 -458 747
rect 3892 799 3944 809
rect -369 616 -313 626
rect -369 470 -313 480
rect 3747 616 3803 626
rect 3747 470 3803 480
rect 2254 439 3238 449
rect 1850 387 2254 439
rect 1850 368 1902 387
rect 2254 377 3238 387
rect 1532 316 1902 368
rect 196 297 1180 307
rect 1532 297 1584 316
rect 1180 245 1584 297
rect 196 235 1180 245
rect -369 204 -313 214
rect -369 58 -313 68
rect 3747 204 3803 214
rect 3747 58 3803 68
rect -510 -53 -458 -43
rect 3892 9 3944 747
rect 3892 -53 3944 -43
<< via2 >>
rect -369 480 -367 616
rect -367 480 -315 616
rect -315 480 -313 616
rect 3747 480 3749 616
rect 3749 480 3801 616
rect 3801 480 3803 616
rect -369 68 -367 204
rect -367 68 -315 204
rect -315 68 -313 204
rect 3747 68 3749 204
rect 3749 68 3801 204
rect 3801 68 3803 204
<< metal3 >>
rect -379 616 -303 621
rect 3737 616 3813 621
rect -379 480 -369 616
rect -313 480 -303 616
rect 3733 480 3743 616
rect 3807 480 3817 616
rect -379 475 -303 480
rect 3737 475 3813 480
rect -371 372 -311 475
rect -371 312 3805 372
rect 3745 209 3805 312
rect -379 204 -303 209
rect 3737 204 3813 209
rect -383 68 -373 204
rect -309 68 -299 204
rect 3737 68 3747 204
rect 3803 68 3813 204
rect -379 63 -303 68
rect 3737 63 3813 68
<< via3 >>
rect 3743 480 3747 616
rect 3747 480 3803 616
rect 3803 480 3807 616
rect -373 68 -369 204
rect -369 68 -313 204
rect -313 68 -309 204
<< metal4 >>
rect 3742 616 3808 617
rect 3742 480 3743 616
rect 3807 480 3808 616
rect 3742 479 3808 480
rect 3745 372 3805 479
rect -371 312 3805 372
rect -371 205 -311 312
rect -374 204 -308 205
rect -374 68 -373 204
rect -309 68 -308 204
rect -374 67 -308 68
use sky130_fd_pr__nfet_01v8_4VSDG9  sky130_fd_pr__nfet_01v8_4VSDG9_0
timestamp 1717432527
transform 1 0 3819 0 1 548
box -73 -106 73 106
use sky130_fd_pr__nfet_01v8_4VSDG9  sky130_fd_pr__nfet_01v8_4VSDG9_1
timestamp 1717432527
transform 1 0 -385 0 1 548
box -73 -106 73 106
use sky130_fd_pr__nfet_01v8_4VSDG9  sky130_fd_pr__nfet_01v8_4VSDG9_2
timestamp 1717432527
transform 1 0 -385 0 1 136
box -73 -106 73 106
use sky130_fd_pr__nfet_01v8_4VSDG9  sky130_fd_pr__nfet_01v8_4VSDG9_4
timestamp 1717432527
transform 1 0 3819 0 1 136
box -73 -106 73 106
use sky130_fd_pr__nfet_01v8_BAH34H  sky130_fd_pr__nfet_01v8_BAH34H_0
timestamp 1717432527
transform 1 0 1717 0 -1 548
box -2087 -168 2087 168
use sky130_fd_pr__nfet_01v8_N7TR4F  sky130_fd_pr__nfet_01v8_N7TR4F_1
timestamp 1717428712
transform 1 0 1717 0 1 167
box -2087 -137 2087 137
<< labels >>
flabel metal4 3774 404 3774 404 0 FreeSans 160 0 0 0 D4
port 0 nsew
flabel metal3 3771 267 3771 267 0 FreeSans 160 0 0 0 D3
port 1 nsew
flabel metal1 3872 406 3872 406 0 FreeSans 160 0 0 0 AVSS
port 2 nsew
flabel metal2 3923 426 3923 426 0 FreeSans 160 0 0 0 S
port 3 nsew
flabel metal1 1876 291 1876 291 0 FreeSans 160 0 0 0 plus
port 4 nsew
flabel metal2 1873 388 1873 388 0 FreeSans 160 0 0 0 minus
port 5 nsew
<< end >>
