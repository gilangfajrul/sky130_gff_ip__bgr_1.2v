magic
tech sky130A
magscale 1 2
timestamp 1720116957
<< nmos >>
rect -2629 -90 -29 90
rect 29 -90 2629 90
<< ndiff >>
rect -2687 78 -2629 90
rect -2687 -78 -2675 78
rect -2641 -78 -2629 78
rect -2687 -90 -2629 -78
rect -29 78 29 90
rect -29 -78 -17 78
rect 17 -78 29 78
rect -29 -90 29 -78
rect 2629 78 2687 90
rect 2629 -78 2641 78
rect 2675 -78 2687 78
rect 2629 -90 2687 -78
<< ndiffc >>
rect -2675 -78 -2641 78
rect -17 -78 17 78
rect 2641 -78 2675 78
<< poly >>
rect -1987 162 -671 178
rect -1987 145 -1971 162
rect -2629 128 -1971 145
rect -687 145 -671 162
rect 671 162 1987 178
rect 671 145 687 162
rect -687 128 -29 145
rect -2629 90 -29 128
rect 29 128 687 145
rect 1971 145 1987 162
rect 1971 128 2629 145
rect 29 90 2629 128
rect -2629 -128 -29 -90
rect -2629 -145 -1971 -128
rect -1987 -162 -1971 -145
rect -687 -145 -29 -128
rect 29 -128 2629 -90
rect 29 -145 687 -128
rect -687 -162 -671 -145
rect -1987 -178 -671 -162
rect 671 -162 687 -145
rect 1971 -145 2629 -128
rect 1971 -162 1987 -145
rect 671 -178 1987 -162
<< polycont >>
rect -1971 128 -687 162
rect 687 128 1971 162
rect -1971 -162 -687 -128
rect 687 -162 1971 -128
<< locali >>
rect -1987 128 -1971 162
rect -687 128 -671 162
rect 671 128 687 162
rect 1971 128 1987 162
rect -2675 78 -2641 94
rect -2675 -94 -2641 -78
rect -17 78 17 94
rect -17 -94 17 -78
rect 2641 78 2675 94
rect 2641 -94 2675 -78
rect -1987 -162 -1971 -128
rect -687 -162 -671 -128
rect 671 -162 687 -128
rect 1971 -162 1987 -128
<< viali >>
rect -1971 128 -687 162
rect 687 128 1971 162
rect -2675 -78 -2641 78
rect -17 -78 17 78
rect 2641 -78 2675 78
rect -1971 -162 -687 -128
rect 687 -162 1971 -128
<< metal1 >>
rect -1983 162 -675 168
rect -1983 128 -1971 162
rect -687 128 -675 162
rect -1983 122 -675 128
rect 675 162 1983 168
rect 675 128 687 162
rect 1971 128 1983 162
rect 675 122 1983 128
rect -2681 78 -2635 90
rect -2681 -78 -2675 78
rect -2641 -78 -2635 78
rect -2681 -90 -2635 -78
rect -23 78 23 90
rect -23 -78 -17 78
rect 17 -78 23 78
rect -23 -90 23 -78
rect 2635 78 2681 90
rect 2635 -78 2641 78
rect 2675 -78 2681 78
rect 2635 -90 2681 -78
rect -1983 -128 -675 -122
rect -1983 -162 -1971 -128
rect -687 -162 -675 -128
rect -1983 -168 -675 -162
rect 675 -128 1983 -122
rect 675 -162 687 -128
rect 1971 -162 1983 -128
rect 675 -168 1983 -162
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.9 l 13 m 1 nf 2 diffcov 100 polycov 50 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
