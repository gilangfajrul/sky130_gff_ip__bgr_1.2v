magic
tech sky130A
magscale 1 2
timestamp 1717511434
<< checkpaint >>
rect 5002 -9752 7944 -9434
rect 5002 -13364 10138 -9752
rect 7196 -13682 10138 -13364
<< error_s >>
rect 298 -241 333 -207
rect 299 -260 333 -241
rect 200 -390 207 -372
rect 129 -521 187 -515
rect 129 -555 141 -521
rect 129 -561 187 -555
rect 129 -841 187 -835
rect 129 -875 141 -841
rect 129 -881 187 -875
rect 129 -949 187 -943
rect 129 -972 141 -949
rect 129 -989 187 -972
rect 101 -1017 200 -1000
rect 129 -1269 187 -1263
rect 129 -1303 141 -1269
rect 129 -1309 187 -1303
rect 318 -1617 333 -260
rect 352 -294 387 -260
rect 352 -1617 386 -294
rect 498 -362 556 -356
rect 498 -396 510 -362
rect 498 -402 556 -396
rect 1236 -468 1294 -462
rect 1236 -502 1248 -468
rect 1236 -508 1294 -502
rect 498 -574 556 -568
rect 498 -608 510 -574
rect 498 -614 556 -608
rect 498 -682 556 -676
rect 1236 -680 1294 -674
rect 498 -716 510 -682
rect 1236 -714 1248 -680
rect 498 -722 556 -716
rect 1236 -720 1294 -714
rect 1236 -788 1294 -782
rect 1236 -822 1248 -788
rect 1236 -828 1294 -822
rect 498 -894 556 -888
rect 498 -928 510 -894
rect 498 -934 556 -928
rect 668 -953 702 -935
rect 1090 -953 1124 -935
rect 668 -989 738 -953
rect 498 -1002 556 -996
rect 498 -1036 510 -1002
rect 685 -1023 756 -989
rect 498 -1042 556 -1036
rect 498 -1214 556 -1208
rect 498 -1248 510 -1214
rect 498 -1254 556 -1248
rect 498 -1322 556 -1316
rect 498 -1356 510 -1322
rect 498 -1362 556 -1356
rect 498 -1534 556 -1528
rect 498 -1568 510 -1534
rect 498 -1574 556 -1568
rect 352 -1651 367 -1617
rect 685 -1670 755 -1023
rect 867 -1091 925 -1085
rect 867 -1125 879 -1091
rect 867 -1131 925 -1125
rect 867 -1285 925 -1279
rect 867 -1319 879 -1285
rect 867 -1325 925 -1319
rect 867 -1393 925 -1387
rect 867 -1427 879 -1393
rect 867 -1433 925 -1427
rect 867 -1587 925 -1581
rect 867 -1621 879 -1587
rect 867 -1627 925 -1621
rect 685 -1706 738 -1670
rect 1054 -1723 1124 -953
rect 1236 -1000 1294 -994
rect 1236 -1034 1248 -1000
rect 1236 -1040 1294 -1034
rect 1406 -1059 1440 -1041
rect 1406 -1095 1476 -1059
rect 1236 -1108 1294 -1102
rect 1236 -1142 1248 -1108
rect 1423 -1129 1494 -1095
rect 1236 -1148 1294 -1142
rect 1236 -1320 1294 -1314
rect 1236 -1354 1248 -1320
rect 1236 -1360 1294 -1354
rect 1236 -1428 1294 -1422
rect 1236 -1462 1248 -1428
rect 1236 -1468 1294 -1462
rect 1236 -1640 1294 -1634
rect 1236 -1674 1248 -1640
rect 1236 -1680 1294 -1674
rect 1054 -1759 1107 -1723
rect 1423 -1776 1493 -1129
rect 1605 -1197 1663 -1191
rect 1605 -1231 1617 -1197
rect 1605 -1237 1663 -1231
rect 1605 -1391 1663 -1385
rect 1605 -1425 1617 -1391
rect 1605 -1431 1663 -1425
rect 1605 -1499 1663 -1493
rect 1605 -1533 1617 -1499
rect 1605 -1539 1663 -1533
rect 1605 -1693 1663 -1687
rect 1605 -1727 1617 -1693
rect 1605 -1733 1663 -1727
rect 1423 -1812 1476 -1776
rect 5895 -10804 5930 -10770
rect 5896 -10823 5930 -10804
rect 5730 -11332 5800 -11330
rect 5915 -11962 5930 -10823
rect 5949 -10857 5984 -10823
rect 5949 -11962 5983 -10857
rect 6079 -11385 6149 -11383
rect 5949 -11996 5964 -11962
rect 6264 -12015 6279 -10823
rect 6298 -12015 6332 -10769
rect 6444 -10832 6502 -10826
rect 6444 -10866 6456 -10832
rect 6444 -10872 6502 -10866
rect 6444 -11026 6502 -11020
rect 6444 -11060 6456 -11026
rect 6444 -11066 6502 -11060
rect 6444 -11134 6502 -11128
rect 6444 -11168 6456 -11134
rect 6444 -11174 6502 -11168
rect 6614 -11315 6648 -11297
rect 6444 -11328 6502 -11322
rect 6444 -11362 6456 -11328
rect 6614 -11351 6684 -11315
rect 6444 -11368 6502 -11362
rect 6631 -11385 6702 -11351
rect 6982 -11385 7017 -11351
rect 6444 -11436 6502 -11430
rect 6444 -11470 6456 -11436
rect 6444 -11476 6502 -11470
rect 6444 -11630 6502 -11624
rect 6444 -11664 6456 -11630
rect 6444 -11670 6502 -11664
rect 6444 -11738 6502 -11732
rect 6444 -11772 6456 -11738
rect 6444 -11778 6502 -11772
rect 6444 -11932 6502 -11926
rect 6444 -11966 6456 -11932
rect 6444 -11972 6502 -11966
rect 6298 -12049 6313 -12015
rect 6631 -12068 6701 -11385
rect 6983 -11404 7017 -11385
rect 6813 -11453 6871 -11447
rect 6813 -11487 6825 -11453
rect 6813 -11493 6871 -11487
rect 6813 -11665 6871 -11659
rect 6813 -11699 6825 -11665
rect 6813 -11705 6871 -11699
rect 6813 -11773 6871 -11767
rect 6813 -11807 6825 -11773
rect 6813 -11813 6871 -11807
rect 6813 -11985 6871 -11979
rect 6813 -12019 6825 -11985
rect 6813 -12025 6871 -12019
rect 6631 -12104 6684 -12068
rect 7002 -12121 7017 -11404
rect 7036 -11438 7071 -11404
rect 7036 -12121 7070 -11438
rect 7352 -11457 7386 -11439
rect 7352 -11493 7422 -11457
rect 7182 -11506 7240 -11500
rect 7182 -11540 7194 -11506
rect 7369 -11527 7440 -11493
rect 7720 -11527 7755 -11493
rect 7182 -11546 7240 -11540
rect 7182 -11718 7240 -11712
rect 7182 -11752 7194 -11718
rect 7182 -11758 7240 -11752
rect 7182 -11826 7240 -11820
rect 7182 -11860 7194 -11826
rect 7182 -11866 7240 -11860
rect 7182 -12038 7240 -12032
rect 7182 -12072 7194 -12038
rect 7182 -12078 7240 -12072
rect 7036 -12155 7051 -12121
rect 7369 -12174 7439 -11527
rect 7721 -11546 7755 -11527
rect 7551 -11595 7609 -11589
rect 7551 -11629 7563 -11595
rect 7551 -11635 7609 -11629
rect 7551 -11789 7609 -11783
rect 7551 -11823 7563 -11789
rect 7551 -11829 7609 -11823
rect 7551 -11897 7609 -11891
rect 7551 -11931 7563 -11897
rect 7551 -11937 7609 -11931
rect 7551 -12091 7609 -12085
rect 7551 -12125 7563 -12091
rect 7551 -12131 7609 -12125
rect 7369 -12210 7422 -12174
rect 7740 -12227 7755 -11546
rect 7774 -11580 7809 -11546
rect 7774 -12227 7808 -11580
rect 7920 -11648 7978 -11642
rect 7920 -11682 7932 -11648
rect 7920 -11688 7978 -11682
rect 7920 -11842 7978 -11836
rect 7920 -11876 7932 -11842
rect 7920 -11882 7978 -11876
rect 7920 -11950 7978 -11944
rect 7920 -11984 7932 -11950
rect 7920 -11990 7978 -11984
rect 7920 -12144 7978 -12138
rect 7920 -12178 7932 -12144
rect 7920 -12184 7978 -12178
rect 7774 -12261 7789 -12227
rect 8109 -12280 8124 -11546
rect 8143 -12280 8177 -11492
rect 8273 -11703 8343 -11701
rect 8143 -12314 8158 -12280
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
use sky130_fd_pr__cap_mim_m3_1_JDQXT2  XC1
timestamp 0
transform 1 0 3731 0 1 -5305
box -1886 -6640 1886 6640
use sky130_fd_pr__pfet_01v8_M47XPL  XM1
timestamp 0
transform 1 0 6842 0 1 -11736
box -211 -421 211 421
use sky130_fd_pr__pfet_01v8_M47XPL  XM2
timestamp 0
transform 1 0 7211 0 1 -11789
box -211 -421 211 421
use sky130_fd_pr__nfet_01v8_9XY3GD  XM3
timestamp 0
transform 1 0 6473 0 1 -11399
box -211 -705 211 705
use sky130_fd_pr__nfet_01v8_9XY3GD  XM4
timestamp 0
transform 1 0 8667 0 1 -11717
box -211 -705 211 705
use sky130_fd_pr__nfet_01v8_PTX3GD  XM5
timestamp 0
transform 1 0 896 0 1 -1356
box -211 -403 211 403
use sky130_fd_pr__nfet_01v8_PTX3GD  XM6
timestamp 0
transform 1 0 7580 0 1 -11860
box -211 -403 211 403
use sky130_fd_pr__nfet_01v8_PTX3GD  XM7
timestamp 0
transform 1 0 7949 0 1 -11913
box -211 -403 211 403
use sky130_fd_pr__pfet_01v8_M47T9Z  XM8
timestamp 0
transform 1 0 158 0 1 -912
box -211 -741 211 741
use sky130_fd_pr__pfet_01v8_M47T9Z  XM9
timestamp 0
transform 1 0 527 0 1 -965
box -211 -741 211 741
use sky130_fd_pr__pfet_01v8_M47T9Z  XM10
timestamp 0
transform 1 0 1265 0 1 -1071
box -211 -741 211 741
use sky130_fd_pr__nfet_01v8_PTX3GD  XM11
timestamp 0
transform 1 0 1634 0 1 -1462
box -211 -403 211 403
use sky130_fd_pr__res_high_po_0p35_Q7UHRC  XR1
timestamp 0
transform 1 0 5765 0 1 -11366
box -201 -632 201 632
use sky130_fd_pr__res_high_po_0p35_Q7UHRC  XR2
timestamp 0
transform 1 0 6114 0 1 -11419
box -201 -632 201 632
use sky130_fd_pr__res_high_po_0p35_Q7UHRC  XR4
timestamp 0
transform 1 0 8308 0 1 -11737
box -201 -632 201 632
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 out
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 -
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 +
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 GND
port 4 nsew
<< end >>
