magic
tech sky130A
magscale 1 2
timestamp 1762689433
<< metal1 >>
rect 1577 10482 1587 10534
rect 1639 10482 1649 10534
rect 5869 10050 5879 10102
rect 5931 10050 5941 10102
rect -1283 9945 -1231 9951
rect 3035 9909 3087 9915
rect -1283 9114 -1231 9893
rect 1669 9857 1675 9909
rect 1727 9906 1733 9909
rect 3029 9906 3035 9909
rect 1727 9860 3035 9906
rect 1727 9857 1733 9860
rect 3029 9857 3035 9860
rect 3087 9857 3093 9909
rect 3035 9851 3087 9857
rect 3339 9853 3345 9905
rect 3397 9853 5879 9905
rect 5931 9853 5937 9905
rect 1284 9771 1290 9823
rect 1342 9771 3665 9823
rect 3717 9771 3723 9823
rect 6213 9651 6269 9657
rect 6269 9595 8977 9651
rect 9033 9595 9039 9651
rect 6213 9589 6269 9595
rect -1283 9056 -1231 9062
rect 2613 8981 2623 9033
rect 2675 8981 2685 9033
rect 3345 8514 3397 8520
rect 3397 8462 8048 8514
rect 8100 8462 8106 8514
rect 3345 8456 3397 8462
rect 3934 8422 3986 8428
rect 2880 8370 2886 8422
rect 2938 8370 3934 8422
rect 3934 8364 3986 8370
rect 3035 8254 3087 8260
rect 2799 8205 3035 8251
rect 3035 8196 3087 8202
<< via1 >>
rect 1587 10482 1639 10534
rect 5879 10050 5931 10102
rect -1283 9893 -1231 9945
rect 1675 9857 1727 9909
rect 3035 9857 3087 9909
rect 3345 9853 3397 9905
rect 5879 9853 5931 9905
rect 1290 9771 1342 9823
rect 3665 9771 3717 9823
rect 6213 9595 6269 9651
rect 8977 9595 9033 9651
rect -1283 9062 -1231 9114
rect 2623 8981 2675 9033
rect 3345 8462 3397 8514
rect 8048 8462 8100 8514
rect 2886 8370 2938 8422
rect 3934 8370 3986 8422
rect 3035 8202 3087 8254
<< metal2 >>
rect 1587 10534 1639 10544
rect 1290 10482 1587 10534
rect -1285 9947 -1229 9957
rect -1289 9893 -1285 9945
rect -1229 9893 -1225 9945
rect -1285 9881 -1229 9891
rect 1290 9823 1342 10482
rect 1587 10472 1639 10482
rect 5787 10536 5843 10782
rect 5787 10480 6269 10536
rect 1678 9915 1724 10255
rect 5879 10102 5931 10112
rect 1675 9909 1727 9915
rect 3035 9909 3087 9915
rect 3029 9857 3035 9909
rect 3087 9857 3093 9909
rect 3345 9905 3397 9911
rect 1675 9851 1727 9857
rect 3035 9851 3087 9857
rect 1290 9765 1342 9771
rect -1289 9062 -1283 9114
rect -1231 9062 -722 9114
rect 2621 9035 2677 9045
rect 2621 8969 2677 8979
rect 2886 8422 2938 8879
rect 2886 8364 2938 8370
rect 3038 8254 3084 9851
rect 3345 8514 3397 9853
rect 5879 9905 5931 10050
rect 5879 9847 5931 9853
rect 3665 9823 3717 9829
rect 3665 9249 3717 9771
rect 6213 9651 6269 10480
rect 8977 9651 9033 9657
rect 6207 9595 6213 9651
rect 6269 9595 6275 9651
rect 8977 9280 9033 9595
rect 8048 8514 8100 8520
rect 3339 8462 3345 8514
rect 3397 8462 3403 8514
rect 3928 8370 3934 8422
rect 3986 8370 3992 8422
rect 3029 8202 3035 8254
rect 3087 8202 3093 8254
rect 3934 8115 3986 8370
rect 8048 8118 8100 8462
<< via2 >>
rect -1285 9945 -1229 9947
rect -1285 9893 -1283 9945
rect -1283 9893 -1231 9945
rect -1231 9893 -1229 9945
rect -1285 9891 -1229 9893
rect 2621 9033 2677 9035
rect 2621 8981 2623 9033
rect 2623 8981 2675 9033
rect 2675 8981 2677 9033
rect 2621 8979 2677 8981
<< metal3 >>
rect -1305 9952 -1205 9969
rect -1305 9886 -1290 9952
rect -1226 9886 -1205 9952
rect -1305 9869 -1205 9886
rect 2611 9037 2687 9040
rect 2611 9035 3710 9037
rect 2611 8979 2621 9035
rect 2677 8979 3710 9035
rect 2611 8977 3710 8979
rect 2611 8974 2687 8977
<< via3 >>
rect -1290 9947 -1226 9952
rect -1290 9891 -1285 9947
rect -1285 9891 -1229 9947
rect -1229 9891 -1226 9947
rect -1290 9886 -1226 9891
<< metal4 >>
rect -1384 9952 -1207 9967
rect -1384 9886 -1290 9952
rect -1226 9886 -1207 9952
rect -1384 9871 -1207 9886
use cap_op  cap_op_0
timestamp 1718554435
transform 1 0 -5171 0 1 11901
box -12037 -11160 3906 3480
use differential_pair  differential_pair_0
timestamp 1720116957
transform 1 0 4032 0 1 8666
box -606 -124 5240 892
use nmos_tail_current  nmos_tail_current_0
timestamp 1720118050
transform -1 0 8043 0 -1 8201
box -321 -141 8599 1579
use pmos_current_bgr_2  pmos_current_bgr_2_0
timestamp 1720112176
transform 1 0 1636 0 1 11374
box -250 -1450 4496 516
use resistor_op_tt  resistor_op_tt_0
timestamp 1720284839
transform 0 -1 5238 -1 0 9265
box -417 2220 767 6092
<< end >>
