magic
tech sky130A
magscale 1 2
timestamp 1716351939
<< error_p >>
rect -450 1588 -380 1590
rect -284 1588 -214 1590
rect -118 1588 -48 1590
rect 48 1588 118 1590
rect 214 1588 284 1590
rect 380 1588 450 1590
rect -450 552 -380 554
rect -284 552 -214 554
rect -118 552 -48 554
rect 48 552 118 554
rect 214 552 284 554
rect 380 552 450 554
rect -450 -484 -380 -482
rect -284 -484 -214 -482
rect -118 -484 -48 -482
rect 48 -484 118 -482
rect 214 -484 284 -482
rect 380 -484 450 -482
rect -450 -1520 -380 -1518
rect -284 -1520 -214 -1518
rect -118 -1520 -48 -1518
rect 48 -1520 118 -1518
rect 214 -1520 284 -1518
rect 380 -1520 450 -1518
<< nwell >>
rect -677 -2195 677 2195
<< nsubdiff >>
rect -641 2125 -545 2159
rect 545 2125 641 2159
rect -641 2063 -607 2125
rect 607 2063 641 2125
rect -641 -2125 -607 -2063
rect 607 -2125 641 -2063
rect -641 -2159 -545 -2125
rect 545 -2159 641 -2125
<< nsubdiffcont >>
rect -545 2125 545 2159
rect -641 -2063 -607 2063
rect 607 -2063 641 2063
rect -545 -2159 545 -2125
<< xpolycontact >>
rect -450 1588 -380 2020
rect -450 1088 -380 1520
rect -284 1588 -214 2020
rect -284 1088 -214 1520
rect -118 1588 -48 2020
rect -118 1088 -48 1520
rect 48 1588 118 2020
rect 48 1088 118 1520
rect 214 1588 284 2020
rect 214 1088 284 1520
rect 380 1588 450 2020
rect 380 1088 450 1520
rect -450 552 -380 984
rect -450 52 -380 484
rect -284 552 -214 984
rect -284 52 -214 484
rect -118 552 -48 984
rect -118 52 -48 484
rect 48 552 118 984
rect 48 52 118 484
rect 214 552 284 984
rect 214 52 284 484
rect 380 552 450 984
rect 380 52 450 484
rect -450 -484 -380 -52
rect -450 -984 -380 -552
rect -284 -484 -214 -52
rect -284 -984 -214 -552
rect -118 -484 -48 -52
rect -118 -984 -48 -552
rect 48 -484 118 -52
rect 48 -984 118 -552
rect 214 -484 284 -52
rect 214 -984 284 -552
rect 380 -484 450 -52
rect 380 -984 450 -552
rect -450 -1520 -380 -1088
rect -450 -2020 -380 -1588
rect -284 -1520 -214 -1088
rect -284 -2020 -214 -1588
rect -118 -1520 -48 -1088
rect -118 -2020 -48 -1588
rect 48 -1520 118 -1088
rect 48 -2020 118 -1588
rect 214 -1520 284 -1088
rect 214 -2020 284 -1588
rect 380 -1520 450 -1088
rect 380 -2020 450 -1588
<< ppolyres >>
rect -450 1520 -380 1588
rect -284 1520 -214 1588
rect -118 1520 -48 1588
rect 48 1520 118 1588
rect 214 1520 284 1588
rect 380 1520 450 1588
rect -450 484 -380 552
rect -284 484 -214 552
rect -118 484 -48 552
rect 48 484 118 552
rect 214 484 284 552
rect 380 484 450 552
rect -450 -552 -380 -484
rect -284 -552 -214 -484
rect -118 -552 -48 -484
rect 48 -552 118 -484
rect 214 -552 284 -484
rect 380 -552 450 -484
rect -450 -1588 -380 -1520
rect -284 -1588 -214 -1520
rect -118 -1588 -48 -1520
rect 48 -1588 118 -1520
rect 214 -1588 284 -1520
rect 380 -1588 450 -1520
<< locali >>
rect -561 2125 -545 2159
rect 545 2125 561 2159
rect -641 2063 -607 2079
rect 607 2063 641 2079
rect -641 -2079 -607 -2063
rect 607 -2079 641 -2063
rect -561 -2159 -545 -2125
rect 545 -2159 561 -2125
<< viali >>
rect -434 1605 -396 2002
rect -268 1605 -230 2002
rect -102 1605 -64 2002
rect 64 1605 102 2002
rect 230 1605 268 2002
rect 396 1605 434 2002
rect -434 1106 -396 1503
rect -268 1106 -230 1503
rect -102 1106 -64 1503
rect 64 1106 102 1503
rect 230 1106 268 1503
rect 396 1106 434 1503
rect -434 569 -396 966
rect -268 569 -230 966
rect -102 569 -64 966
rect 64 569 102 966
rect 230 569 268 966
rect 396 569 434 966
rect -434 70 -396 467
rect -268 70 -230 467
rect -102 70 -64 467
rect 64 70 102 467
rect 230 70 268 467
rect 396 70 434 467
rect -434 -467 -396 -70
rect -268 -467 -230 -70
rect -102 -467 -64 -70
rect 64 -467 102 -70
rect 230 -467 268 -70
rect 396 -467 434 -70
rect -434 -966 -396 -569
rect -268 -966 -230 -569
rect -102 -966 -64 -569
rect 64 -966 102 -569
rect 230 -966 268 -569
rect 396 -966 434 -569
rect -434 -1503 -396 -1106
rect -268 -1503 -230 -1106
rect -102 -1503 -64 -1106
rect 64 -1503 102 -1106
rect 230 -1503 268 -1106
rect 396 -1503 434 -1106
rect -434 -2002 -396 -1605
rect -268 -2002 -230 -1605
rect -102 -2002 -64 -1605
rect 64 -2002 102 -1605
rect 230 -2002 268 -1605
rect 396 -2002 434 -1605
<< metal1 >>
rect -440 2002 -390 2014
rect -440 1605 -434 2002
rect -396 1605 -390 2002
rect -440 1593 -390 1605
rect -274 2002 -224 2014
rect -274 1605 -268 2002
rect -230 1605 -224 2002
rect -274 1593 -224 1605
rect -108 2002 -58 2014
rect -108 1605 -102 2002
rect -64 1605 -58 2002
rect -108 1593 -58 1605
rect 58 2002 108 2014
rect 58 1605 64 2002
rect 102 1605 108 2002
rect 58 1593 108 1605
rect 224 2002 274 2014
rect 224 1605 230 2002
rect 268 1605 274 2002
rect 224 1593 274 1605
rect 390 2002 440 2014
rect 390 1605 396 2002
rect 434 1605 440 2002
rect 390 1593 440 1605
rect -440 1503 -390 1515
rect -440 1106 -434 1503
rect -396 1106 -390 1503
rect -440 1094 -390 1106
rect -274 1503 -224 1515
rect -274 1106 -268 1503
rect -230 1106 -224 1503
rect -274 1094 -224 1106
rect -108 1503 -58 1515
rect -108 1106 -102 1503
rect -64 1106 -58 1503
rect -108 1094 -58 1106
rect 58 1503 108 1515
rect 58 1106 64 1503
rect 102 1106 108 1503
rect 58 1094 108 1106
rect 224 1503 274 1515
rect 224 1106 230 1503
rect 268 1106 274 1503
rect 224 1094 274 1106
rect 390 1503 440 1515
rect 390 1106 396 1503
rect 434 1106 440 1503
rect 390 1094 440 1106
rect -440 966 -390 978
rect -440 569 -434 966
rect -396 569 -390 966
rect -440 557 -390 569
rect -274 966 -224 978
rect -274 569 -268 966
rect -230 569 -224 966
rect -274 557 -224 569
rect -108 966 -58 978
rect -108 569 -102 966
rect -64 569 -58 966
rect -108 557 -58 569
rect 58 966 108 978
rect 58 569 64 966
rect 102 569 108 966
rect 58 557 108 569
rect 224 966 274 978
rect 224 569 230 966
rect 268 569 274 966
rect 224 557 274 569
rect 390 966 440 978
rect 390 569 396 966
rect 434 569 440 966
rect 390 557 440 569
rect -440 467 -390 479
rect -440 70 -434 467
rect -396 70 -390 467
rect -440 58 -390 70
rect -274 467 -224 479
rect -274 70 -268 467
rect -230 70 -224 467
rect -274 58 -224 70
rect -108 467 -58 479
rect -108 70 -102 467
rect -64 70 -58 467
rect -108 58 -58 70
rect 58 467 108 479
rect 58 70 64 467
rect 102 70 108 467
rect 58 58 108 70
rect 224 467 274 479
rect 224 70 230 467
rect 268 70 274 467
rect 224 58 274 70
rect 390 467 440 479
rect 390 70 396 467
rect 434 70 440 467
rect 390 58 440 70
rect -440 -70 -390 -58
rect -440 -467 -434 -70
rect -396 -467 -390 -70
rect -440 -479 -390 -467
rect -274 -70 -224 -58
rect -274 -467 -268 -70
rect -230 -467 -224 -70
rect -274 -479 -224 -467
rect -108 -70 -58 -58
rect -108 -467 -102 -70
rect -64 -467 -58 -70
rect -108 -479 -58 -467
rect 58 -70 108 -58
rect 58 -467 64 -70
rect 102 -467 108 -70
rect 58 -479 108 -467
rect 224 -70 274 -58
rect 224 -467 230 -70
rect 268 -467 274 -70
rect 224 -479 274 -467
rect 390 -70 440 -58
rect 390 -467 396 -70
rect 434 -467 440 -70
rect 390 -479 440 -467
rect -440 -569 -390 -557
rect -440 -966 -434 -569
rect -396 -966 -390 -569
rect -440 -978 -390 -966
rect -274 -569 -224 -557
rect -274 -966 -268 -569
rect -230 -966 -224 -569
rect -274 -978 -224 -966
rect -108 -569 -58 -557
rect -108 -966 -102 -569
rect -64 -966 -58 -569
rect -108 -978 -58 -966
rect 58 -569 108 -557
rect 58 -966 64 -569
rect 102 -966 108 -569
rect 58 -978 108 -966
rect 224 -569 274 -557
rect 224 -966 230 -569
rect 268 -966 274 -569
rect 224 -978 274 -966
rect 390 -569 440 -557
rect 390 -966 396 -569
rect 434 -966 440 -569
rect 390 -978 440 -966
rect -440 -1106 -390 -1094
rect -440 -1503 -434 -1106
rect -396 -1503 -390 -1106
rect -440 -1515 -390 -1503
rect -274 -1106 -224 -1094
rect -274 -1503 -268 -1106
rect -230 -1503 -224 -1106
rect -274 -1515 -224 -1503
rect -108 -1106 -58 -1094
rect -108 -1503 -102 -1106
rect -64 -1503 -58 -1106
rect -108 -1515 -58 -1503
rect 58 -1106 108 -1094
rect 58 -1503 64 -1106
rect 102 -1503 108 -1106
rect 58 -1515 108 -1503
rect 224 -1106 274 -1094
rect 224 -1503 230 -1106
rect 268 -1503 274 -1106
rect 224 -1515 274 -1503
rect 390 -1106 440 -1094
rect 390 -1503 396 -1106
rect 434 -1503 440 -1106
rect 390 -1515 440 -1503
rect -440 -1605 -390 -1593
rect -440 -2002 -434 -1605
rect -396 -2002 -390 -1605
rect -440 -2014 -390 -2002
rect -274 -1605 -224 -1593
rect -274 -2002 -268 -1605
rect -230 -2002 -224 -1605
rect -274 -2014 -224 -2002
rect -108 -1605 -58 -1593
rect -108 -2002 -102 -1605
rect -64 -2002 -58 -1605
rect -108 -2014 -58 -2002
rect 58 -1605 108 -1593
rect 58 -2002 64 -1605
rect 102 -2002 108 -1605
rect 58 -2014 108 -2002
rect 224 -1605 274 -1593
rect 224 -2002 230 -1605
rect 268 -2002 274 -1605
rect 224 -2014 274 -2002
rect 390 -1605 440 -1593
rect 390 -2002 396 -1605
rect 434 -2002 440 -1605
rect 390 -2014 440 -2002
<< properties >>
string FIXED_BBOX -624 -2142 624 2142
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.350 l 0.5 m 4 nx 6 wmin 0.350 lmin 0.50 rho 319.8 val 1.57k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 0 wmax 0.350 vias 1 n_guard 1 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
