magic
tech sky130A
magscale 1 2
timestamp 1717913728
<< nmos >>
rect -229 -131 -29 69
rect 29 -131 229 69
<< ndiff >>
rect -287 57 -229 69
rect -287 -119 -275 57
rect -241 -119 -229 57
rect -287 -131 -229 -119
rect -29 57 29 69
rect -29 -119 -17 57
rect 17 -119 29 57
rect -29 -131 29 -119
rect 229 57 287 69
rect 229 -119 241 57
rect 275 -119 287 57
rect 229 -131 287 -119
<< ndiffc >>
rect -275 -119 -241 57
rect -17 -119 17 57
rect 241 -119 275 57
<< poly >>
rect -229 141 -29 157
rect -229 107 -213 141
rect -45 107 -29 141
rect -229 69 -29 107
rect 29 141 229 157
rect 29 107 45 141
rect 213 107 229 141
rect 29 69 229 107
rect -229 -157 -29 -131
rect 29 -157 229 -131
<< polycont >>
rect -213 107 -45 141
rect 45 107 213 141
<< locali >>
rect -229 107 -213 141
rect -45 107 -29 141
rect 29 107 45 141
rect 213 107 229 141
rect -275 57 -241 73
rect -275 -135 -241 -119
rect -17 57 17 73
rect -17 -135 17 -119
rect 241 57 275 73
rect 241 -135 275 -119
<< viali >>
rect -213 107 -45 141
rect 45 107 213 141
rect -275 -119 -241 57
rect -17 -119 17 57
rect 241 -119 275 57
<< metal1 >>
rect -225 141 -33 147
rect -225 107 -213 141
rect -45 107 -33 141
rect -225 101 -33 107
rect 33 141 225 147
rect 33 107 45 141
rect 213 107 225 141
rect 33 101 225 107
rect -281 57 -235 69
rect -281 -119 -275 57
rect -241 -119 -235 57
rect -281 -131 -235 -119
rect -23 57 23 69
rect -23 -119 -17 57
rect 17 -119 23 57
rect -23 -131 23 -119
rect 235 57 281 69
rect 235 -119 241 57
rect 275 -119 281 57
rect 235 -131 281 -119
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 1 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
