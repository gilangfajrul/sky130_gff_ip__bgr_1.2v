magic
tech sky130A
magscale 1 2
timestamp 1716468452
<< psubdiff >>
rect -194 1508 -134 1542
rect 8412 1508 8472 1542
rect -194 1478 -160 1508
rect 8438 1478 8472 1508
rect -194 -70 -160 -40
rect 8438 -70 8472 -40
rect -194 -104 -134 -70
rect 8412 -104 8472 -70
<< psubdiffcont >>
rect -134 1508 8412 1542
rect -194 -40 -160 1478
rect 8438 -40 8472 1478
rect -134 -104 8412 -70
<< poly >>
rect -123 1429 -4 1481
rect 1040 1436 3068 1478
rect -34 1410 -4 1429
rect 8282 1429 8401 1481
rect 8282 1410 8312 1429
rect 54 1042 8224 1184
rect -34 797 -4 816
rect -123 745 -4 797
rect 8304 791 8401 797
rect -123 641 -4 693
rect 54 648 8224 790
rect 8282 745 8401 791
rect 8282 647 8401 693
rect 8304 641 8401 647
rect 54 254 8224 396
rect -34 9 -4 28
rect -123 -43 -4 9
rect 8282 9 8312 28
rect 5210 -40 7238 2
rect 8282 -43 8401 9
<< locali >>
rect -194 1508 -134 1542
rect 8412 1508 8472 1542
rect -194 1478 -160 1508
rect 8438 1478 8472 1508
rect -80 1410 -46 1436
rect 8324 1410 8358 1436
rect -80 790 -46 816
rect 8324 790 8358 828
rect -80 624 -46 648
rect 8324 614 8358 648
rect -80 2 -46 28
rect 8324 2 8358 28
rect -194 -70 -160 -40
rect 8438 -70 8472 -40
rect -194 -104 -134 -70
rect 8412 -104 8472 -70
<< viali >>
rect 4055 1508 4111 1542
rect -194 -36 -160 1474
rect -110 1436 -38 1474
rect 1054 1436 3054 1470
rect 8316 1436 8388 1474
rect -110 752 -38 790
rect 8316 752 8388 790
rect -110 648 -38 686
rect 8316 648 8388 686
rect -110 -36 -38 2
rect 5224 -32 7224 2
rect 8316 -36 8388 2
rect 8438 -36 8472 1474
rect 4167 -104 4223 -70
<< metal1 >>
rect 4043 1542 4123 1548
rect 4043 1508 4055 1542
rect 4111 1508 4123 1542
rect 4043 1502 4123 1508
rect -200 1480 -154 1486
rect -200 1474 -26 1480
rect -200 -36 -194 1474
rect -160 1436 -110 1474
rect -38 1436 -26 1474
rect -160 1430 -26 1436
rect 2 1470 3066 1476
rect 2 1444 1054 1470
rect -160 796 -154 1430
rect -86 1410 -40 1430
rect 2 1408 48 1444
rect 1042 1436 1054 1444
rect 3054 1436 3066 1470
rect 1042 1430 3066 1436
rect 4060 1408 4106 1502
rect 8432 1480 8478 1486
rect 8304 1474 8478 1480
rect 8304 1436 8316 1474
rect 8388 1436 8438 1474
rect 8304 1430 8438 1436
rect 8318 1410 8364 1430
rect 4060 1016 4106 1374
rect 4159 1222 4169 1398
rect 4221 1222 4231 1398
rect 8217 1222 8227 1398
rect 8279 1222 8289 1398
rect 33 816 48 827
rect 4060 816 4112 1016
rect 4166 816 4218 1016
rect 8217 828 8227 1004
rect 8279 828 8289 1004
rect 8324 824 8358 828
rect -86 796 -40 816
rect -160 790 -26 796
rect -160 752 -110 790
rect -38 752 -26 790
rect -160 746 -26 752
rect -160 692 -154 746
rect 10 742 48 816
rect 8318 796 8364 824
rect 8432 796 8438 1430
rect 8304 790 8438 796
rect 8304 752 8316 790
rect 8388 752 8438 790
rect 8304 746 8438 752
rect 10 696 8276 742
rect -160 686 -26 692
rect -160 648 -110 686
rect -38 648 -26 686
rect -160 642 -26 648
rect -160 8 -154 642
rect -86 614 -40 642
rect -11 609 61 610
rect -11 434 -1 609
rect 51 434 61 609
rect 4060 422 4112 622
rect 4166 422 4218 622
rect 8230 612 8276 696
rect 8432 692 8438 746
rect 8304 686 8438 692
rect 8304 648 8316 686
rect 8388 648 8438 686
rect 8304 642 8438 648
rect 8318 613 8364 642
rect -11 40 -1 216
rect 51 40 61 216
rect 4047 40 4057 216
rect 4109 40 4119 216
rect -86 8 -40 28
rect -160 2 -26 8
rect -160 -36 -110 2
rect -38 -36 -26 2
rect -200 -42 -26 -36
rect -200 -48 -154 -42
rect 4172 -64 4218 422
rect 5212 2 7236 8
rect 5212 -32 5224 2
rect 7224 -6 7236 2
rect 8230 -6 8276 30
rect 8318 8 8364 28
rect 8432 8 8438 642
rect 7224 -32 8276 -6
rect 5212 -38 8276 -32
rect 8304 2 8438 8
rect 8304 -36 8316 2
rect 8388 -36 8438 2
rect 8472 -36 8478 1474
rect 8304 -42 8478 -36
rect 8432 -48 8478 -42
rect 4155 -70 4235 -64
rect 4155 -104 4167 -70
rect 4223 -104 4235 -70
rect 4155 -110 4235 -104
<< via1 >>
rect 4169 1222 4221 1398
rect 8227 1222 8279 1398
rect 4112 816 4166 1016
rect 8227 828 8279 1004
rect -1 434 51 609
rect 4112 422 4166 622
rect -1 40 51 216
rect 4057 40 4109 216
<< metal2 >>
rect 4169 1398 4221 1408
rect 4169 1140 4221 1222
rect 8225 1398 8281 1408
rect 8225 1212 8281 1222
rect -155 1135 8379 1140
rect -155 1086 8435 1135
rect -155 352 -101 1086
rect 4111 1016 4167 1026
rect 4111 806 4167 816
rect 8227 1004 8279 1014
rect 8227 747 8279 828
rect -1 691 8279 747
rect -1 609 51 691
rect -1 424 51 434
rect 4111 622 4167 632
rect 4111 412 4167 422
rect 8381 352 8435 1086
rect -155 298 8435 352
rect -3 216 53 226
rect -3 30 53 40
rect 4057 216 4109 298
rect 8381 293 8435 298
rect 4057 30 4109 40
<< via2 >>
rect 8225 1222 8227 1398
rect 8227 1222 8279 1398
rect 8279 1222 8281 1398
rect 4111 816 4112 1016
rect 4112 816 4166 1016
rect 4166 816 4167 1016
rect 4111 422 4112 622
rect 4112 422 4166 622
rect 4166 422 4167 622
rect -3 40 -1 216
rect -1 40 51 216
rect 51 40 53 216
<< metal3 >>
rect 8215 1398 8291 1403
rect 8215 1222 8225 1398
rect 8281 1222 8291 1398
rect 8215 1144 8291 1222
rect 8215 1082 8433 1144
rect 4101 1016 4177 1021
rect 4097 816 4107 1016
rect 4171 816 4181 1016
rect 4101 811 4177 816
rect 8371 750 8433 1082
rect -155 688 8433 750
rect -155 356 -93 688
rect 4101 622 4177 627
rect 4097 422 4107 622
rect 4171 422 4181 622
rect 4101 417 4177 422
rect -155 294 63 356
rect -13 216 63 294
rect -13 40 -3 216
rect 53 40 63 216
rect -13 35 63 40
<< via3 >>
rect 4107 816 4111 1016
rect 4111 816 4167 1016
rect 4167 816 4171 1016
rect 4107 422 4111 622
rect 4111 422 4167 622
rect 4167 422 4171 622
<< metal4 >>
rect 4106 1016 4172 1017
rect 4106 816 4107 1016
rect 4171 816 4172 1016
rect 4106 622 4172 816
rect 4106 422 4107 622
rect 4171 422 4172 622
rect 4106 421 4172 422
use sky130_fd_pr__nfet_01v8_HZDFY5  sky130_fd_pr__nfet_01v8_HZDFY5_0
timestamp 1716275522
transform 1 0 8297 0 1 128
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_HZDFY5  sky130_fd_pr__nfet_01v8_HZDFY5_1
timestamp 1716275522
transform 1 0 8297 0 1 1310
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_HZDFY5  sky130_fd_pr__nfet_01v8_HZDFY5_2
timestamp 1716275522
transform 1 0 8297 0 1 916
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_HZDFY5  sky130_fd_pr__nfet_01v8_HZDFY5_3
timestamp 1716275522
transform 1 0 8297 0 1 522
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_HZDFY5  sky130_fd_pr__nfet_01v8_HZDFY5_4
timestamp 1716275522
transform -1 0 -19 0 -1 1310
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_HZDFY5  sky130_fd_pr__nfet_01v8_HZDFY5_5
timestamp 1716275522
transform 1 0 -19 0 1 128
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_HZDFY5  sky130_fd_pr__nfet_01v8_HZDFY5_6
timestamp 1716275522
transform 1 0 -19 0 1 522
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_HZDFY5  sky130_fd_pr__nfet_01v8_HZDFY5_7
timestamp 1716275522
transform 1 0 -19 0 1 916
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_P5G96Q  sky130_fd_pr__nfet_01v8_P5G96Q_0
timestamp 1716212328
transform 1 0 6224 0 1 1310
box -2058 -126 2058 126
use sky130_fd_pr__nfet_01v8_P5G96Q  sky130_fd_pr__nfet_01v8_P5G96Q_1
timestamp 1716212328
transform 1 0 2054 0 1 128
box -2058 -126 2058 126
use sky130_fd_pr__nfet_01v8_P5G96Q  sky130_fd_pr__nfet_01v8_P5G96Q_2
timestamp 1716212328
transform 1 0 6224 0 1 128
box -2058 -126 2058 126
use sky130_fd_pr__nfet_01v8_P5G96Q  sky130_fd_pr__nfet_01v8_P5G96Q_3
timestamp 1716212328
transform 1 0 2054 0 1 1310
box -2058 -126 2058 126
use sky130_fd_pr__nfet_01v8_P5G96Q  sky130_fd_pr__nfet_01v8_P5G96Q_4
timestamp 1716212328
transform 1 0 6224 0 1 522
box -2058 -126 2058 126
use sky130_fd_pr__nfet_01v8_P5G96Q  sky130_fd_pr__nfet_01v8_P5G96Q_5
timestamp 1716212328
transform 1 0 2054 0 1 522
box -2058 -126 2058 126
use sky130_fd_pr__nfet_01v8_P5G96Q  sky130_fd_pr__nfet_01v8_P5G96Q_6
timestamp 1716212328
transform 1 0 6224 0 1 916
box -2058 -126 2058 126
use sky130_fd_pr__nfet_01v8_P5G96Q  sky130_fd_pr__nfet_01v8_P5G96Q_7
timestamp 1716212328
transform 1 0 2054 0 1 916
box -2058 -126 2058 126
<< end >>
