.param i_tail = 20.0e-06
.param lrz = 3.72e+01
.param mrz = 1.00e+00
.param lrs = 3.73e-01
.param mrs = 1.00e+00
.param mc = 4.00e+00
.param wc = 3.09e-01
.param w0 = 12
.param l0 = 5
.param nf0 = 1.00
.param w1 = 3
.param l1 = 5
.param nf1 = 1.00
.param w2 = 2.5
.param l2 = 5
.param nf2 = 1.00
.param w3 = 1.5
.param l3 = 5
.param nf3 = 1.00
.param w4 = 0.03
.param l4 = 0.60
.param nf4 = 1.00
