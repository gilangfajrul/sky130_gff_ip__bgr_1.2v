magic
tech sky130A
magscale 1 2
timestamp 1762701392
<< metal3 >>
rect -4165 3612 -333 3640
rect -4165 188 -417 3612
rect -353 188 -333 3612
rect -4165 160 -333 188
rect 333 3612 4165 3640
rect 333 188 4081 3612
rect 4145 188 4165 3612
rect 333 160 4165 188
rect -4165 -188 -333 -160
rect -4165 -3612 -417 -188
rect -353 -3612 -333 -188
rect -4165 -3640 -333 -3612
rect 333 -188 4165 -160
rect 333 -3612 4081 -188
rect 4145 -3612 4165 -188
rect 333 -3640 4165 -3612
<< via3 >>
rect -417 188 -353 3612
rect 4081 188 4145 3612
rect -417 -3612 -353 -188
rect 4081 -3612 4145 -188
<< mimcap >>
rect -4125 3560 -725 3600
rect -4125 240 -4085 3560
rect -765 240 -725 3560
rect -4125 200 -725 240
rect 373 3560 3773 3600
rect 373 240 413 3560
rect 3733 240 3773 3560
rect 373 200 3773 240
rect -4125 -240 -725 -200
rect -4125 -3560 -4085 -240
rect -765 -3560 -725 -240
rect -4125 -3600 -725 -3560
rect 373 -240 3773 -200
rect 373 -3560 413 -240
rect 3733 -3560 3773 -240
rect 373 -3600 3773 -3560
<< mimcapcontact >>
rect -4085 240 -765 3560
rect 413 240 3733 3560
rect -4085 -3560 -765 -240
rect 413 -3560 3733 -240
<< metal4 >>
rect -2477 3561 -2373 3800
rect -433 3612 -337 3628
rect -4086 3560 -764 3561
rect -4086 240 -4085 3560
rect -765 240 -764 3560
rect -4086 239 -764 240
rect -2477 -239 -2373 239
rect -433 188 -417 3612
rect -353 188 -337 3612
rect 2021 3561 2125 3800
rect 4065 3612 4161 3628
rect 412 3560 3734 3561
rect 412 240 413 3560
rect 3733 240 3734 3560
rect 412 239 3734 240
rect -433 172 -337 188
rect -433 -188 -337 -172
rect -4086 -240 -764 -239
rect -4086 -3560 -4085 -240
rect -765 -3560 -764 -240
rect -4086 -3561 -764 -3560
rect -2477 -3800 -2373 -3561
rect -433 -3612 -417 -188
rect -353 -3612 -337 -188
rect 2021 -239 2125 239
rect 4065 188 4081 3612
rect 4145 188 4161 3612
rect 4065 172 4161 188
rect 4065 -188 4161 -172
rect 412 -240 3734 -239
rect 412 -3560 413 -240
rect 3733 -3560 3734 -240
rect 412 -3561 3734 -3560
rect -433 -3628 -337 -3612
rect 2021 -3800 2125 -3561
rect 4065 -3612 4081 -188
rect 4145 -3612 4161 -188
rect 4065 -3628 4161 -3612
<< labels >>
rlabel via3 -385 -1900 -385 -1900 0 C2_0_0
port 1 nsew
rlabel mimcapcontact -2425 -1900 -2425 -1900 0 C1_0
port 2 nsew
rlabel via3 -385 1900 -385 1900 0 C2_0_1
port 3 nsew
rlabel via3 4113 -1900 4113 -1900 0 C2_1_0
port 4 nsew
rlabel mimcapcontact 2073 -1900 2073 -1900 0 C1_1
port 5 nsew
rlabel via3 4113 1900 4113 1900 0 C2_1_1
port 6 nsew
<< properties >>
string FIXED_BBOX 333 160 3813 3640
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 17 l 17 val 590.92 carea 2.00 cperi 0.19 class capacitor nx 2 ny 2 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 0 tconnect 1 ccov 100 stack 1 doports 1
<< end >>
