magic
tech sky130A
magscale 1 2
timestamp 1762846550
<< metal1 >>
rect 4519 868 4563 903
rect 4404 626 4414 802
rect 4466 626 4476 802
rect 5016 732 5026 784
rect 5110 732 5120 784
rect 5274 732 5284 784
rect 5368 732 5378 784
rect 112 150 122 326
rect 174 150 184 326
rect 4404 150 4414 326
rect 4466 150 4476 326
rect 4815 198 4825 374
rect 4877 198 4887 374
rect 5032 -91 5080 70
rect 154 -410 164 -358
rect 561 -410 571 -358
rect 10 -1239 259 -1189
<< via1 >>
rect 4414 626 4466 802
rect 5026 732 5110 784
rect 5284 732 5368 784
rect 122 150 174 326
rect 4414 150 4466 326
rect 4825 198 4877 374
rect 164 -410 561 -358
<< metal2 >>
rect 4414 802 4466 812
rect 5026 784 5110 794
rect 5284 784 5368 794
rect 4466 732 5026 784
rect 5110 732 5284 784
rect 5368 732 5374 784
rect 5026 722 5110 732
rect 5284 722 5368 732
rect 4414 616 4466 626
rect 4825 374 4877 384
rect 122 326 174 336
rect 122 -348 174 150
rect 4414 326 4466 336
rect 4466 234 4825 306
rect 4825 188 4877 198
rect 4414 140 4466 150
rect 122 -358 561 -348
rect 122 -410 164 -358
rect 122 -420 561 -410
use nmos_startup  nmos_startup_0
timestamp 1720119402
transform 1 0 4926 0 1 179
box -204 -154 746 692
use pmos_startup  pmos_startup_0
timestamp 1720267898
transform -1 0 4417 0 -1 444
box -176 -494 4422 430
use resistorstart  resistorstart_0
timestamp 1718868641
transform 1 0 33 0 1 -1528
box -53 -53 21855 1511
<< labels >>
flabel metal1 77 -1212 77 -1212 0 FreeSans 1600 0 0 0 avss
port 0 nsew
flabel metal2 4652 749 4652 749 0 FreeSans 1600 0 0 0 out
port 1 nsew
flabel metal1 4539 886 4539 886 0 FreeSans 1600 0 0 0 vdde
port 2 nsew
<< end >>
