magic
tech sky130A
magscale 1 2
timestamp 1717265618
<< error_p >>
rect -2123 -15 2123 236
<< nwell >>
rect -2123 -15 2123 347
rect -2123 -380 2123 -18
<< pmos >>
rect -2029 47 -29 247
rect 29 47 2029 247
rect -2029 -318 -29 -118
rect 29 -318 2029 -118
<< pdiff >>
rect -2087 235 -2029 247
rect -2087 59 -2075 235
rect -2041 59 -2029 235
rect -2087 47 -2029 59
rect -29 235 29 247
rect -29 59 -17 235
rect 17 59 29 235
rect -29 47 29 59
rect 2029 235 2087 247
rect 2029 59 2041 235
rect 2075 59 2087 235
rect 2029 47 2087 59
rect -2087 -130 -2029 -118
rect -2087 -306 -2075 -130
rect -2041 -306 -2029 -130
rect -2087 -318 -2029 -306
rect -29 -130 29 -118
rect -29 -306 -17 -130
rect 17 -306 29 -130
rect -29 -318 29 -306
rect 2029 -130 2087 -118
rect 2029 -306 2041 -130
rect 2075 -306 2087 -130
rect 2029 -318 2087 -306
<< pdiffc >>
rect -2075 59 -2041 235
rect -17 59 17 235
rect 2041 59 2075 235
rect -2075 -306 -2041 -130
rect -17 -306 17 -130
rect 2041 -306 2075 -130
<< poly >>
rect -2029 328 -29 344
rect -2029 294 -2013 328
rect -45 294 -29 328
rect -2029 247 -29 294
rect 29 328 2029 344
rect 29 294 45 328
rect 2013 294 2029 328
rect 29 247 2029 294
rect -2029 21 -29 47
rect 29 21 2029 47
rect -2029 -37 -29 -21
rect -2029 -71 -2013 -37
rect -45 -71 -29 -37
rect -2029 -118 -29 -71
rect 29 -37 2029 -21
rect 29 -71 45 -37
rect 2013 -71 2029 -37
rect 29 -118 2029 -71
rect -2029 -344 -29 -318
rect 29 -344 2029 -318
<< polycont >>
rect -2013 294 -45 328
rect 45 294 2013 328
rect -2013 -71 -45 -37
rect 45 -71 2013 -37
<< locali >>
rect -2029 294 -2013 328
rect -45 294 -29 328
rect 29 294 45 328
rect 2013 294 2029 328
rect -2075 235 -2041 251
rect -2075 43 -2041 59
rect -17 235 17 251
rect -17 43 17 59
rect 2041 235 2075 251
rect 2041 43 2075 59
rect -2029 -71 -2013 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 2013 -71 2029 -37
rect -2075 -130 -2041 -114
rect -2075 -322 -2041 -306
rect -17 -130 17 -114
rect -17 -322 17 -306
rect 2041 -130 2075 -114
rect 2041 -322 2075 -306
<< viali >>
rect -2013 294 -45 328
rect 45 294 2013 328
rect -2075 59 -2041 235
rect -17 59 17 235
rect 2041 59 2075 235
rect -2013 -71 -45 -37
rect 45 -71 2013 -37
rect -2075 -306 -2041 -130
rect -17 -306 17 -130
rect 2041 -306 2075 -130
<< metal1 >>
rect -2025 328 -33 334
rect -2025 294 -2013 328
rect -45 294 -33 328
rect -2025 288 -33 294
rect 33 328 2025 334
rect 33 294 45 328
rect 2013 294 2025 328
rect 33 288 2025 294
rect -2081 235 -2035 247
rect -2081 59 -2075 235
rect -2041 59 -2035 235
rect -2081 47 -2035 59
rect -23 235 23 247
rect -23 59 -17 235
rect 17 59 23 235
rect -23 47 23 59
rect 2035 235 2081 247
rect 2035 59 2041 235
rect 2075 59 2081 235
rect 2035 47 2081 59
rect -2025 -37 -33 -31
rect -2025 -71 -2013 -37
rect -45 -71 -33 -37
rect -2025 -77 -33 -71
rect 33 -37 2025 -31
rect 33 -71 45 -37
rect 2013 -71 2025 -37
rect 33 -77 2025 -71
rect -2081 -130 -2035 -118
rect -2081 -306 -2075 -130
rect -2041 -306 -2035 -130
rect -2081 -318 -2035 -306
rect -23 -130 23 -118
rect -23 -306 -17 -130
rect 17 -306 23 -130
rect -23 -318 23 -306
rect 2035 -130 2081 -118
rect 2035 -306 2041 -130
rect 2075 -306 2081 -130
rect 2035 -318 2081 -306
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 10 m 2 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
