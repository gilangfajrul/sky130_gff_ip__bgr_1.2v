magic
tech sky130A
magscale 1 2
timestamp 1716599695
<< nwell >>
rect 45 1386 95 1602
rect 4376 1512 4431 1562
rect 4381 1396 4431 1512
rect 13125 1511 13201 1563
rect 4381 1385 4443 1396
rect 4381 1346 4441 1385
rect 146 1269 4274 1321
rect 4380 1314 4432 1341
rect 4369 1262 4432 1314
rect 21725 981 21775 1033
rect 21725 931 21827 981
rect 21867 931 26111 981
rect 26061 848 26111 931
rect 45 599 4221 649
rect 4381 599 4431 694
rect 45 516 95 599
rect 4380 349 4432 448
<< viali >>
rect 140 1895 178 1929
rect 25978 1895 26016 1929
rect 140 -17 178 17
rect 25978 -17 26016 17
<< metal1 >>
rect 128 1929 190 1935
rect 128 1895 140 1929
rect 178 1895 190 1929
rect 128 1889 190 1895
rect 25966 1929 26028 1935
rect 25966 1895 25978 1929
rect 26016 1895 26028 1929
rect 25966 1889 26028 1895
rect 128 1721 178 1889
rect 4332 1678 4481 1728
rect 8673 1678 8822 1728
rect 13009 1678 13158 1728
rect 17342 1678 17491 1728
rect 21673 1678 21822 1728
rect 25978 1722 26028 1889
rect 45 1512 140 1562
rect 4336 1512 4431 1562
rect 45 1064 95 1512
rect 4381 1396 4431 1512
rect 4466 1511 4476 1563
rect 4552 1511 4562 1563
rect 8586 1511 8596 1563
rect 8672 1511 8682 1563
rect 8717 1512 8812 1562
rect 13008 1512 13103 1562
rect 8717 1396 8767 1512
rect 4381 1387 4476 1396
rect 4381 1346 4469 1387
rect 8672 1346 8767 1396
rect 8802 1345 8812 1397
rect 8888 1345 8898 1397
rect 12922 1345 12932 1397
rect 13008 1345 13018 1397
rect 13053 1396 13103 1512
rect 13138 1511 13148 1563
rect 13224 1511 13234 1563
rect 17258 1511 17268 1563
rect 17344 1511 17354 1563
rect 17389 1512 17484 1562
rect 21680 1512 21775 1562
rect 17389 1396 17439 1512
rect 13053 1346 13148 1396
rect 17344 1346 17439 1396
rect 17474 1345 17484 1397
rect 17560 1345 17570 1397
rect 21594 1345 21604 1397
rect 21680 1345 21690 1397
rect 21725 1396 21775 1512
rect 21810 1511 21820 1563
rect 21896 1511 21906 1563
rect 21725 1346 21820 1396
rect 130 1179 140 1231
rect 216 1179 226 1231
rect 4250 1179 4260 1231
rect 4336 1179 4346 1231
rect 4381 1180 4476 1230
rect 8672 1180 8767 1230
rect 4381 1064 4431 1180
rect 45 1014 140 1064
rect 4336 1014 4431 1064
rect 4466 1013 4476 1065
rect 4552 1013 4562 1065
rect 8586 1013 8596 1065
rect 8672 1013 8682 1065
rect 8717 1064 8767 1180
rect 8802 1179 8812 1231
rect 8888 1179 8898 1231
rect 12922 1179 12932 1231
rect 13008 1179 13018 1231
rect 13053 1180 13148 1230
rect 17344 1180 17439 1230
rect 13053 1064 13103 1180
rect 8717 1014 8812 1064
rect 13008 1014 13103 1064
rect 13138 1013 13148 1065
rect 13224 1013 13234 1065
rect 17258 1013 17268 1065
rect 17344 1013 17354 1065
rect 17389 1064 17439 1180
rect 17474 1179 17484 1231
rect 17560 1179 17570 1231
rect 21594 1179 21604 1231
rect 21680 1179 21690 1231
rect 21810 1179 21820 1231
rect 21896 1179 21906 1231
rect 17389 1014 17484 1064
rect 21680 1014 21775 1064
rect 21725 981 21775 1014
rect 21810 1013 21820 1065
rect 21896 1013 21906 1065
rect 25930 1013 25940 1065
rect 26016 1013 26026 1065
rect 21725 931 26111 981
rect 130 847 140 899
rect 216 847 226 899
rect 4250 847 4260 899
rect 4336 847 4346 899
rect 4381 848 4501 898
rect 8674 848 8769 898
rect 4250 681 4260 733
rect 4336 681 4346 733
rect 4381 649 4431 848
rect 4466 681 4476 733
rect 4552 681 4562 733
rect 8586 681 8596 733
rect 8672 681 8682 733
rect 8719 732 8769 848
rect 8802 847 8812 899
rect 8888 847 8898 899
rect 12922 847 12932 899
rect 13008 847 13018 899
rect 13053 848 13148 898
rect 17344 848 17439 898
rect 13053 732 13103 848
rect 8719 682 8814 732
rect 13008 682 13103 732
rect 13138 681 13148 733
rect 13224 681 13234 733
rect 17258 681 17268 733
rect 17344 681 17354 733
rect 17389 732 17439 848
rect 17474 847 17484 899
rect 17560 847 17570 899
rect 21594 847 21604 899
rect 21680 847 21690 899
rect 26061 898 26111 931
rect 21725 848 21820 898
rect 26016 848 26111 898
rect 21725 732 21775 848
rect 17389 682 17484 732
rect 21680 682 21775 732
rect 21810 681 21820 733
rect 21896 681 21906 733
rect 25930 681 25940 733
rect 26016 681 26026 733
rect 45 599 4431 649
rect 45 566 95 599
rect 45 516 140 566
rect 4336 516 4431 566
rect 130 349 140 401
rect 216 349 226 401
rect 4250 349 4260 401
rect 4336 349 4346 401
rect 4381 400 4431 516
rect 4466 515 4476 567
rect 4552 515 4562 567
rect 8586 515 8596 567
rect 8672 515 8682 567
rect 8717 516 8812 566
rect 13008 516 13103 566
rect 8717 400 8767 516
rect 4381 350 4476 400
rect 8672 350 8767 400
rect 8802 349 8812 401
rect 8888 349 8898 401
rect 12922 349 12932 401
rect 13008 349 13018 401
rect 13053 400 13103 516
rect 13138 515 13148 567
rect 13224 515 13234 567
rect 17258 515 17268 567
rect 17344 515 17354 567
rect 17389 516 17484 566
rect 21680 516 21775 566
rect 17389 400 17439 516
rect 13053 350 13148 400
rect 17344 350 17439 400
rect 17474 349 17484 401
rect 17560 349 17570 401
rect 21594 349 21604 401
rect 21680 349 21690 401
rect 21725 400 21775 516
rect 21725 350 21820 400
rect 4324 184 4473 234
rect 8678 184 8827 234
rect 13008 184 13157 234
rect 17334 184 17483 234
rect 21661 184 21810 234
rect 128 23 178 184
rect 25978 23 26028 189
rect 128 17 190 23
rect 128 -17 140 17
rect 178 -17 190 17
rect 128 -23 190 -17
rect 25966 17 26028 23
rect 25966 -17 25978 17
rect 26016 -17 26028 17
rect 25966 -23 26028 -17
<< via1 >>
rect 4476 1511 4552 1563
rect 8596 1511 8672 1563
rect 8812 1345 8888 1397
rect 12932 1345 13008 1397
rect 13148 1511 13224 1563
rect 17268 1511 17344 1563
rect 17484 1345 17560 1397
rect 21604 1345 21680 1397
rect 21820 1511 21896 1563
rect 140 1179 216 1231
rect 4260 1179 4336 1231
rect 4476 1013 4552 1065
rect 8596 1013 8672 1065
rect 8812 1179 8888 1231
rect 12932 1179 13008 1231
rect 13148 1013 13224 1065
rect 17268 1013 17344 1065
rect 17484 1179 17560 1231
rect 21604 1179 21680 1231
rect 21820 1179 21896 1231
rect 21820 1013 21896 1065
rect 25940 1013 26016 1065
rect 140 847 216 899
rect 4260 847 4336 899
rect 4260 681 4336 733
rect 4476 681 4552 733
rect 8596 681 8672 733
rect 8812 847 8888 899
rect 12932 847 13008 899
rect 13148 681 13224 733
rect 17268 681 17344 733
rect 17484 847 17560 899
rect 21604 847 21680 899
rect 21820 681 21896 733
rect 25940 681 26016 733
rect 140 349 216 401
rect 4260 349 4336 401
rect 4476 515 4552 567
rect 8596 515 8672 567
rect 8812 349 8888 401
rect 12932 349 13008 401
rect 13148 515 13224 567
rect 17268 515 17344 567
rect 17484 349 17560 401
rect 21604 349 21680 401
<< metal2 >>
rect 4476 1563 4552 1573
rect 4380 1511 4476 1563
rect 4380 1321 4432 1511
rect 4476 1501 4552 1511
rect 8596 1563 8672 1573
rect 13148 1563 13224 1573
rect 8672 1511 8768 1563
rect 8596 1501 8672 1511
rect 8716 1397 8768 1511
rect 13052 1511 13148 1563
rect 8812 1397 8888 1407
rect 8716 1345 8812 1397
rect 8812 1335 8888 1345
rect 12932 1397 13008 1407
rect 13052 1397 13104 1511
rect 13148 1501 13224 1511
rect 17268 1563 17344 1573
rect 21820 1563 21896 1573
rect 17344 1511 17440 1563
rect 17268 1501 17344 1511
rect 13008 1345 13104 1397
rect 17388 1397 17440 1511
rect 21724 1511 21820 1563
rect 17484 1397 17560 1407
rect 17388 1345 17484 1397
rect 12932 1335 13008 1345
rect 17484 1335 17560 1345
rect 21604 1397 21680 1407
rect 21724 1397 21776 1511
rect 21820 1501 21896 1511
rect 21680 1345 21776 1397
rect 21604 1335 21680 1345
rect 44 1269 4432 1321
rect 44 1231 96 1269
rect 140 1231 216 1241
rect 44 1179 140 1231
rect 140 1169 216 1179
rect 4260 1231 4336 1241
rect 8812 1231 8888 1241
rect 4336 1179 4432 1231
rect 4260 1169 4336 1179
rect 4380 1065 4432 1179
rect 8716 1179 8812 1231
rect 4476 1065 4552 1075
rect 4380 1013 4476 1065
rect 4476 1003 4552 1013
rect 8596 1065 8672 1075
rect 8716 1065 8768 1179
rect 8812 1169 8888 1179
rect 12932 1231 13008 1241
rect 17484 1231 17560 1241
rect 13008 1179 13104 1231
rect 12932 1169 13008 1179
rect 8672 1013 8768 1065
rect 13052 1065 13104 1179
rect 17388 1179 17484 1231
rect 13148 1065 13224 1075
rect 13052 1013 13148 1065
rect 8596 1003 8672 1013
rect 13148 1003 13224 1013
rect 17268 1065 17344 1075
rect 17388 1065 17440 1179
rect 17484 1169 17560 1179
rect 21604 1231 21680 1241
rect 21820 1233 21896 1243
rect 21680 1179 21776 1231
rect 21604 1169 21680 1179
rect 17344 1013 17440 1065
rect 21724 1065 21776 1179
rect 21820 1167 21896 1177
rect 21820 1065 21896 1075
rect 21724 1013 21820 1065
rect 17268 1003 17344 1013
rect 21820 1003 21896 1013
rect 25940 1065 26016 1075
rect 26016 1013 26112 1065
rect 25940 1003 26016 1013
rect 140 899 216 909
rect 44 847 140 899
rect 44 401 96 847
rect 140 837 216 847
rect 4260 899 4336 909
rect 8812 899 8888 909
rect 4336 847 4432 899
rect 4260 837 4336 847
rect 4260 735 4336 745
rect 4380 733 4432 847
rect 8716 847 8812 899
rect 4476 733 4552 743
rect 4380 681 4476 733
rect 4260 669 4336 679
rect 4476 671 4552 681
rect 8596 733 8672 743
rect 8716 733 8768 847
rect 8812 837 8888 847
rect 12932 899 13008 909
rect 17484 899 17560 909
rect 13008 847 13104 899
rect 12932 837 13008 847
rect 8672 681 8768 733
rect 13052 733 13104 847
rect 17388 847 17484 899
rect 13148 733 13224 743
rect 13052 681 13148 733
rect 8596 671 8672 681
rect 13148 671 13224 681
rect 17268 733 17344 743
rect 17388 733 17440 847
rect 17484 837 17560 847
rect 21604 899 21680 909
rect 21680 847 21776 899
rect 21604 837 21680 847
rect 17344 681 17440 733
rect 21724 733 21776 847
rect 21820 733 21896 743
rect 21724 681 21820 733
rect 17268 671 17344 681
rect 21820 671 21896 681
rect 25940 733 26016 743
rect 26060 733 26112 1013
rect 26016 681 26112 733
rect 25940 671 26016 681
rect 4476 567 4552 577
rect 4380 515 4476 567
rect 140 401 216 411
rect 44 349 140 401
rect 140 339 216 349
rect 4260 401 4336 411
rect 4380 401 4432 515
rect 4476 505 4552 515
rect 8596 567 8672 577
rect 13148 567 13224 577
rect 8672 515 8768 567
rect 8596 505 8672 515
rect 4336 349 4432 401
rect 8716 401 8768 515
rect 13052 515 13148 567
rect 8812 401 8888 411
rect 8716 349 8812 401
rect 4260 339 4336 349
rect 8812 339 8888 349
rect 12932 401 13008 411
rect 13052 401 13104 515
rect 13148 505 13224 515
rect 17268 567 17344 577
rect 17344 515 17440 567
rect 17268 505 17344 515
rect 13008 349 13104 401
rect 17388 401 17440 515
rect 17484 401 17560 411
rect 17388 349 17484 401
rect 12932 339 13008 349
rect 17484 339 17560 349
rect 21604 401 21680 411
rect 21604 339 21680 349
<< via2 >>
rect 21820 1231 21896 1233
rect 21820 1179 21896 1231
rect 21820 1177 21896 1179
rect 4260 733 4336 735
rect 4260 681 4336 733
rect 4260 679 4336 681
<< metal3 >>
rect 21717 1233 21906 1238
rect 21717 1177 21820 1233
rect 21896 1177 21906 1233
rect 21717 1172 21906 1177
rect 21717 989 21783 1172
rect 4373 923 21783 989
rect 4373 740 4439 923
rect 4250 735 4439 740
rect 4250 679 4260 735
rect 4336 679 4439 735
rect 4250 674 4439 679
use sky130_fd_pr__res_high_po_0p35_NUNB3Q  sky130_fd_pr__res_high_po_0p35_NUNB3Q_0
timestamp 1716568865
transform 0 -1 13078 1 0 956
box -1009 -13131 1009 13131
<< end >>
