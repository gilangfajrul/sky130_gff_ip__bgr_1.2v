magic
tech sky130A
magscale 1 2
timestamp 1717227652
<< nwell >>
rect 464 1614 2262 2520
<< nsubdiff >>
rect 500 2450 560 2484
rect 2166 2450 2226 2484
rect 500 2424 534 2450
rect 2192 2424 2226 2450
rect 500 1684 534 1710
rect 2192 1684 2226 1710
rect 500 1650 560 1684
rect 2166 1650 2226 1684
<< nsubdiffcont >>
rect 560 2450 2166 2484
rect 500 1710 534 2424
rect 2192 1710 2226 2424
rect 560 1650 2166 1684
<< poly >>
rect 646 2164 676 2196
rect 584 2148 676 2164
rect 584 2114 600 2148
rect 634 2114 676 2148
rect 584 2098 676 2114
rect 2050 2164 2080 2170
rect 2050 2148 2142 2164
rect 2050 2114 2092 2148
rect 2126 2114 2142 2148
rect 2050 2098 2142 2114
rect 2050 2040 2142 2056
rect 584 2020 676 2036
rect 584 1986 600 2020
rect 634 1986 676 2020
rect 584 1970 676 1986
rect 646 1938 676 1970
rect 2050 2006 2092 2040
rect 2126 2006 2142 2040
rect 2050 1990 2142 2006
rect 2050 1964 2081 1990
<< polycont >>
rect 600 2114 634 2148
rect 2092 2114 2126 2148
rect 600 1986 634 2020
rect 2092 2006 2126 2040
<< locali >>
rect 500 2450 560 2484
rect 2166 2450 2226 2484
rect 500 2424 534 2450
rect 2192 2424 2226 2450
rect 600 2148 634 2196
rect 600 2098 634 2114
rect 2092 2148 2126 2193
rect 2092 2098 2126 2114
rect 2092 2040 2126 2056
rect 600 2020 634 2036
rect 600 1938 634 1986
rect 2092 1939 2126 2006
rect 500 1684 534 1710
rect 2192 1684 2226 1710
rect 500 1650 560 1684
rect 2166 1650 2226 1684
<< viali >>
rect 1346 2450 1380 2484
rect 500 2114 534 2148
rect 600 2114 634 2148
rect 2092 2114 2126 2148
rect 2192 2114 2226 2148
rect 500 1986 534 2020
rect 600 1986 634 2020
rect 2092 2006 2126 2040
rect 2192 2006 2226 2040
rect 1346 1650 1380 1684
rect 1346 1649 1380 1650
<< metal1 >>
rect 1334 2484 1392 2490
rect 1334 2450 1346 2484
rect 1380 2450 1392 2484
rect 1334 2384 1392 2450
rect 1327 2208 1337 2384
rect 1389 2208 1399 2384
rect 1985 2208 1995 2384
rect 2047 2208 2057 2384
rect 594 2154 640 2196
rect 488 2148 640 2154
rect 488 2114 500 2148
rect 534 2114 600 2148
rect 634 2114 640 2148
rect 488 2108 640 2114
rect 594 2102 640 2108
rect 682 2090 728 2208
rect 2086 2154 2132 2207
rect 2086 2148 2238 2154
rect 880 2090 1188 2114
rect 1538 2090 1846 2115
rect 2086 2114 2092 2148
rect 2126 2114 2192 2148
rect 2226 2114 2238 2148
rect 2086 2108 2238 2114
rect 2086 2102 2132 2108
rect 682 2044 2044 2090
rect 594 2026 640 2032
rect 488 2020 640 2026
rect 880 2021 1188 2044
rect 1538 2022 1846 2044
rect 488 1986 500 2020
rect 534 1986 600 2020
rect 634 1986 640 2020
rect 488 1980 640 1986
rect 594 1938 640 1980
rect 1998 1931 2044 2044
rect 2086 2046 2132 2052
rect 2086 2040 2238 2046
rect 2086 2006 2092 2040
rect 2126 2006 2192 2040
rect 2226 2006 2238 2040
rect 2086 2000 2238 2006
rect 2086 1932 2132 2000
rect 669 1750 679 1926
rect 731 1750 741 1926
rect 1327 1750 1337 1926
rect 1389 1750 1399 1926
rect 1340 1684 1386 1750
rect 1340 1649 1346 1684
rect 1380 1649 1386 1684
rect 1340 1637 1386 1649
<< via1 >>
rect 1337 2208 1389 2384
rect 1995 2208 2047 2384
rect 679 1750 731 1926
rect 1337 1750 1389 1926
<< metal2 >>
rect 1335 2384 1391 2394
rect 1335 2198 1391 2208
rect 1995 2384 2047 2394
rect 1995 2093 2047 2208
rect 679 2041 2047 2093
rect 679 1926 731 2041
rect 679 1740 731 1750
rect 1335 1926 1391 1936
rect 1335 1740 1391 1750
<< via2 >>
rect 1335 2208 1337 2384
rect 1337 2208 1389 2384
rect 1389 2208 1391 2384
rect 1335 1750 1337 1926
rect 1337 1750 1389 1926
rect 1389 1750 1391 1926
<< metal3 >>
rect 1325 2384 1401 2389
rect 1325 2208 1335 2384
rect 1391 2208 1401 2384
rect 1325 2203 1401 2208
rect 1333 1931 1393 2203
rect 1325 1926 1401 1931
rect 1325 1750 1335 1926
rect 1391 1750 1401 1926
rect 1325 1745 1401 1750
use sky130_fd_pr__pfet_01v8_2XU96L  sky130_fd_pr__pfet_01v8_2XU96L_1 ~/chipalooza/sky130_gff_ip__bgr_1.2v/magic
timestamp 1717000582
transform 1 0 661 0 1 1838
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XU96L  sky130_fd_pr__pfet_01v8_2XU96L_2
timestamp 1717000582
transform 1 0 661 0 1 2296
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XU96L  sky130_fd_pr__pfet_01v8_2XU96L_3
timestamp 1717000582
transform 1 0 2065 0 1 2296
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XU96L  sky130_fd_pr__pfet_01v8_2XU96L_4
timestamp 1717000582
transform 1 0 2065 0 1 1838
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_9X8F2A  sky130_fd_pr__pfet_01v8_9X8F2A_0
timestamp 1717222322
transform 1 0 1363 0 1 1874
box -723 -198 723 164
use sky130_fd_pr__pfet_01v8_CVDFWD  sky130_fd_pr__pfet_01v8_CVDFWD_0
timestamp 1717222322
transform 1 0 1363 0 1 2260
box -723 -164 723 198
<< labels >>
flabel metal1 1353 2428 1353 2428 0 FreeSans 160 0 0 0 VDD
port 2 nsew
flabel metal2 2017 2125 2017 2125 0 FreeSans 160 0 0 0 D2
port 3 nsew
flabel metal1 2027 2000 2027 2000 0 FreeSans 160 0 0 0 D1
port 5 nsew
<< end >>
