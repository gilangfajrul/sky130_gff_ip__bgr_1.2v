magic
tech sky130A
magscale 1 2
timestamp 1718727926
<< dnwell >>
rect -18177 13834 9526 23101
rect -18177 -28 -1264 13834
rect 8926 -27 9526 13834
rect 0 -28 9526 -27
rect -18177 -628 9526 -28
<< nwell >>
rect -18257 22896 9606 23182
rect -18257 -422 -17971 22896
rect -16702 14626 -2985 17677
rect 9320 -422 9606 22896
rect -18257 -708 9606 -422
<< pwell >>
rect -1450 14508 8723 17815
<< nsubdiff >>
rect -18220 23125 9569 23145
rect -18220 23091 -18140 23125
rect 9489 23091 9569 23125
rect -18220 23071 9569 23091
rect -18220 23065 -18146 23071
rect -18220 -591 -18200 23065
rect -18166 -591 -18146 23065
rect -18220 -597 -18146 -591
rect 9495 23065 9569 23071
rect 9495 -591 9515 23065
rect 9549 -591 9569 23065
rect 9495 -597 9569 -591
rect -18220 -617 9569 -597
rect -18220 -651 -18140 -617
rect 9489 -651 9569 -617
rect -18220 -671 9569 -651
<< nsubdiffcont >>
rect -18140 23091 9489 23125
rect -18200 -591 -18166 23065
rect 9515 -591 9549 23065
rect -18140 -651 9489 -617
<< locali >>
rect -18200 23091 -18140 23125
rect 9489 23091 9549 23125
rect -18200 23065 -18166 23091
rect 9515 23065 9549 23091
rect -18200 -617 -18166 -591
rect 9515 -617 9549 -591
rect -18200 -651 -18140 -617
rect 9489 -651 9549 -617
<< viali >>
rect -17337 20867 -16940 20901
rect -12825 19303 -12600 19337
rect -14371 15664 -7986 15698
rect -7585 15658 -5316 15692
rect -10222 15558 -7986 15592
rect -5650 15552 -5281 15586
rect -7960 15110 -7926 15459
rect -7577 15131 -7543 15480
<< metal1 >>
rect -17347 22334 -17337 22386
rect -16940 22334 -16930 22386
rect -17582 22169 -16928 22219
rect -17582 20757 -17532 22169
rect -3 22002 7 22054
rect 404 22002 414 22054
rect 4333 21836 4343 21888
rect 4740 21836 4750 21888
rect -17365 21329 -17355 21399
rect -16923 21329 -16913 21399
rect -17312 21166 -17302 21231
rect -17118 21166 -17108 21231
rect -17161 21165 -17118 21166
rect -17347 21024 -17337 21058
rect -17349 21006 -17337 21024
rect -16940 21024 -16930 21058
rect -16940 21006 -16928 21024
rect -17349 20901 -16928 21006
rect -17349 20867 -17337 20901
rect -16940 20867 -16928 20901
rect -17349 20861 -16928 20867
rect -17582 20707 -13228 20757
rect -13278 17800 -13228 20707
rect -13011 20440 -12592 20655
rect -13150 19598 -12592 19670
rect -13150 19209 -13078 19598
rect -13011 19442 -13001 19494
rect -12604 19491 -12594 19494
rect -12604 19442 -12588 19491
rect -12836 19343 -12588 19442
rect -12837 19337 -12588 19343
rect -12837 19303 -12825 19337
rect -12600 19303 -12588 19337
rect -12837 19297 -12588 19303
rect -13150 19137 -7820 19209
rect -16774 17750 -13228 17800
rect -16774 17069 -16724 17750
rect -16774 17019 -16389 17069
rect -16435 16745 -16389 17019
rect -8353 15704 -7938 15705
rect -14383 15698 -7938 15704
rect -14383 15664 -14371 15698
rect -7986 15664 -7938 15698
rect -14383 15658 -7938 15664
rect -17911 15546 -12226 15619
rect -8353 15598 -7938 15658
rect -10234 15592 -7938 15598
rect -10234 15558 -10222 15592
rect -7986 15558 -7938 15592
rect -10234 15552 -7938 15558
rect -12286 15171 -12240 15546
rect -11736 15462 -11726 15514
rect -10742 15462 -10732 15514
rect -9678 15462 -9668 15514
rect -8684 15462 -8674 15514
rect -8353 15492 -7938 15552
rect -7892 15618 -7820 19137
rect -7770 18045 -7544 18111
rect -7770 17226 -7704 18045
rect -2235 17322 -2110 17841
rect -7780 17160 -7770 17226
rect -7704 17160 -7694 17226
rect -2245 17197 -2235 17322
rect -2110 17197 -2100 17322
rect 39 17269 99 17293
rect 31 17262 99 17269
rect -2235 17191 -2110 17197
rect -1450 17171 -1059 17223
rect 39 17209 99 17262
rect -7723 16989 -7717 17049
rect -7657 16989 -2858 17049
rect -3305 16784 -3245 16989
rect -3305 16218 -3245 16458
rect -2918 16308 -2858 16989
rect -2390 16608 -2338 16614
rect -1450 16608 -1398 17171
rect -303 17149 99 17209
rect -990 16609 -944 16873
rect -2338 16556 -1398 16608
rect -993 16603 -941 16609
rect -2390 16550 -2338 16556
rect -1003 16551 -993 16603
rect -941 16551 -931 16603
rect -993 16545 -941 16551
rect -303 16396 -243 17149
rect -2745 16336 -2739 16396
rect -2679 16336 -243 16396
rect -2918 16248 -247 16308
rect -3305 16158 -342 16218
rect -402 15872 -342 16158
rect -307 15960 -247 16248
rect 8530 16158 8576 16531
rect 8535 15992 8787 16061
rect -307 15900 4073 15960
rect -402 15812 3934 15872
rect -7595 15698 -7585 15701
rect -7597 15652 -7585 15698
rect -7236 15698 -7226 15701
rect -5650 15698 -5269 15699
rect -7236 15692 -5269 15698
rect -5316 15658 -5269 15692
rect -7595 15649 -7585 15652
rect -7236 15652 -5269 15658
rect -7236 15649 -7226 15652
rect -7892 15546 -7334 15618
rect -5662 15586 -5269 15652
rect -2394 15603 -2334 15609
rect -5662 15552 -5650 15586
rect -5281 15552 -5269 15586
rect -5662 15546 -5269 15552
rect -8353 15480 -7537 15492
rect -8353 15473 -7586 15480
rect -7966 15459 -7586 15473
rect -7966 15110 -7960 15459
rect -7926 15131 -7586 15459
rect -7534 15131 -7524 15480
rect -7380 15464 -7334 15546
rect -3271 15543 -2394 15603
rect -3271 15283 -3211 15543
rect -2394 15537 -2334 15543
rect 3874 15381 3934 15812
rect 4013 15523 4073 15900
rect 8369 15874 8379 15934
rect 8439 15874 8449 15934
rect 8369 15767 8449 15874
rect 4878 15670 4888 15722
rect 5872 15670 5882 15722
rect 6936 15670 6946 15722
rect 7930 15670 7940 15722
rect 8694 15635 8787 15992
rect 8550 15567 8787 15635
rect 8550 15566 8763 15567
rect 4003 15463 4013 15523
rect 4073 15463 4083 15523
rect 3868 15329 3878 15381
rect 3930 15329 3940 15381
rect 2982 15242 3155 15323
rect 3235 15242 3245 15323
rect -7926 15110 -7537 15131
rect -994 15112 -934 15118
rect -7966 15098 -7537 15110
rect -7926 14626 -7586 15098
rect -2641 15052 -994 15112
rect -934 15052 -924 15112
rect 3610 15102 4274 15268
rect -7387 14645 -7327 15013
rect -2641 14645 -2581 15052
rect -994 15046 -934 15052
rect -376 15009 -48 15059
rect -2234 14929 -2109 14935
rect -2244 14804 -2234 14929
rect -2109 14804 -893 14929
rect -2234 14798 -2109 14804
rect -8047 13355 -7469 14626
rect -7387 14585 -2581 14645
rect -1018 14170 -893 14804
rect -375 14526 -325 15009
rect 3610 14951 3776 15102
rect 2924 14935 3776 14951
rect 2924 14819 3018 14935
rect 3161 14819 3776 14935
rect 2924 14785 3776 14819
rect -376 14520 -324 14526
rect -376 14462 -324 14468
rect -1018 14039 -893 14045
rect -8047 12777 4635 13355
rect 5213 12777 5219 13355
rect 397 11390 407 12166
rect 459 11390 469 12166
rect 4507 12162 4579 12168
rect 4042 12100 4052 12152
rect 4228 12100 4238 12152
rect 4579 12090 9169 12162
rect 4507 12084 4579 12090
rect 4042 11842 4052 11894
rect 4228 11842 4238 11894
rect 4628 11713 4638 11765
rect 5208 11713 5218 11765
rect 5606 11634 9204 11680
rect 5606 11298 5652 11634
rect 4272 11227 4428 11273
rect 5261 11252 5652 11298
rect 397 10396 407 11172
rect 459 10396 469 11172
rect 4042 10668 4052 10720
rect 4228 10668 4238 10720
rect 4042 10410 4052 10462
rect 4228 10410 4238 10462
rect 4205 10350 4322 10361
rect 786 9200 852 10345
rect 1678 9346 1744 10340
rect 2567 9462 2633 10342
rect 3481 9585 3547 10326
rect 4205 9787 4324 10350
rect 4382 9939 4428 11227
rect 4814 10373 5032 10757
rect 4814 10155 9201 10373
rect 4382 9893 9196 9939
rect 4205 9668 9196 9787
rect 3481 9519 9186 9585
rect 2567 9396 9186 9462
rect 1678 9280 9184 9346
rect 786 9134 9184 9200
rect 2011 6034 2021 6715
rect 2701 6034 2711 6715
rect 623 1870 633 2550
rect 1313 1870 1323 2550
<< via1 >>
rect -17337 22334 -16940 22386
rect 7 22002 404 22054
rect 4343 21836 4740 21888
rect -17355 21329 -16923 21399
rect -17302 21166 -17118 21231
rect -17337 21006 -16940 21058
rect -13001 19442 -12604 19494
rect -11726 15462 -10742 15514
rect -9668 15462 -8684 15514
rect -7770 17160 -7704 17226
rect -2235 17197 -2110 17322
rect -7717 16989 -7657 17049
rect -2390 16556 -2338 16608
rect -993 16551 -941 16603
rect -2739 16336 -2679 16396
rect -7585 15692 -7236 15701
rect -7585 15658 -7236 15692
rect -7585 15649 -7236 15658
rect -7586 15131 -7577 15480
rect -7577 15131 -7543 15480
rect -7543 15131 -7534 15480
rect -2394 15543 -2334 15603
rect 8379 15874 8439 15934
rect 4888 15670 5872 15722
rect 6946 15670 7930 15722
rect 4013 15463 4073 15523
rect 3878 15329 3930 15381
rect 3155 15242 3235 15323
rect -994 15052 -934 15112
rect -2234 14804 -2109 14929
rect 3018 14819 3161 14935
rect -376 14468 -324 14520
rect -1018 14045 -893 14170
rect 4635 12777 5213 13355
rect 407 11390 459 12166
rect 4052 12100 4228 12152
rect 4507 12090 4579 12162
rect 4052 11842 4228 11894
rect 4638 11713 5208 11765
rect 407 10396 459 11172
rect 4052 10668 4228 10720
rect 4052 10410 4228 10462
rect 2021 6034 2701 6715
rect 633 1870 1313 2550
<< metal2 >>
rect -17337 22388 -16940 22398
rect -17337 22322 -16940 22332
rect 7 22054 404 22064
rect 7 21992 404 22002
rect -368 21836 -145 21888
rect -8683 21668 -8673 21724
rect -8617 21668 -8607 21724
rect -17573 21399 -16923 21409
rect -17573 21329 -17355 21399
rect -17573 21319 -16923 21329
rect -17573 20863 -17439 21319
rect -17302 21231 -17118 21241
rect -17302 21156 -17118 21166
rect -17337 21060 -16940 21070
rect -17337 20994 -16940 21004
rect -17573 20729 -13166 20863
rect -13300 19358 -13166 20729
rect -13001 19496 -12604 19506
rect -13001 19430 -12604 19440
rect -13300 19224 -7680 19358
rect -368 19320 -302 21836
rect 332 19443 404 21992
rect 4343 21888 4740 21898
rect 4343 21826 4740 21836
rect 4668 19610 4740 21826
rect 4668 19538 8636 19610
rect 8708 19538 8717 19610
rect 8497 19443 8569 19453
rect 332 19371 8497 19443
rect 8569 19371 8578 19443
rect 8497 19361 8569 19371
rect 8313 19320 8369 19325
rect -368 19315 8374 19320
rect -368 19259 8313 19315
rect 8369 19259 8378 19315
rect -368 19254 8374 19259
rect 8313 19249 8369 19254
rect -8041 17772 -8027 17838
rect -7961 17772 -7947 17838
rect -8041 17523 -7947 17772
rect -8041 17467 -8022 17523
rect -7966 17467 -7947 17523
rect -7814 17645 -7680 19224
rect -7814 17526 -1288 17645
rect -7814 17511 -1417 17526
rect -8041 17447 -7947 17467
rect -1422 17402 -1417 17511
rect -1293 17402 -1288 17526
rect -1422 17397 -1288 17402
rect -1417 17393 -1293 17397
rect -2235 17322 -2110 17332
rect -7770 17226 -7704 17236
rect -2241 17197 -2235 17322
rect -2110 17197 -2104 17322
rect -2235 17187 -2110 17197
rect -7770 17150 -7704 17160
rect 41 17058 97 17068
rect -7717 17049 -7657 17055
rect -8011 16989 -7717 17049
rect -12324 16975 -12268 16985
rect -7717 16983 -7657 16989
rect 41 16872 97 16882
rect -12324 16789 -12268 16799
rect -2394 16612 -2334 16621
rect -996 16612 -932 16622
rect -2396 16556 -2394 16608
rect -2334 16556 -2332 16608
rect -2394 16543 -2334 16552
rect -1006 16547 -997 16607
rect -932 16547 -928 16607
rect -996 16532 -932 16542
rect -3105 16434 -142 16494
rect -2739 16396 -2679 16406
rect -2739 16326 -2679 16336
rect 4157 15914 4209 16280
rect 8379 15934 8439 15944
rect -1198 15866 -1132 15871
rect -1935 15861 -1132 15866
rect -10241 15524 -10169 15797
rect -1935 15795 -1920 15861
rect -1854 15795 -1198 15861
rect -1935 15790 -1132 15795
rect -1198 15785 -1132 15790
rect 1425 15862 4209 15914
rect 8372 15876 8379 15932
rect 8439 15876 8446 15932
rect 8379 15864 8439 15874
rect -7586 15701 -7236 15711
rect -7586 15649 -7585 15701
rect -7586 15543 -7236 15649
rect 1425 15610 1477 15862
rect 4888 15724 5872 15734
rect 4888 15658 5872 15668
rect 6946 15724 7930 15734
rect 6946 15658 7930 15668
rect -2400 15601 -2394 15603
rect -2334 15601 -2328 15603
rect -2401 15545 -2394 15601
rect -2334 15545 -2327 15601
rect -2400 15543 -2394 15545
rect -2334 15543 -2328 15545
rect -11726 15514 -8684 15524
rect -10742 15462 -9668 15514
rect -11726 15452 -8684 15462
rect -7586 15480 -7467 15543
rect -7534 15131 -7467 15480
rect 3154 15523 4073 15533
rect 3154 15463 4013 15523
rect 3154 15453 4073 15463
rect 3154 15333 3234 15453
rect 3874 15385 3934 15395
rect 3154 15330 3235 15333
rect 3155 15323 3235 15330
rect 3874 15315 3934 15325
rect 3155 15232 3235 15242
rect -7586 15121 -7534 15131
rect -996 15114 -932 15124
rect -1000 15052 -996 15112
rect -932 15052 -928 15112
rect -996 15040 -932 15050
rect 1425 14976 1477 15065
rect 1425 14945 3160 14976
rect -2234 14929 -2109 14939
rect 1425 14935 3161 14945
rect 1425 14924 3018 14935
rect 3018 14809 3161 14819
rect -2234 14794 -2109 14804
rect -2526 14664 1356 14674
rect -2526 14659 1285 14664
rect -2526 14603 -2518 14659
rect -2462 14603 1285 14659
rect -2526 14598 1285 14603
rect 1351 14598 1356 14664
rect -2526 14588 1356 14598
rect 4306 14584 4376 14593
rect 3774 14583 4377 14584
rect -1446 14520 -318 14521
rect -1446 14468 -376 14520
rect -324 14468 -318 14520
rect -1446 14461 -318 14468
rect 3774 14513 4306 14583
rect 4376 14513 4377 14583
rect 3774 14512 4377 14513
rect -1446 7351 -1386 14461
rect -1024 14045 -1018 14170
rect -893 14045 -887 14170
rect 405 14110 461 14119
rect 402 14054 405 14057
rect 461 14054 464 14057
rect -1018 9475 -893 14045
rect 402 12166 464 14054
rect 402 11390 407 12166
rect 459 11390 464 12166
rect 402 11172 464 11390
rect 402 10396 407 11172
rect 459 10396 464 11172
rect 402 10384 464 10396
rect 655 12873 727 12883
rect 655 10386 727 12801
rect 1547 12849 1619 12859
rect 2439 12842 2511 12847
rect 2435 12780 2444 12842
rect 2506 12780 2515 12842
rect 1547 10396 1619 12777
rect 2439 10396 2511 12780
rect 2262 9476 2458 9491
rect 3304 9476 3429 12166
rect 3774 10730 3846 14512
rect 4306 14503 4376 14512
rect 4754 14447 4816 14451
rect 3904 14442 4821 14447
rect 3904 14380 4754 14442
rect 4816 14380 4821 14442
rect 3904 14375 4821 14380
rect 3904 11904 3976 14375
rect 4754 14371 4816 14375
rect 4635 13355 5213 13361
rect 4052 12152 4507 12162
rect 4228 12100 4507 12152
rect 4052 12090 4507 12100
rect 4579 12090 4585 12162
rect 3904 11894 4240 11904
rect 3904 11842 4052 11894
rect 4228 11842 4240 11894
rect 3904 11832 4240 11842
rect 4635 11765 5213 12777
rect 4635 11755 4638 11765
rect 5208 11755 5213 11765
rect 4638 11703 5208 11713
rect 4627 11019 9178 11539
rect 5787 10892 9204 10964
rect 3774 10720 4240 10730
rect 3774 10668 4052 10720
rect 4228 10668 4240 10720
rect 3774 10658 4240 10668
rect 5787 10472 5859 10892
rect 4052 10462 5859 10472
rect 4228 10410 5859 10462
rect 4052 10400 5859 10410
rect 2262 9475 3429 9476
rect -1018 9351 3429 9475
rect -1018 9350 2458 9351
rect 2262 9335 2458 9350
rect -1446 7282 -1386 7291
rect 2291 6725 2416 9335
rect 3679 9024 3803 9033
rect 3679 8740 3803 8900
rect 2021 6715 2701 6725
rect 2021 6024 2701 6034
rect 633 2550 1313 2560
rect 633 1860 1313 1870
<< via2 >>
rect -17337 22386 -16940 22388
rect -17337 22334 -16940 22386
rect -17337 22332 -16940 22334
rect -8673 21668 -8617 21724
rect -17298 21170 -17122 21226
rect -17337 21058 -16940 21060
rect -17337 21006 -16940 21058
rect -17337 21004 -16940 21006
rect -13001 19494 -12604 19496
rect -13001 19442 -12604 19494
rect -13001 19440 -12604 19442
rect 8636 19538 8708 19610
rect 8497 19371 8569 19443
rect 8313 19259 8369 19315
rect -8027 17772 -7961 17838
rect -8022 17467 -7966 17523
rect -1417 17402 -1293 17526
rect -7770 17160 -7704 17226
rect -2235 17197 -2110 17322
rect -12324 16799 -12268 16975
rect 41 16882 97 17058
rect -2394 16608 -2334 16612
rect -2394 16556 -2390 16608
rect -2390 16556 -2338 16608
rect -2338 16556 -2334 16608
rect -996 16607 -932 16612
rect -2394 16552 -2334 16556
rect -997 16603 -932 16607
rect -997 16551 -993 16603
rect -993 16551 -941 16603
rect -941 16551 -932 16603
rect -997 16547 -932 16551
rect -996 16542 -932 16547
rect -2739 16336 -2679 16396
rect -1920 15795 -1854 15861
rect -1198 15795 -1132 15861
rect 8381 15876 8437 15932
rect 4888 15722 5872 15724
rect 4888 15670 5872 15722
rect 4888 15668 5872 15670
rect 6946 15722 7930 15724
rect 6946 15670 7930 15722
rect 6946 15668 7930 15670
rect -2392 15545 -2336 15601
rect 4013 15463 4073 15523
rect 3874 15381 3934 15385
rect 3874 15329 3878 15381
rect 3878 15329 3930 15381
rect 3930 15329 3934 15381
rect 3874 15325 3934 15329
rect -996 15112 -932 15114
rect -996 15052 -994 15112
rect -994 15052 -934 15112
rect -934 15052 -932 15112
rect -996 15050 -932 15052
rect -2229 14809 -2114 14924
rect -2518 14603 -2462 14659
rect 1285 14598 1351 14664
rect 4306 14513 4376 14583
rect 405 14054 461 14110
rect 655 12801 727 12873
rect 1547 12777 1619 12849
rect 2444 12780 2506 12842
rect 4754 14380 4816 14442
rect -1446 7291 -1386 7351
rect 3679 8900 3803 9024
rect 633 1870 1313 2550
<< metal3 >>
rect -17957 22388 -16930 22393
rect -17957 22332 -17337 22388
rect -16940 22332 -16930 22388
rect -17957 22327 -16930 22332
rect -17957 22311 -17506 22327
rect -17582 20785 -17506 22311
rect -8678 21724 -8612 21734
rect -8678 21668 -8673 21724
rect -8617 21668 -8612 21724
rect -8678 21646 -8612 21668
rect -17433 21580 -8612 21646
rect -17433 21230 -17368 21580
rect -17308 21230 -17112 21231
rect -17433 21226 -17112 21230
rect -17433 21170 -17298 21226
rect -17122 21170 -17112 21226
rect -17433 21165 -17112 21170
rect -17347 21064 -16930 21065
rect -17347 21000 -17337 21064
rect -16940 21000 -16930 21064
rect -17347 20999 -16930 21000
rect -17582 20709 -13258 20785
rect -13334 19222 -13258 20709
rect -13011 19500 -12594 19501
rect -13011 19436 -13001 19500
rect -12604 19436 -12594 19500
rect -13011 19435 -12594 19436
rect -8782 19271 -8688 21580
rect 8603 19615 8723 19623
rect 8603 19533 8631 19615
rect 8713 19533 8723 19615
rect 8603 19526 8723 19533
rect 8471 19443 8591 19453
rect 8471 19438 8497 19443
rect 8569 19438 8591 19443
rect 8471 19366 8492 19438
rect 8574 19366 8591 19438
rect 8471 19356 8591 19366
rect 8285 19319 8397 19331
rect -13334 19146 -12258 19222
rect -8782 19177 -7947 19271
rect 8285 19255 8309 19319
rect 8373 19255 8397 19319
rect 8285 19243 8397 19255
rect -12334 16975 -12258 19146
rect -8041 17838 -7947 19177
rect -8041 17772 -8027 17838
rect -7961 17772 -7947 17838
rect -8041 17767 -7947 17772
rect -8212 17602 -187 17666
rect 3478 17650 3560 17835
rect -8212 17158 -8148 17602
rect -8041 17523 -1841 17541
rect -8041 17467 -8022 17523
rect -7966 17467 -1841 17523
rect -8041 17447 -1841 17467
rect -2240 17322 -2105 17327
rect -7780 17226 -7694 17231
rect -7780 17160 -7770 17226
rect -7704 17160 -7694 17226
rect -2240 17197 -2235 17322
rect -2110 17197 -2105 17322
rect -2240 17192 -2105 17197
rect -7780 17155 -7694 17160
rect -12334 16799 -12324 16975
rect -12268 16799 -12258 16975
rect -12334 16794 -12258 16799
rect -7770 14664 -7704 17155
rect -2399 16612 -2329 16617
rect -2399 16552 -2394 16612
rect -2334 16552 -2329 16612
rect -2399 16547 -2329 16552
rect -2749 16396 -2669 16401
rect -3118 16336 -2739 16396
rect -2679 16336 -2669 16396
rect -2749 16331 -2669 16336
rect -2394 15606 -2334 16547
rect -2397 15601 -2331 15606
rect -2397 15545 -2392 15601
rect -2336 15545 -2331 15601
rect -2397 15540 -2331 15545
rect -2234 14929 -2109 17192
rect -1935 15861 -1841 17447
rect -1935 15795 -1920 15861
rect -1854 15795 -1841 15861
rect -1935 15790 -1841 15795
rect -2239 14924 -2104 14929
rect -2239 14809 -2229 14924
rect -2114 14809 -2104 14924
rect -2239 14804 -2104 14809
rect -7770 14659 -2452 14664
rect -7770 14603 -2518 14659
rect -2462 14603 -2452 14659
rect -7770 14598 -2452 14603
rect -1682 9067 -1586 17602
rect -1682 8973 -1681 9067
rect -1587 8973 -1586 9067
rect -1682 8972 -1586 8973
rect -1422 17526 -1288 17531
rect -1422 17402 -1417 17526
rect -1293 17402 -1288 17526
rect -1422 16002 -1288 17402
rect -251 17184 -187 17602
rect 3468 17568 3478 17650
rect 3560 17568 3570 17650
rect -251 17120 107 17184
rect 31 17058 107 17120
rect 31 16882 41 17058
rect 97 16882 107 17058
rect 31 16877 107 16882
rect -1019 16612 -909 16629
rect -1019 16607 -996 16612
rect -1019 16547 -997 16607
rect -1019 16542 -996 16547
rect -932 16542 -909 16612
rect -1019 16527 -909 16542
rect -1422 15927 6516 16002
rect 8379 15937 8439 16827
rect 8636 16112 8708 16113
rect 8631 16042 8637 16112
rect 8707 16042 8713 16112
rect -1422 9029 -1288 15927
rect -1198 15866 4878 15867
rect -1208 15861 4878 15866
rect -1208 15795 -1198 15861
rect -1132 15795 4878 15861
rect -1208 15790 4878 15795
rect 4801 15729 4878 15790
rect 6441 15729 6516 15927
rect 8376 15932 8442 15937
rect 8376 15876 8381 15932
rect 8437 15876 8442 15932
rect 8376 15871 8442 15876
rect 4801 15724 5882 15729
rect 4801 15668 4888 15724
rect 5872 15668 5882 15724
rect 4801 15663 5882 15668
rect 6441 15724 7940 15729
rect 6441 15668 6946 15724
rect 7930 15668 7940 15724
rect 6441 15664 7940 15668
rect 6881 15663 7940 15664
rect 4003 15523 4083 15528
rect 4003 15463 4013 15523
rect 4073 15463 4348 15523
rect 4003 15458 4083 15463
rect 3850 15390 3958 15403
rect 3850 15320 3869 15390
rect 3939 15320 3958 15390
rect 3850 15307 3958 15320
rect -1019 15114 -910 15131
rect -1019 15050 -996 15114
rect -932 15050 -910 15114
rect -1019 15027 -910 15050
rect 1280 14664 2512 14669
rect 1280 14598 1285 14664
rect 1351 14598 2512 14664
rect 1280 14593 2512 14598
rect 1745 14115 1809 14120
rect 400 14114 1810 14115
rect 400 14110 1745 14114
rect 400 14054 405 14110
rect 461 14054 1745 14110
rect 400 14050 1745 14054
rect 1809 14050 1810 14114
rect 400 14049 1810 14050
rect 1745 14044 1809 14049
rect 628 12878 754 12891
rect 628 12796 650 12878
rect 732 12796 754 12878
rect 628 12783 754 12796
rect 1521 12854 1645 12866
rect 1521 12772 1542 12854
rect 1624 12772 1645 12854
rect 2439 12842 2511 14593
rect 4284 14583 4397 14599
rect 4284 14513 4306 14583
rect 4376 14513 4397 14583
rect 4284 14497 4397 14513
rect 8636 14447 8708 16042
rect 4749 14442 8708 14447
rect 4749 14380 4754 14442
rect 4816 14380 8708 14442
rect 4749 14375 8708 14380
rect 2439 12780 2444 12842
rect 2506 12780 2511 12842
rect 2439 12775 2511 12780
rect 1521 12759 1645 12772
rect -1422 9024 3808 9029
rect -1681 8967 -1587 8972
rect -1422 8900 3679 9024
rect 3803 8900 3808 9024
rect -1422 8895 3808 8900
rect -1470 7356 -1362 7366
rect -1470 7286 -1451 7356
rect -1381 7286 -1362 7356
rect -1470 7275 -1362 7286
rect 623 2550 1323 2555
rect 623 1870 633 2550
rect 1313 1870 1323 2550
rect 623 1865 1323 1870
<< via3 >>
rect -17337 21060 -16940 21064
rect -17337 21004 -16940 21060
rect -17337 21000 -16940 21004
rect -13001 19496 -12604 19500
rect -13001 19440 -12604 19496
rect -13001 19436 -12604 19440
rect 8631 19610 8713 19615
rect 8631 19538 8636 19610
rect 8636 19538 8708 19610
rect 8708 19538 8713 19610
rect 8631 19533 8713 19538
rect 8492 19371 8497 19438
rect 8497 19371 8569 19438
rect 8569 19371 8574 19438
rect 8492 19366 8574 19371
rect 8309 19315 8373 19319
rect 8309 19259 8313 19315
rect 8313 19259 8369 19315
rect 8369 19259 8373 19315
rect 8309 19255 8373 19259
rect -1681 8973 -1587 9067
rect 3478 17568 3560 17650
rect -996 16542 -932 16612
rect 8637 16042 8707 16112
rect 3869 15385 3939 15390
rect 3869 15325 3874 15385
rect 3874 15325 3934 15385
rect 3934 15325 3939 15385
rect 3869 15320 3939 15325
rect -996 15050 -932 15114
rect 1745 14050 1809 14114
rect 650 12873 732 12878
rect 650 12801 655 12873
rect 655 12801 727 12873
rect 727 12801 732 12873
rect 650 12796 732 12801
rect 1542 12849 1624 12854
rect 1542 12777 1547 12849
rect 1547 12777 1619 12849
rect 1619 12777 1624 12849
rect 1542 12772 1624 12777
rect 4306 14513 4376 14583
rect -1451 7351 -1381 7356
rect -1451 7291 -1446 7351
rect -1446 7291 -1386 7351
rect -1386 7291 -1381 7351
rect -1451 7286 -1381 7291
rect 633 1870 1313 2550
<< metal4 >>
rect -17338 21064 -16939 21065
rect -17338 21000 -17337 21064
rect -16940 21000 -16939 21064
rect -17338 20999 -16939 21000
rect -17054 20907 -16940 20999
rect -17054 20793 -13226 20907
rect -13340 19387 -13226 20793
rect 8630 19615 8714 19616
rect 8630 19533 8631 19615
rect 8713 19533 8714 19615
rect 8630 19532 8714 19533
rect -13002 19500 -12603 19501
rect -13002 19499 -13001 19500
rect -13028 19436 -13001 19499
rect -12604 19436 -12603 19500
rect -13028 19435 -12603 19436
rect 8491 19438 8575 19439
rect -13028 19387 -12914 19435
rect -13340 19273 -12914 19387
rect 8491 19366 8492 19438
rect 8574 19366 8575 19438
rect 8491 19365 8575 19366
rect 8308 19319 8374 19320
rect -13340 17916 -13226 19273
rect 8308 19255 8309 19319
rect 8373 19255 8374 19319
rect -17736 17802 -13226 17916
rect -7760 19116 -5020 19182
rect -17736 15344 -16724 17802
rect -7760 17721 -7694 19116
rect 8308 18138 8374 19255
rect -7760 17655 -1487 17721
rect -17736 14332 -15401 15344
rect -16413 2198 -15401 14332
rect -1553 14318 -1487 17655
rect 3477 17650 3561 17651
rect 3477 17568 3478 17650
rect 3560 17568 3561 17650
rect -997 16612 -931 16613
rect -997 16542 -996 16612
rect -932 16542 -931 16612
rect -997 16541 -931 16542
rect -994 15115 -934 16541
rect -997 15114 -931 15115
rect -997 15050 -996 15114
rect -932 15050 -931 15114
rect -997 15049 -931 15050
rect 3477 14542 3561 17568
rect 1547 14470 3561 14542
rect -1553 14252 727 14318
rect -15226 12214 -1917 13224
rect 655 12879 727 14252
rect 649 12878 733 12879
rect 649 12796 650 12878
rect 732 12796 733 12878
rect 1547 12855 1619 14470
rect 3653 14115 3719 17854
rect 8497 15924 8569 19365
rect 8636 16112 8708 19532
rect 8636 16042 8637 16112
rect 8707 16042 8708 16112
rect 8636 16041 8708 16042
rect 8497 15852 8633 15924
rect 3868 15390 3940 15391
rect 3868 15320 3869 15390
rect 3939 15385 3940 15390
rect 3939 15325 4384 15385
rect 3939 15320 3940 15325
rect 3868 15319 3940 15320
rect 8561 14584 8633 15852
rect 4305 14583 8633 14584
rect 4305 14513 4306 14583
rect 4376 14513 8633 14583
rect 4305 14512 8633 14513
rect 1744 14114 3719 14115
rect 1744 14050 1745 14114
rect 1809 14050 3719 14114
rect 1744 14049 3719 14050
rect 649 12795 733 12796
rect 1541 12854 1625 12855
rect 1541 12772 1542 12854
rect 1624 12772 1625 12854
rect 1541 12771 1625 12772
rect -1830 9067 -1586 9068
rect -1830 8973 -1681 9067
rect -1587 8973 -1586 9067
rect -1830 8972 -1586 8973
rect -1452 7356 -1380 7357
rect -1452 7286 -1451 7356
rect -1381 7286 -1380 7356
rect -1452 7285 -1380 7286
rect -1446 7210 -1386 7285
rect -1807 7114 -1386 7210
rect -14358 2550 1314 2551
rect -14358 1870 633 2550
rect 1313 1870 1314 2550
rect -14358 1869 1314 1870
rect -14358 1536 -1847 1869
use bjt  bjt_0
timestamp 1718348362
transform 0 -1 7195 1 0 1540
box -387 -387 7324 7279
use cap_op  cap_op_0
timestamp 1718554435
transform 1 0 -5617 0 1 11002
box -12037 -11160 3906 3480
use differential_pair  differential_pair_0
timestamp 1717432846
transform 1 0 4692 0 1 15013
box -567 -89 4001 858
use digital  digital_0
timestamp 1718522076
transform 0 1 3934 1 0 10121
box -202 -4018 2522 1619
use nmos_startup  nmos_startup_0
timestamp 1717696245
transform 1 0 -1078 0 1 16928
box -204 -148 746 686
use nmos_tail_current  nmos_tail_current_0
timestamp 1717870580
transform 1 0 100 0 1 16054
box -315 -141 8593 1579
use pmos_current_bgr  pmos_current_bgr_0
timestamp 1717985588
transform 1 0 -16475 0 1 17121
box -227 -1493 8585 556
use pmos_current_bgr_2  pmos_current_bgr_2_0
timestamp 1717930986
transform -1 0 -3210 0 1 17072
box -225 -1450 4471 516
use pmos_iptat  pmos_iptat_0
timestamp 1717930986
transform 1 0 -12328 0 1 14730
box -191 -104 4438 898
use pmos_startup  pmos_startup_0
timestamp 1717930986
transform -1 0 -3176 0 1 15183
box -191 -509 4437 439
use res_trim  res_trim_0
timestamp 1718517160
transform 0 -1 8672 1 0 17734
box -31 -51 1533 16353
use resist_const  resist_const_0
timestamp 1717597558
transform 1 0 -19769 0 1 24804
box 2248 -3973 28492 -2077
use resistor_op_tt  resistor_op_tt_0
timestamp 1717870769
transform 0 -1 5318 1 0 15108
box -441 2216 791 5516
use resistorstart  resistorstart_0
timestamp 1717756107
transform 1 0 -13132 0 -1 20778
box -53 -53 21855 1511
<< labels >>
flabel metal2 9110 11276 9110 11276 0 FreeSans 1600 0 0 0 AVDD
port 0 nsew
flabel metal1 9110 10277 9110 10277 0 FreeSans 1600 0 0 0 DVDD
port 1 nsew
flabel metal1 9025 12135 9025 12135 0 FreeSans 1600 0 0 0 VBGTC
port 4 nsew
flabel metal1 8928 9914 8928 9914 0 FreeSans 1600 0 0 0 VENA
port 5 nsew
flabel metal1 8992 9711 8992 9711 0 FreeSans 1600 0 0 0 DVSS
port 6 nsew
flabel metal1 8963 9542 8963 9542 0 FreeSans 1600 0 0 0 TRIM0
port 7 nsew
flabel metal1 8956 9419 8956 9419 0 FreeSans 1600 0 0 0 TRIM1
port 8 nsew
flabel metal1 8975 9310 8975 9310 0 FreeSans 1600 0 0 0 TRIM2
port 9 nsew
flabel metal1 8962 9147 8962 9147 0 FreeSans 1600 0 0 0 TRIM3
port 10 nsew
flabel metal4 -17674 17728 -17674 17728 0 FreeSans 1600 0 0 0 AVSS
port 11 nsew
flabel metal2 9133 10922 9133 10922 0 FreeSans 1600 0 0 0 VBGSC
port 2 nsew
flabel metal1 9134 11659 9134 11659 0 FreeSans 1600 0 0 0 ENA
port 3 nsew
flabel metal1 -17884 15577 -17884 15577 0 FreeSans 1600 0 0 0 IPTAT
port 12 nsew
flabel metal3 -17907 22357 -17907 22357 0 FreeSans 1600 0 0 0 VREF
port 14 nsew
<< end >>
