magic
tech sky130A
magscale 1 2
timestamp 1717222322
<< nwell >>
rect -723 -198 723 164
<< pmos >>
rect -629 -136 -29 64
rect 29 -136 629 64
<< pdiff >>
rect -687 52 -629 64
rect -687 -124 -675 52
rect -641 -124 -629 52
rect -687 -136 -629 -124
rect -29 52 29 64
rect -29 -124 -17 52
rect 17 -124 29 52
rect -29 -136 29 -124
rect 629 52 687 64
rect 629 -124 641 52
rect 675 -124 687 52
rect 629 -136 687 -124
<< pdiffc >>
rect -675 -124 -641 52
rect -17 -124 17 52
rect 641 -124 675 52
<< poly >>
rect -487 145 -171 161
rect -487 128 -471 145
rect -629 111 -471 128
rect -187 128 -171 145
rect 171 145 487 161
rect 171 128 187 145
rect -187 111 -29 128
rect -629 64 -29 111
rect 29 111 187 128
rect 471 128 487 145
rect 471 111 629 128
rect 29 64 629 111
rect -629 -162 -29 -136
rect 29 -162 629 -136
<< polycont >>
rect -471 111 -187 145
rect 187 111 471 145
<< locali >>
rect -487 111 -471 145
rect -187 111 -171 145
rect 171 111 187 145
rect 471 111 487 145
rect -675 52 -641 68
rect -675 -140 -641 -124
rect -17 52 17 68
rect -17 -140 17 -124
rect 641 52 675 68
rect 641 -140 675 -124
<< viali >>
rect -471 111 -187 145
rect 187 111 471 145
rect -675 -124 -641 52
rect -17 -124 17 52
rect 641 -124 675 52
<< metal1 >>
rect -483 145 -175 151
rect -483 111 -471 145
rect -187 111 -175 145
rect -483 105 -175 111
rect 175 145 483 151
rect 175 111 187 145
rect 471 111 483 145
rect 175 105 483 111
rect -681 52 -635 64
rect -681 -124 -675 52
rect -641 -124 -635 52
rect -681 -136 -635 -124
rect -23 52 23 64
rect -23 -124 -17 52
rect 17 -124 23 52
rect -23 -136 23 -124
rect 635 52 681 64
rect 635 -124 641 52
rect 675 -124 681 52
rect 635 -136 681 -124
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 3 m 1 nf 2 diffcov 100 polycov 50 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
