magic
tech sky130A
magscale 1 2
timestamp 1717930986
<< nwell >>
rect -191 -509 4437 439
<< nsubdiff >>
rect -155 369 -95 403
rect 4341 369 4401 403
rect -155 343 -121 369
rect 4367 343 4401 369
rect -155 -439 -121 -413
rect 4367 -439 4401 -413
rect -155 -473 -95 -439
rect 4341 -473 4401 -439
<< nsubdiffcont >>
rect -95 369 4341 403
rect -155 -413 -121 343
rect 4367 -413 4401 343
rect -95 -473 4341 -439
<< poly >>
rect 6 -2 36 93
rect -56 -18 36 -2
rect -56 -52 -40 -18
rect -6 -52 36 -18
rect -56 -68 36 -52
rect 6 -152 36 -68
rect 4210 -2 4240 91
rect 4210 -18 4302 -2
rect 4210 -52 4252 -18
rect 4286 -52 4302 -18
rect 4210 -68 4302 -52
rect 4210 -147 4240 -68
<< polycont >>
rect -40 -52 -6 -18
rect 4252 -52 4286 -18
<< locali >>
rect -155 369 -95 403
rect 4341 369 4401 403
rect -155 343 -121 369
rect 4367 343 4401 369
rect -40 -18 -6 -2
rect -40 -68 -6 -52
rect 4252 -18 4286 -2
rect 4252 -68 4286 -52
rect -155 -439 -121 -413
rect 4367 -439 4401 -413
rect -155 -473 -95 -439
rect 4341 -473 4401 -439
<< viali >>
rect 2106 369 2140 403
rect -155 -52 -121 -18
rect -40 -52 -6 -18
rect 4252 -52 4286 -18
rect 4367 -52 4401 -18
rect 2106 -473 2140 -439
<< metal1 >>
rect 2094 403 2152 409
rect 2094 369 2106 403
rect 2140 369 2152 403
rect 2094 288 2152 369
rect 2087 112 2097 288
rect 2149 112 2159 288
rect -46 -12 0 101
rect 42 59 88 101
rect 42 13 620 59
rect 1594 13 2669 59
rect 4158 -12 4204 101
rect -167 -18 0 -12
rect -167 -52 -155 -18
rect -121 -52 -40 -18
rect -6 -52 0 -18
rect -167 -58 0 -52
rect -46 -83 0 -58
rect 3872 -58 4204 -12
rect 4246 -12 4292 107
rect 4246 -18 4413 -12
rect 4246 -52 4252 -18
rect 4286 -52 4367 -18
rect 4401 -52 4413 -18
rect 4246 -58 4413 -52
rect 3872 -83 3918 -58
rect -46 -129 598 -83
rect 2648 -129 3918 -83
rect -46 -171 0 -129
rect 42 -179 88 -129
rect 4246 -175 4292 -58
rect 2087 -358 2097 -182
rect 2149 -358 2159 -182
rect 2094 -439 2152 -358
rect 4158 -406 4204 -360
rect 2094 -473 2106 -439
rect 2140 -473 2152 -439
rect 2094 -479 2152 -473
<< via1 >>
rect 2097 112 2149 288
rect 2097 -358 2149 -182
<< metal2 >>
rect 2097 288 2149 298
rect 2097 -182 2149 112
rect 2097 -368 2149 -358
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_1
timestamp 1717765832
transform 1 0 4225 0 1 -270
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_2
timestamp 1717765832
transform 1 0 21 0 1 200
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_3
timestamp 1717765832
transform 1 0 4225 0 1 200
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_4
timestamp 1717765832
transform 1 0 21 0 1 -270
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_8RMJP2  sky130_fd_pr__pfet_01v8_8RMJP2_0
timestamp 1717765832
transform 1 0 2123 0 1 -234
box -2123 -198 2123 164
use sky130_fd_pr__pfet_01v8_CVRJBD  sky130_fd_pr__pfet_01v8_CVRJBD_1
timestamp 1717765832
transform 1 0 2123 0 1 164
box -2123 -164 2123 198
<< labels >>
flabel metal1 62 24 62 24 0 FreeSans 1600 0 0 0 D3
port 1 nsew
flabel metal1 4184 50 4184 50 0 FreeSans 1600 0 0 0 D2
port 2 nsew
flabel metal1 4180 -390 4180 -390 0 FreeSans 1600 0 0 0 D4
port 3 nsew
flabel metal1 2116 -418 2116 -418 0 FreeSans 1600 0 0 0 VDDE
port 4 nsew
<< end >>
