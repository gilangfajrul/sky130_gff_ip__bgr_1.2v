magic
tech sky130A
magscale 1 2
timestamp 1717755416
<< pwell >>
rect -616 -15290 616 15290
<< psubdiff >>
rect -580 15220 -484 15254
rect 484 15220 580 15254
rect -580 15158 -546 15220
rect 546 15158 580 15220
rect -580 -15220 -546 -15158
rect 546 -15220 580 -15158
rect -580 -15254 -484 -15220
rect 484 -15254 580 -15220
<< psubdiffcont >>
rect -484 15220 484 15254
rect -580 -15158 -546 15158
rect 546 -15158 580 15158
rect -484 -15254 484 -15220
<< xpolycontact >>
rect -450 14692 -380 15124
rect -450 10892 -380 11324
rect -284 14692 -214 15124
rect -284 10892 -214 11324
rect -118 14692 -48 15124
rect -118 10892 -48 11324
rect 48 14692 118 15124
rect 48 10892 118 11324
rect 214 14692 284 15124
rect 214 10892 284 11324
rect 380 14692 450 15124
rect 380 10892 450 11324
rect -450 10356 -380 10788
rect -450 6556 -380 6988
rect -284 10356 -214 10788
rect -284 6556 -214 6988
rect -118 10356 -48 10788
rect -118 6556 -48 6988
rect 48 10356 118 10788
rect 48 6556 118 6988
rect 214 10356 284 10788
rect 214 6556 284 6988
rect 380 10356 450 10788
rect 380 6556 450 6988
rect -450 6020 -380 6452
rect -450 2220 -380 2652
rect -284 6020 -214 6452
rect -284 2220 -214 2652
rect -118 6020 -48 6452
rect -118 2220 -48 2652
rect 48 6020 118 6452
rect 48 2220 118 2652
rect 214 6020 284 6452
rect 214 2220 284 2652
rect 380 6020 450 6452
rect 380 2220 450 2652
rect -450 1684 -380 2116
rect -450 -2116 -380 -1684
rect -284 1684 -214 2116
rect -284 -2116 -214 -1684
rect -118 1684 -48 2116
rect -118 -2116 -48 -1684
rect 48 1684 118 2116
rect 48 -2116 118 -1684
rect 214 1684 284 2116
rect 214 -2116 284 -1684
rect 380 1684 450 2116
rect 380 -2116 450 -1684
rect -450 -2652 -380 -2220
rect -450 -6452 -380 -6020
rect -284 -2652 -214 -2220
rect -284 -6452 -214 -6020
rect -118 -2652 -48 -2220
rect -118 -6452 -48 -6020
rect 48 -2652 118 -2220
rect 48 -6452 118 -6020
rect 214 -2652 284 -2220
rect 214 -6452 284 -6020
rect 380 -2652 450 -2220
rect 380 -6452 450 -6020
rect -450 -6988 -380 -6556
rect -450 -10788 -380 -10356
rect -284 -6988 -214 -6556
rect -284 -10788 -214 -10356
rect -118 -6988 -48 -6556
rect -118 -10788 -48 -10356
rect 48 -6988 118 -6556
rect 48 -10788 118 -10356
rect 214 -6988 284 -6556
rect 214 -10788 284 -10356
rect 380 -6988 450 -6556
rect 380 -10788 450 -10356
rect -450 -11324 -380 -10892
rect -450 -15124 -380 -14692
rect -284 -11324 -214 -10892
rect -284 -15124 -214 -14692
rect -118 -11324 -48 -10892
rect -118 -15124 -48 -14692
rect 48 -11324 118 -10892
rect 48 -15124 118 -14692
rect 214 -11324 284 -10892
rect 214 -15124 284 -14692
rect 380 -11324 450 -10892
rect 380 -15124 450 -14692
<< ppolyres >>
rect -450 11324 -380 14692
rect -284 11324 -214 14692
rect -118 11324 -48 14692
rect 48 11324 118 14692
rect 214 11324 284 14692
rect 380 11324 450 14692
rect -450 6988 -380 10356
rect -284 6988 -214 10356
rect -118 6988 -48 10356
rect 48 6988 118 10356
rect 214 6988 284 10356
rect 380 6988 450 10356
rect -450 2652 -380 6020
rect -284 2652 -214 6020
rect -118 2652 -48 6020
rect 48 2652 118 6020
rect 214 2652 284 6020
rect 380 2652 450 6020
rect -450 -1684 -380 1684
rect -284 -1684 -214 1684
rect -118 -1684 -48 1684
rect 48 -1684 118 1684
rect 214 -1684 284 1684
rect 380 -1684 450 1684
rect -450 -6020 -380 -2652
rect -284 -6020 -214 -2652
rect -118 -6020 -48 -2652
rect 48 -6020 118 -2652
rect 214 -6020 284 -2652
rect 380 -6020 450 -2652
rect -450 -10356 -380 -6988
rect -284 -10356 -214 -6988
rect -118 -10356 -48 -6988
rect 48 -10356 118 -6988
rect 214 -10356 284 -6988
rect 380 -10356 450 -6988
rect -450 -14692 -380 -11324
rect -284 -14692 -214 -11324
rect -118 -14692 -48 -11324
rect 48 -14692 118 -11324
rect 214 -14692 284 -11324
rect 380 -14692 450 -11324
<< locali >>
rect -580 15220 -484 15254
rect 484 15220 580 15254
rect -580 15158 -546 15220
rect 546 15158 580 15220
rect -580 -15220 -546 -15158
rect 546 -15220 580 -15158
rect -580 -15254 -484 -15220
rect 484 -15254 580 -15220
<< viali >>
rect -434 14709 -396 15106
rect -268 14709 -230 15106
rect -102 14709 -64 15106
rect 64 14709 102 15106
rect 230 14709 268 15106
rect 396 14709 434 15106
rect -434 10910 -396 11307
rect -268 10910 -230 11307
rect -102 10910 -64 11307
rect 64 10910 102 11307
rect 230 10910 268 11307
rect 396 10910 434 11307
rect -434 10373 -396 10770
rect -268 10373 -230 10770
rect -102 10373 -64 10770
rect 64 10373 102 10770
rect 230 10373 268 10770
rect 396 10373 434 10770
rect -434 6574 -396 6971
rect -268 6574 -230 6971
rect -102 6574 -64 6971
rect 64 6574 102 6971
rect 230 6574 268 6971
rect 396 6574 434 6971
rect -434 6037 -396 6434
rect -268 6037 -230 6434
rect -102 6037 -64 6434
rect 64 6037 102 6434
rect 230 6037 268 6434
rect 396 6037 434 6434
rect -434 2238 -396 2635
rect -268 2238 -230 2635
rect -102 2238 -64 2635
rect 64 2238 102 2635
rect 230 2238 268 2635
rect 396 2238 434 2635
rect -434 1701 -396 2098
rect -268 1701 -230 2098
rect -102 1701 -64 2098
rect 64 1701 102 2098
rect 230 1701 268 2098
rect 396 1701 434 2098
rect -434 -2098 -396 -1701
rect -268 -2098 -230 -1701
rect -102 -2098 -64 -1701
rect 64 -2098 102 -1701
rect 230 -2098 268 -1701
rect 396 -2098 434 -1701
rect -434 -2635 -396 -2238
rect -268 -2635 -230 -2238
rect -102 -2635 -64 -2238
rect 64 -2635 102 -2238
rect 230 -2635 268 -2238
rect 396 -2635 434 -2238
rect -434 -6434 -396 -6037
rect -268 -6434 -230 -6037
rect -102 -6434 -64 -6037
rect 64 -6434 102 -6037
rect 230 -6434 268 -6037
rect 396 -6434 434 -6037
rect -434 -6971 -396 -6574
rect -268 -6971 -230 -6574
rect -102 -6971 -64 -6574
rect 64 -6971 102 -6574
rect 230 -6971 268 -6574
rect 396 -6971 434 -6574
rect -434 -10770 -396 -10373
rect -268 -10770 -230 -10373
rect -102 -10770 -64 -10373
rect 64 -10770 102 -10373
rect 230 -10770 268 -10373
rect 396 -10770 434 -10373
rect -434 -11307 -396 -10910
rect -268 -11307 -230 -10910
rect -102 -11307 -64 -10910
rect 64 -11307 102 -10910
rect 230 -11307 268 -10910
rect 396 -11307 434 -10910
rect -434 -15106 -396 -14709
rect -268 -15106 -230 -14709
rect -102 -15106 -64 -14709
rect 64 -15106 102 -14709
rect 230 -15106 268 -14709
rect 396 -15106 434 -14709
<< metal1 >>
rect -440 15106 -390 15118
rect -440 14709 -434 15106
rect -396 14709 -390 15106
rect -440 14697 -390 14709
rect -274 15106 -224 15118
rect -274 14709 -268 15106
rect -230 14709 -224 15106
rect -274 14697 -224 14709
rect -108 15106 -58 15118
rect -108 14709 -102 15106
rect -64 14709 -58 15106
rect -108 14697 -58 14709
rect 58 15106 108 15118
rect 58 14709 64 15106
rect 102 14709 108 15106
rect 58 14697 108 14709
rect 224 15106 274 15118
rect 224 14709 230 15106
rect 268 14709 274 15106
rect 224 14697 274 14709
rect 390 15106 440 15118
rect 390 14709 396 15106
rect 434 14709 440 15106
rect 390 14697 440 14709
rect -440 11307 -390 11319
rect -440 10910 -434 11307
rect -396 10910 -390 11307
rect -440 10898 -390 10910
rect -274 11307 -224 11319
rect -274 10910 -268 11307
rect -230 10910 -224 11307
rect -274 10898 -224 10910
rect -108 11307 -58 11319
rect -108 10910 -102 11307
rect -64 10910 -58 11307
rect -108 10898 -58 10910
rect 58 11307 108 11319
rect 58 10910 64 11307
rect 102 10910 108 11307
rect 58 10898 108 10910
rect 224 11307 274 11319
rect 224 10910 230 11307
rect 268 10910 274 11307
rect 224 10898 274 10910
rect 390 11307 440 11319
rect 390 10910 396 11307
rect 434 10910 440 11307
rect 390 10898 440 10910
rect -440 10770 -390 10782
rect -440 10373 -434 10770
rect -396 10373 -390 10770
rect -440 10361 -390 10373
rect -274 10770 -224 10782
rect -274 10373 -268 10770
rect -230 10373 -224 10770
rect -274 10361 -224 10373
rect -108 10770 -58 10782
rect -108 10373 -102 10770
rect -64 10373 -58 10770
rect -108 10361 -58 10373
rect 58 10770 108 10782
rect 58 10373 64 10770
rect 102 10373 108 10770
rect 58 10361 108 10373
rect 224 10770 274 10782
rect 224 10373 230 10770
rect 268 10373 274 10770
rect 224 10361 274 10373
rect 390 10770 440 10782
rect 390 10373 396 10770
rect 434 10373 440 10770
rect 390 10361 440 10373
rect -440 6971 -390 6983
rect -440 6574 -434 6971
rect -396 6574 -390 6971
rect -440 6562 -390 6574
rect -274 6971 -224 6983
rect -274 6574 -268 6971
rect -230 6574 -224 6971
rect -274 6562 -224 6574
rect -108 6971 -58 6983
rect -108 6574 -102 6971
rect -64 6574 -58 6971
rect -108 6562 -58 6574
rect 58 6971 108 6983
rect 58 6574 64 6971
rect 102 6574 108 6971
rect 58 6562 108 6574
rect 224 6971 274 6983
rect 224 6574 230 6971
rect 268 6574 274 6971
rect 224 6562 274 6574
rect 390 6971 440 6983
rect 390 6574 396 6971
rect 434 6574 440 6971
rect 390 6562 440 6574
rect -440 6434 -390 6446
rect -440 6037 -434 6434
rect -396 6037 -390 6434
rect -440 6025 -390 6037
rect -274 6434 -224 6446
rect -274 6037 -268 6434
rect -230 6037 -224 6434
rect -274 6025 -224 6037
rect -108 6434 -58 6446
rect -108 6037 -102 6434
rect -64 6037 -58 6434
rect -108 6025 -58 6037
rect 58 6434 108 6446
rect 58 6037 64 6434
rect 102 6037 108 6434
rect 58 6025 108 6037
rect 224 6434 274 6446
rect 224 6037 230 6434
rect 268 6037 274 6434
rect 224 6025 274 6037
rect 390 6434 440 6446
rect 390 6037 396 6434
rect 434 6037 440 6434
rect 390 6025 440 6037
rect -440 2635 -390 2647
rect -440 2238 -434 2635
rect -396 2238 -390 2635
rect -440 2226 -390 2238
rect -274 2635 -224 2647
rect -274 2238 -268 2635
rect -230 2238 -224 2635
rect -274 2226 -224 2238
rect -108 2635 -58 2647
rect -108 2238 -102 2635
rect -64 2238 -58 2635
rect -108 2226 -58 2238
rect 58 2635 108 2647
rect 58 2238 64 2635
rect 102 2238 108 2635
rect 58 2226 108 2238
rect 224 2635 274 2647
rect 224 2238 230 2635
rect 268 2238 274 2635
rect 224 2226 274 2238
rect 390 2635 440 2647
rect 390 2238 396 2635
rect 434 2238 440 2635
rect 390 2226 440 2238
rect -440 2098 -390 2110
rect -440 1701 -434 2098
rect -396 1701 -390 2098
rect -440 1689 -390 1701
rect -274 2098 -224 2110
rect -274 1701 -268 2098
rect -230 1701 -224 2098
rect -274 1689 -224 1701
rect -108 2098 -58 2110
rect -108 1701 -102 2098
rect -64 1701 -58 2098
rect -108 1689 -58 1701
rect 58 2098 108 2110
rect 58 1701 64 2098
rect 102 1701 108 2098
rect 58 1689 108 1701
rect 224 2098 274 2110
rect 224 1701 230 2098
rect 268 1701 274 2098
rect 224 1689 274 1701
rect 390 2098 440 2110
rect 390 1701 396 2098
rect 434 1701 440 2098
rect 390 1689 440 1701
rect -440 -1701 -390 -1689
rect -440 -2098 -434 -1701
rect -396 -2098 -390 -1701
rect -440 -2110 -390 -2098
rect -274 -1701 -224 -1689
rect -274 -2098 -268 -1701
rect -230 -2098 -224 -1701
rect -274 -2110 -224 -2098
rect -108 -1701 -58 -1689
rect -108 -2098 -102 -1701
rect -64 -2098 -58 -1701
rect -108 -2110 -58 -2098
rect 58 -1701 108 -1689
rect 58 -2098 64 -1701
rect 102 -2098 108 -1701
rect 58 -2110 108 -2098
rect 224 -1701 274 -1689
rect 224 -2098 230 -1701
rect 268 -2098 274 -1701
rect 224 -2110 274 -2098
rect 390 -1701 440 -1689
rect 390 -2098 396 -1701
rect 434 -2098 440 -1701
rect 390 -2110 440 -2098
rect -440 -2238 -390 -2226
rect -440 -2635 -434 -2238
rect -396 -2635 -390 -2238
rect -440 -2647 -390 -2635
rect -274 -2238 -224 -2226
rect -274 -2635 -268 -2238
rect -230 -2635 -224 -2238
rect -274 -2647 -224 -2635
rect -108 -2238 -58 -2226
rect -108 -2635 -102 -2238
rect -64 -2635 -58 -2238
rect -108 -2647 -58 -2635
rect 58 -2238 108 -2226
rect 58 -2635 64 -2238
rect 102 -2635 108 -2238
rect 58 -2647 108 -2635
rect 224 -2238 274 -2226
rect 224 -2635 230 -2238
rect 268 -2635 274 -2238
rect 224 -2647 274 -2635
rect 390 -2238 440 -2226
rect 390 -2635 396 -2238
rect 434 -2635 440 -2238
rect 390 -2647 440 -2635
rect -440 -6037 -390 -6025
rect -440 -6434 -434 -6037
rect -396 -6434 -390 -6037
rect -440 -6446 -390 -6434
rect -274 -6037 -224 -6025
rect -274 -6434 -268 -6037
rect -230 -6434 -224 -6037
rect -274 -6446 -224 -6434
rect -108 -6037 -58 -6025
rect -108 -6434 -102 -6037
rect -64 -6434 -58 -6037
rect -108 -6446 -58 -6434
rect 58 -6037 108 -6025
rect 58 -6434 64 -6037
rect 102 -6434 108 -6037
rect 58 -6446 108 -6434
rect 224 -6037 274 -6025
rect 224 -6434 230 -6037
rect 268 -6434 274 -6037
rect 224 -6446 274 -6434
rect 390 -6037 440 -6025
rect 390 -6434 396 -6037
rect 434 -6434 440 -6037
rect 390 -6446 440 -6434
rect -440 -6574 -390 -6562
rect -440 -6971 -434 -6574
rect -396 -6971 -390 -6574
rect -440 -6983 -390 -6971
rect -274 -6574 -224 -6562
rect -274 -6971 -268 -6574
rect -230 -6971 -224 -6574
rect -274 -6983 -224 -6971
rect -108 -6574 -58 -6562
rect -108 -6971 -102 -6574
rect -64 -6971 -58 -6574
rect -108 -6983 -58 -6971
rect 58 -6574 108 -6562
rect 58 -6971 64 -6574
rect 102 -6971 108 -6574
rect 58 -6983 108 -6971
rect 224 -6574 274 -6562
rect 224 -6971 230 -6574
rect 268 -6971 274 -6574
rect 224 -6983 274 -6971
rect 390 -6574 440 -6562
rect 390 -6971 396 -6574
rect 434 -6971 440 -6574
rect 390 -6983 440 -6971
rect -440 -10373 -390 -10361
rect -440 -10770 -434 -10373
rect -396 -10770 -390 -10373
rect -440 -10782 -390 -10770
rect -274 -10373 -224 -10361
rect -274 -10770 -268 -10373
rect -230 -10770 -224 -10373
rect -274 -10782 -224 -10770
rect -108 -10373 -58 -10361
rect -108 -10770 -102 -10373
rect -64 -10770 -58 -10373
rect -108 -10782 -58 -10770
rect 58 -10373 108 -10361
rect 58 -10770 64 -10373
rect 102 -10770 108 -10373
rect 58 -10782 108 -10770
rect 224 -10373 274 -10361
rect 224 -10770 230 -10373
rect 268 -10770 274 -10373
rect 224 -10782 274 -10770
rect 390 -10373 440 -10361
rect 390 -10770 396 -10373
rect 434 -10770 440 -10373
rect 390 -10782 440 -10770
rect -440 -10910 -390 -10898
rect -440 -11307 -434 -10910
rect -396 -11307 -390 -10910
rect -440 -11319 -390 -11307
rect -274 -10910 -224 -10898
rect -274 -11307 -268 -10910
rect -230 -11307 -224 -10910
rect -274 -11319 -224 -11307
rect -108 -10910 -58 -10898
rect -108 -11307 -102 -10910
rect -64 -11307 -58 -10910
rect -108 -11319 -58 -11307
rect 58 -10910 108 -10898
rect 58 -11307 64 -10910
rect 102 -11307 108 -10910
rect 58 -11319 108 -11307
rect 224 -10910 274 -10898
rect 224 -11307 230 -10910
rect 268 -11307 274 -10910
rect 224 -11319 274 -11307
rect 390 -10910 440 -10898
rect 390 -11307 396 -10910
rect 434 -11307 440 -10910
rect 390 -11319 440 -11307
rect -440 -14709 -390 -14697
rect -440 -15106 -434 -14709
rect -396 -15106 -390 -14709
rect -440 -15118 -390 -15106
rect -274 -14709 -224 -14697
rect -274 -15106 -268 -14709
rect -230 -15106 -224 -14709
rect -274 -15118 -224 -15106
rect -108 -14709 -58 -14697
rect -108 -15106 -102 -14709
rect -64 -15106 -58 -14709
rect -108 -15118 -58 -15106
rect 58 -14709 108 -14697
rect 58 -15106 64 -14709
rect 102 -15106 108 -14709
rect 58 -15118 108 -15106
rect 224 -14709 274 -14697
rect 224 -15106 230 -14709
rect 268 -15106 274 -14709
rect 224 -15118 274 -15106
rect 390 -14709 440 -14697
rect 390 -15106 396 -14709
rect 434 -15106 440 -14709
rect 390 -15118 440 -15106
<< properties >>
string FIXED_BBOX -563 -15237 563 15237
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.350 l 17 m 7 nx 6 wmin 0.350 lmin 0.50 rho 319.8 val 16.646k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
