* NGSPICE file created from bgr_op5_block_rev2.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_CJRLGR a_n287_n255# a_n229_n343# a_229_n255# a_229_55#
+ a_n29_n255# a_n287_55# a_n29_55# a_29_n343# VSUBS
X0 a_229_55# a_29_n343# a_n29_55# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1 a_n29_n255# a_n229_n343# a_n287_n255# VSUBS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2 a_229_n255# a_29_n343# a_n29_n255# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3 a_n29_55# a_n229_n343# a_n287_55# VSUBS sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
C0 a_n229_n343# a_29_n343# 0.14779f
C1 a_229_n255# VSUBS 0.114051f
C2 a_n287_n255# VSUBS 0.114051f
C3 a_229_55# VSUBS 0.114051f
C4 a_n287_55# VSUBS 0.114051f
C5 a_29_n343# VSUBS 0.824774f
C6 a_n229_n343# VSUBS 0.824774f
.ends

.subckt sky130_fd_pr__nfet_01v8_6H9P4D a_n73_n100# a_15_n100# a_n15_n126# VSUBS
X0 a_15_n100# a_n15_n126# a_n73_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
C0 a_n73_n100# a_15_n100# 0.162113f
C1 a_15_n100# VSUBS 0.118371f
C2 a_n73_n100# VSUBS 0.118371f
.ends

.subckt nmos_startup AVSS D1 G1
Xsky130_fd_pr__nfet_01v8_CJRLGR_0 D1 G1 D1 D1 AVSS D1 AVSS G1 AVSS sky130_fd_pr__nfet_01v8_CJRLGR
Xsky130_fd_pr__nfet_01v8_6H9P4D_0 D1 D1 D1 AVSS sky130_fd_pr__nfet_01v8_6H9P4D
Xsky130_fd_pr__nfet_01v8_6H9P4D_1 D1 D1 D1 AVSS sky130_fd_pr__nfet_01v8_6H9P4D
Xsky130_fd_pr__nfet_01v8_6H9P4D_3 D1 D1 D1 AVSS sky130_fd_pr__nfet_01v8_6H9P4D
Xsky130_fd_pr__nfet_01v8_6H9P4D_4 D1 D1 D1 AVSS sky130_fd_pr__nfet_01v8_6H9P4D
C0 AVSS G1 0.758576f
C1 D1 G1 0.466067f
C2 AVSS D1 0.381248f
C3 AVSS 0 -0.306076f
C4 D1 0 1.748479f
C5 G1 0 1.308701f
.ends

.subckt sky130_fd_pr__res_high_po_0p35_9NXREG a_380_2220# a_48_1684# a_380_6556# a_546_n2652#
+ a_546_n6988# a_n118_10356# a_214_6020# a_n284_n6452# a_n616_2220# a_n616_6556# a_n616_n6452#
+ a_214_n10788# a_214_2220# a_n284_n2652# a_380_n2116# a_n284_n6988# a_214_6556# a_546_1684#
+ a_n616_n2652# a_n616_n10788# a_48_6020# a_n616_n6988# a_380_10356# a_n118_n6452#
+ a_546_n10788# a_48_2220# a_48_6556# a_n450_n2116# a_n450_1684# a_n118_n2652# a_214_n2116#
+ a_n118_n6988# a_546_6020# a_n450_n10788# a_n450_10356# a_214_10356# a_n284_1684#
+ a_380_n6452# a_380_n10788# a_546_2220# a_546_6556# a_n118_n10788# a_380_n2652# a_n450_6020#
+ a_48_n2116# a_380_n6988# a_n118_1684# a_n450_n6452# a_48_10356# a_n450_2220# a_214_n6452#
+ a_n284_6020# a_n450_6556# a_546_n2116# a_n450_n2652# a_n450_n6988# a_n284_2220#
+ a_380_1684# a_214_n2652# a_546_10356# a_214_n6988# a_n284_6556# a_n118_6020# a_n616_1684#
+ a_n284_n2116# a_48_n6452# a_n284_n10788# a_n616_n2116# a_n284_10356# a_n746_n10918#
+ a_n118_2220# a_214_1684# a_n118_6556# a_n616_10356# a_48_n2652# a_48_n6988# a_380_6020#
+ a_546_n6452# a_n616_6020# a_n118_n2116# a_48_n10788#
X0 a_n284_10356# a_n284_6556# a_n746_n10918# sky130_fd_pr__res_high_po_0p35 l=17
X1 a_380_n6988# a_380_n10788# a_n746_n10918# sky130_fd_pr__res_high_po_0p35 l=17
X2 a_n450_6020# a_n450_2220# a_n746_n10918# sky130_fd_pr__res_high_po_0p35 l=17
X3 a_48_6020# a_48_2220# a_n746_n10918# sky130_fd_pr__res_high_po_0p35 l=17
X4 a_48_10356# a_48_6556# a_n746_n10918# sky130_fd_pr__res_high_po_0p35 l=17
X5 a_n118_n6988# a_n118_n10788# a_n746_n10918# sky130_fd_pr__res_high_po_0p35 l=17
X6 a_n450_10356# a_n450_6556# a_n746_n10918# sky130_fd_pr__res_high_po_0p35 l=17
X7 a_214_n2652# a_214_n6452# a_n746_n10918# sky130_fd_pr__res_high_po_0p35 l=17
X8 a_n118_6020# a_n118_2220# a_n746_n10918# sky130_fd_pr__res_high_po_0p35 l=17
X9 a_n118_10356# a_n118_6556# a_n746_n10918# sky130_fd_pr__res_high_po_0p35 l=17
X10 a_214_1684# a_214_n2116# a_n746_n10918# sky130_fd_pr__res_high_po_0p35 l=17
X11 a_n450_n6988# a_n450_n10788# a_n746_n10918# sky130_fd_pr__res_high_po_0p35 l=17
X12 a_n118_n2652# a_n118_n6452# a_n746_n10918# sky130_fd_pr__res_high_po_0p35 l=17
X13 a_n284_n6988# a_n284_n10788# a_n746_n10918# sky130_fd_pr__res_high_po_0p35 l=17
X14 a_n118_1684# a_n118_n2116# a_n746_n10918# sky130_fd_pr__res_high_po_0p35 l=17
X15 a_n616_n2652# a_n616_n6452# a_n746_n10918# sky130_fd_pr__res_high_po_0p35 l=17
X16 a_n616_n6988# a_n616_n10788# a_n746_n10918# sky130_fd_pr__res_high_po_0p35 l=17
X17 a_n616_6020# a_n616_2220# a_n746_n10918# sky130_fd_pr__res_high_po_0p35 l=17
X18 a_380_6020# a_380_2220# a_n746_n10918# sky130_fd_pr__res_high_po_0p35 l=17
X19 a_48_n6988# a_48_n10788# a_n746_n10918# sky130_fd_pr__res_high_po_0p35 l=17
X20 a_n616_10356# a_n616_6556# a_n746_n10918# sky130_fd_pr__res_high_po_0p35 l=17
X21 a_380_10356# a_380_6556# a_n746_n10918# sky130_fd_pr__res_high_po_0p35 l=17
X22 a_380_n2652# a_380_n6452# a_n746_n10918# sky130_fd_pr__res_high_po_0p35 l=17
X23 a_546_n2652# a_546_n6452# a_n746_n10918# sky130_fd_pr__res_high_po_0p35 l=17
X24 a_n616_1684# a_n616_n2116# a_n746_n10918# sky130_fd_pr__res_high_po_0p35 l=17
X25 a_214_n6988# a_214_n10788# a_n746_n10918# sky130_fd_pr__res_high_po_0p35 l=17
X26 a_546_6020# a_546_2220# a_n746_n10918# sky130_fd_pr__res_high_po_0p35 l=17
X27 a_380_1684# a_380_n2116# a_n746_n10918# sky130_fd_pr__res_high_po_0p35 l=17
X28 a_546_1684# a_546_n2116# a_n746_n10918# sky130_fd_pr__res_high_po_0p35 l=17
X29 a_546_10356# a_546_6556# a_n746_n10918# sky130_fd_pr__res_high_po_0p35 l=17
X30 a_n450_n2652# a_n450_n6452# a_n746_n10918# sky130_fd_pr__res_high_po_0p35 l=17
X31 a_n284_n2652# a_n284_n6452# a_n746_n10918# sky130_fd_pr__res_high_po_0p35 l=17
X32 a_48_n2652# a_48_n6452# a_n746_n10918# sky130_fd_pr__res_high_po_0p35 l=17
X33 a_214_6020# a_214_2220# a_n746_n10918# sky130_fd_pr__res_high_po_0p35 l=17
X34 a_546_n6988# a_546_n10788# a_n746_n10918# sky130_fd_pr__res_high_po_0p35 l=17
X35 a_214_10356# a_214_6556# a_n746_n10918# sky130_fd_pr__res_high_po_0p35 l=17
X36 a_n284_6020# a_n284_2220# a_n746_n10918# sky130_fd_pr__res_high_po_0p35 l=17
X37 a_n450_1684# a_n450_n2116# a_n746_n10918# sky130_fd_pr__res_high_po_0p35 l=17
X38 a_n284_1684# a_n284_n2116# a_n746_n10918# sky130_fd_pr__res_high_po_0p35 l=17
X39 a_48_1684# a_48_n2116# a_n746_n10918# sky130_fd_pr__res_high_po_0p35 l=17
C0 a_n284_1684# a_n118_1684# 0.296258f
C1 a_214_6556# a_48_6556# 0.296258f
C2 a_214_n2116# a_380_n2116# 0.296258f
C3 a_546_2220# a_380_2220# 0.296258f
C4 a_n118_n2652# a_48_n2652# 0.296258f
C5 a_380_n10788# a_546_n10788# 0.296258f
C6 a_n284_6556# a_n118_6556# 0.296258f
C7 a_48_2220# a_214_2220# 0.296258f
C8 a_n118_n6988# a_n284_n6988# 0.296258f
C9 a_214_10356# a_48_10356# 0.296258f
C10 a_n284_1684# a_n450_1684# 0.296258f
C11 a_214_6020# a_48_6020# 0.296258f
C12 a_n450_10356# a_n616_10356# 0.296258f
C13 a_214_n6988# a_48_n6988# 0.296258f
C14 a_n284_6020# a_n450_6020# 0.296258f
C15 a_n284_6556# a_n450_6556# 0.296258f
C16 a_48_2220# a_n118_2220# 0.296258f
C17 a_214_1684# a_380_1684# 0.296258f
C18 a_214_10356# a_380_10356# 0.296258f
C19 a_n450_n2116# a_n616_n2116# 0.296258f
C20 a_n284_10356# a_n118_10356# 0.296258f
C21 a_n118_n6452# a_48_n6452# 0.296258f
C22 a_48_n6988# a_n118_n6988# 0.296258f
C23 a_48_1684# a_214_1684# 0.296258f
C24 a_214_n6452# a_48_n6452# 0.296258f
C25 a_380_n2652# a_214_n2652# 0.296258f
C26 a_n450_n10788# a_n284_n10788# 0.296258f
C27 a_n616_n6452# a_n450_n6452# 0.296258f
C28 a_n284_n2116# a_n118_n2116# 0.296258f
C29 a_n450_6020# a_n616_6020# 0.296258f
C30 a_n118_2220# a_n284_2220# 0.296258f
C31 a_n118_n10788# a_n284_n10788# 0.296258f
C32 a_n450_n2652# a_n284_n2652# 0.296258f
C33 a_n450_n10788# a_n616_n10788# 0.296258f
C34 a_48_1684# a_n118_1684# 0.296258f
C35 a_380_n10788# a_214_n10788# 0.296258f
C36 a_380_n2116# a_546_n2116# 0.296258f
C37 a_n284_n2116# a_n450_n2116# 0.296258f
C38 a_48_n2116# a_n118_n2116# 0.296258f
C39 a_380_n6452# a_214_n6452# 0.296258f
C40 a_380_1684# a_546_1684# 0.296258f
C41 a_380_6556# a_546_6556# 0.296258f
C42 a_380_6020# a_546_6020# 0.296258f
C43 a_48_10356# a_n118_10356# 0.296258f
C44 a_48_n2652# a_214_n2652# 0.296258f
C45 a_n616_6556# a_n450_6556# 0.296258f
C46 a_n118_n2652# a_n284_n2652# 0.296258f
C47 a_380_n6452# a_546_n6452# 0.296258f
C48 a_48_6556# a_n118_6556# 0.296258f
C49 a_546_10356# a_380_10356# 0.296258f
C50 a_n450_2220# a_n284_2220# 0.296258f
C51 a_48_n10788# a_n118_n10788# 0.296258f
C52 a_n284_6020# a_n118_6020# 0.296258f
C53 a_n616_n6988# a_n450_n6988# 0.296258f
C54 a_48_n10788# a_214_n10788# 0.296258f
C55 a_380_2220# a_214_2220# 0.296258f
C56 a_546_n2652# a_380_n2652# 0.296258f
C57 a_380_6556# a_214_6556# 0.296258f
C58 a_380_6020# a_214_6020# 0.296258f
C59 a_n284_n6452# a_n450_n6452# 0.296258f
C60 a_n284_n6452# a_n118_n6452# 0.296258f
C61 a_n616_1684# a_n450_1684# 0.296258f
C62 a_48_6020# a_n118_6020# 0.296258f
C63 a_n450_n2652# a_n616_n2652# 0.296258f
C64 a_214_n6988# a_380_n6988# 0.296258f
C65 a_n450_10356# a_n284_10356# 0.296258f
C66 a_546_n6988# a_380_n6988# 0.296258f
C67 a_n284_n6988# a_n450_n6988# 0.296258f
C68 a_214_n2116# a_48_n2116# 0.296258f
C69 a_n450_2220# a_n616_2220# 0.296258f
C70 a_546_n10788# a_n746_n10918# 0.387223f
C71 a_546_n6988# a_n746_n10918# 0.356961f
C72 a_380_n10788# a_n746_n10918# 0.17691f
C73 a_380_n6988# a_n746_n10918# 0.146647f
C74 a_214_n10788# a_n746_n10918# 0.17691f
C75 a_214_n6988# a_n746_n10918# 0.146647f
C76 a_48_n10788# a_n746_n10918# 0.17691f
C77 a_48_n6988# a_n746_n10918# 0.146647f
C78 a_n118_n10788# a_n746_n10918# 0.17691f
C79 a_n118_n6988# a_n746_n10918# 0.146647f
C80 a_n284_n10788# a_n746_n10918# 0.17691f
C81 a_n284_n6988# a_n746_n10918# 0.146647f
C82 a_n450_n10788# a_n746_n10918# 0.17691f
C83 a_n450_n6988# a_n746_n10918# 0.146647f
C84 a_n616_n10788# a_n746_n10918# 0.387223f
C85 a_n616_n6988# a_n746_n10918# 0.356961f
C86 a_546_n6452# a_n746_n10918# 0.356961f
C87 a_546_n2652# a_n746_n10918# 0.356961f
C88 a_380_n6452# a_n746_n10918# 0.146647f
C89 a_380_n2652# a_n746_n10918# 0.146647f
C90 a_214_n6452# a_n746_n10918# 0.146647f
C91 a_214_n2652# a_n746_n10918# 0.146647f
C92 a_48_n6452# a_n746_n10918# 0.146647f
C93 a_48_n2652# a_n746_n10918# 0.146647f
C94 a_n118_n6452# a_n746_n10918# 0.146647f
C95 a_n118_n2652# a_n746_n10918# 0.146647f
C96 a_n284_n6452# a_n746_n10918# 0.146647f
C97 a_n284_n2652# a_n746_n10918# 0.146647f
C98 a_n450_n6452# a_n746_n10918# 0.146647f
C99 a_n450_n2652# a_n746_n10918# 0.146647f
C100 a_n616_n6452# a_n746_n10918# 0.356961f
C101 a_n616_n2652# a_n746_n10918# 0.356961f
C102 a_546_n2116# a_n746_n10918# 0.356961f
C103 a_546_1684# a_n746_n10918# 0.356961f
C104 a_380_n2116# a_n746_n10918# 0.146647f
C105 a_380_1684# a_n746_n10918# 0.146647f
C106 a_214_n2116# a_n746_n10918# 0.146647f
C107 a_214_1684# a_n746_n10918# 0.146647f
C108 a_48_n2116# a_n746_n10918# 0.146647f
C109 a_48_1684# a_n746_n10918# 0.146647f
C110 a_n118_n2116# a_n746_n10918# 0.146647f
C111 a_n118_1684# a_n746_n10918# 0.146647f
C112 a_n284_n2116# a_n746_n10918# 0.146647f
C113 a_n284_1684# a_n746_n10918# 0.146647f
C114 a_n450_n2116# a_n746_n10918# 0.146647f
C115 a_n450_1684# a_n746_n10918# 0.146647f
C116 a_n616_n2116# a_n746_n10918# 0.356961f
C117 a_n616_1684# a_n746_n10918# 0.356961f
C118 a_546_2220# a_n746_n10918# 0.356961f
C119 a_546_6020# a_n746_n10918# 0.356961f
C120 a_380_2220# a_n746_n10918# 0.146647f
C121 a_380_6020# a_n746_n10918# 0.146647f
C122 a_214_2220# a_n746_n10918# 0.146647f
C123 a_214_6020# a_n746_n10918# 0.146647f
C124 a_48_2220# a_n746_n10918# 0.146647f
C125 a_48_6020# a_n746_n10918# 0.146647f
C126 a_n118_2220# a_n746_n10918# 0.146647f
C127 a_n118_6020# a_n746_n10918# 0.146647f
C128 a_n284_2220# a_n746_n10918# 0.146647f
C129 a_n284_6020# a_n746_n10918# 0.146647f
C130 a_n450_2220# a_n746_n10918# 0.146647f
C131 a_n450_6020# a_n746_n10918# 0.146647f
C132 a_n616_2220# a_n746_n10918# 0.356961f
C133 a_n616_6020# a_n746_n10918# 0.356961f
C134 a_546_6556# a_n746_n10918# 0.356961f
C135 a_546_10356# a_n746_n10918# 0.387223f
C136 a_380_6556# a_n746_n10918# 0.146647f
C137 a_380_10356# a_n746_n10918# 0.17691f
C138 a_214_6556# a_n746_n10918# 0.146647f
C139 a_214_10356# a_n746_n10918# 0.17691f
C140 a_48_6556# a_n746_n10918# 0.146647f
C141 a_48_10356# a_n746_n10918# 0.17691f
C142 a_n118_6556# a_n746_n10918# 0.146647f
C143 a_n118_10356# a_n746_n10918# 0.17691f
C144 a_n284_6556# a_n746_n10918# 0.146647f
C145 a_n284_10356# a_n746_n10918# 0.17691f
C146 a_n450_6556# a_n746_n10918# 0.146647f
C147 a_n450_10356# a_n746_n10918# 0.17691f
C148 a_n616_6556# a_n746_n10918# 0.356961f
C149 a_n616_10356# a_n746_n10918# 0.387223f
.ends

.subckt resistorstart B AVSS A
Xsky130_fd_pr__res_high_po_0p35_9NXREG_0 m1_8663_1119# m1_8663_787# m1_4327_1119#
+ m1_12999_1285# m1_17335_1285# m1_119_456# m1_4327_953# m1_17335_455# m1_8663_123#
+ m1_4327_123# m1_17335_123# m1_21633_953# m1_8663_953# m1_12999_455# m1_12999_1119#
+ m1_17335_455# m1_4327_953# m1_8663_1285# m1_12999_123# AVSS m1_4327_787# m1_17335_123#
+ A m1_17335_621# AVSS m1_8663_787# m1_4327_787# m1_12999_289# m1_8663_289# m1_12999_621#
+ m1_12999_953# m1_17335_621# m1_4327_1285# m1_21633_289# B m1_119_788# m1_8663_455#
+ m1_17335_1119# m1_21633_953# m1_8663_1285# m1_4327_1285# m1_21633_621# m1_12999_1119#
+ m1_4327_289# m1_12999_787# m1_17335_1119# m1_8663_621# m1_17335_289# m1_119_788#
+ m1_8663_289# m1_17335_953# m1_4327_455# m1_4327_289# m1_12999_1285# m1_12999_289#
+ m1_17335_289# m1_8663_455# m1_8663_1119# m1_12999_953# AVSS m1_17335_953# m1_4327_455#
+ m1_4327_621# m1_8663_123# m1_12999_455# m1_17335_787# m1_21633_289# m1_12999_123#
+ m1_119_456# AVSS m1_8663_621# m1_8663_953# m1_4327_621# AVSS m1_12999_787# m1_17335_787#
+ m1_4327_1119# m1_17335_1285# m1_4327_123# m1_12999_621# m1_21633_621# sky130_fd_pr__res_high_po_0p35_9NXREG
C0 m1_21633_953# AVSS 0.423941f
C1 m1_21633_621# AVSS 0.423825f
C2 m1_21633_289# AVSS 0.42396f
C3 m1_17335_1285# AVSS 0.855996f
C4 m1_17335_1119# AVSS 0.301698f
C5 m1_17335_953# AVSS 0.301628f
C6 m1_17335_787# AVSS 0.30161f
C7 m1_17335_621# AVSS 0.30161f
C8 m1_17335_455# AVSS 0.301628f
C9 m1_17335_289# AVSS 0.301698f
C10 m1_17335_123# AVSS 0.855995f
C11 m1_12999_1285# AVSS 0.855996f
C12 m1_12999_1119# AVSS 0.301698f
C13 m1_12999_953# AVSS 0.301628f
C14 m1_12999_787# AVSS 0.30161f
C15 m1_12999_621# AVSS 0.30161f
C16 m1_12999_455# AVSS 0.301628f
C17 m1_12999_289# AVSS 0.301698f
C18 m1_12999_123# AVSS 0.855995f
C19 m1_8663_1285# AVSS 0.855996f
C20 m1_8663_1119# AVSS 0.301698f
C21 m1_8663_953# AVSS 0.301628f
C22 m1_8663_787# AVSS 0.30161f
C23 m1_8663_621# AVSS 0.30161f
C24 m1_8663_455# AVSS 0.301628f
C25 m1_8663_289# AVSS 0.301698f
C26 m1_8663_123# AVSS 0.855996f
C27 m1_4327_1285# AVSS 0.855995f
C28 m1_4327_1119# AVSS 0.301698f
C29 A AVSS 0.185367f
C30 m1_4327_953# AVSS 0.301628f
C31 m1_119_788# AVSS 0.424053f
C32 m1_4327_787# AVSS 0.30161f
C33 m1_4327_621# AVSS 0.30161f
C34 m1_119_456# AVSS 0.424053f
C35 m1_4327_455# AVSS 0.301628f
C36 m1_4327_289# AVSS 0.301698f
C37 B AVSS 0.185367f
C38 m1_4327_123# AVSS 0.855996f
.ends

.subckt sky130_fd_pr__pfet_01v8_CVRJBD a_n2029_n128# a_2029_n64# a_29_n128# a_n2087_n64#
+ w_n2123_n164# a_n29_n64# VSUBS
X0 a_2029_n64# a_29_n128# a_n29_n64# w_n2123_n164# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=10
X1 a_n29_n64# a_n2029_n128# a_n2087_n64# w_n2123_n164# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=10
C0 w_n2123_n164# a_29_n128# 0.823465f
C1 w_n2123_n164# a_n2029_n128# 0.823465f
C2 a_2029_n64# VSUBS 0.149664f
C3 a_n29_n64# VSUBS 0.112935f
C4 a_n2087_n64# VSUBS 0.149664f
C5 a_29_n128# VSUBS 2.76013f
C6 a_n2029_n128# VSUBS 2.76013f
C7 w_n2123_n164# VSUBS 4.61116f
.ends

.subckt sky130_fd_pr__pfet_01v8_8RMJP2 a_n2029_n162# a_n2087_n136# w_n2123_n198# a_29_n162#
+ a_2029_n136# a_n29_n136# VSUBS
X0 a_2029_n136# a_29_n162# a_n29_n136# w_n2123_n198# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=10
X1 a_n29_n136# a_n2029_n162# a_n2087_n136# w_n2123_n198# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=10
C0 w_n2123_n198# a_29_n162# 0.823465f
C1 w_n2123_n198# a_n2029_n162# 0.823465f
C2 a_2029_n136# VSUBS 0.149664f
C3 a_n29_n136# VSUBS 0.112935f
C4 a_n2087_n136# VSUBS 0.149664f
C5 a_29_n162# VSUBS 2.76013f
C6 a_n2029_n162# VSUBS 2.76013f
C7 w_n2123_n198# VSUBS 4.61116f
.ends

.subckt sky130_fd_pr__pfet_01v8_2XUZHN a_n73_n100# w_n109_n162# a_15_n100# a_n15_n126#
+ VSUBS
X0 a_15_n100# a_n15_n126# a_n73_n100# w_n109_n162# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
C0 a_15_n100# a_n73_n100# 0.162113f
C1 a_15_n100# VSUBS 0.111398f
C2 a_n73_n100# VSUBS 0.111398f
C3 w_n109_n162# VSUBS 0.211896f
.ends

.subckt pmos_iptat VDDE D G
Xsky130_fd_pr__pfet_01v8_CVRJBD_1 G D G D VDDE VDDE VSUBS sky130_fd_pr__pfet_01v8_CVRJBD
Xsky130_fd_pr__pfet_01v8_8RMJP2_0 G D VDDE G D VDDE VSUBS sky130_fd_pr__pfet_01v8_8RMJP2
Xsky130_fd_pr__pfet_01v8_2XUZHN_0 D VDDE D D VSUBS sky130_fd_pr__pfet_01v8_2XUZHN
Xsky130_fd_pr__pfet_01v8_2XUZHN_2 D VDDE D D VSUBS sky130_fd_pr__pfet_01v8_2XUZHN
Xsky130_fd_pr__pfet_01v8_2XUZHN_3 D VDDE D D VSUBS sky130_fd_pr__pfet_01v8_2XUZHN
Xsky130_fd_pr__pfet_01v8_2XUZHN_4 D VDDE D D VSUBS sky130_fd_pr__pfet_01v8_2XUZHN
C0 VDDE D 1.599952f
C1 D G 2.061433f
C2 VDDE G 6.186075f
C3 D VSUBS 0.36973f
C4 G VSUBS 5.93504f
C5 VDDE VSUBS 18.917078f
.ends

.subckt sky130_fd_pr__pfet_01v8_2ZH9EN a_15_n200# a_n15_n226# a_n73_n200# w_n109_n262#
+ VSUBS
X0 a_15_n200# a_n15_n226# a_n73_n200# w_n109_n262# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
C0 a_n73_n200# a_15_n200# 0.321048f
C1 a_15_n200# VSUBS 0.193584f
C2 a_n73_n200# VSUBS 0.193584f
C3 w_n109_n262# VSUBS 0.342696f
.ends

.subckt sky130_fd_pr__pfet_01v8_CVH45E a_n429_n228# w_n523_n264# a_29_n228# a_n487_n164#
+ a_n29_n164# a_429_n164# VSUBS
X0 a_429_n164# a_29_n228# a_n29_n164# w_n523_n264# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=2
X1 a_n29_n164# a_n429_n228# a_n487_n164# w_n523_n264# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=2
C0 a_29_n228# w_n523_n264# 0.19694f
C1 a_n429_n228# w_n523_n264# 0.19694f
C2 a_429_n164# VSUBS 0.226031f
C3 a_n29_n164# VSUBS 0.108699f
C4 a_n487_n164# VSUBS 0.226031f
C5 a_29_n228# VSUBS 0.571505f
C6 a_n429_n228# VSUBS 0.571505f
C7 w_n523_n264# VSUBS 1.76356f
.ends

.subckt sky130_fd_pr__pfet_01v8_9XC4R9 a_n429_n262# a_29_n262# a_n487_n236# a_n29_n236#
+ a_429_n236# w_n523_n298# VSUBS
X0 a_n29_n236# a_n429_n262# a_n487_n236# w_n523_n298# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=2
X1 a_429_n236# a_29_n262# a_n29_n236# w_n523_n298# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=2
C0 a_29_n262# w_n523_n298# 0.19694f
C1 a_n429_n262# w_n523_n298# 0.19694f
C2 a_429_n236# VSUBS 0.226031f
C3 a_n29_n236# VSUBS 0.108699f
C4 a_n487_n236# VSUBS 0.226031f
C5 a_29_n262# VSUBS 0.571505f
C6 a_n429_n262# VSUBS 0.571505f
C7 w_n523_n298# VSUBS 1.76356f
.ends

.subckt pmos_ena G AVDD DVDD VDDE
Xsky130_fd_pr__pfet_01v8_2ZH9EN_0 VDDE VDDE VDDE DVDD VSUBS sky130_fd_pr__pfet_01v8_2ZH9EN
Xsky130_fd_pr__pfet_01v8_2ZH9EN_1 VDDE VDDE VDDE DVDD VSUBS sky130_fd_pr__pfet_01v8_2ZH9EN
Xsky130_fd_pr__pfet_01v8_2ZH9EN_2 VDDE VDDE VDDE DVDD VSUBS sky130_fd_pr__pfet_01v8_2ZH9EN
Xsky130_fd_pr__pfet_01v8_2ZH9EN_3 VDDE VDDE VDDE DVDD VSUBS sky130_fd_pr__pfet_01v8_2ZH9EN
Xsky130_fd_pr__pfet_01v8_CVH45E_0 G DVDD G VDDE AVDD VDDE VSUBS sky130_fd_pr__pfet_01v8_CVH45E
Xsky130_fd_pr__pfet_01v8_9XC4R9_0 G G VDDE AVDD VDDE DVDD VSUBS sky130_fd_pr__pfet_01v8_9XC4R9
C0 AVDD G 0.158408f
C1 DVDD G 0.959425f
C2 AVDD VDDE 0.108893f
C3 G VDDE 0.616455f
C4 DVDD VDDE 0.845523f
C5 AVDD VSUBS 0.502599f
C6 VDDE VSUBS 0.804754f
C7 G VSUBS 1.479204f
C8 DVDD VSUBS 7.209626f
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_UG4D4N a_29_n457# a_n287_n369# a_n229_n457# a_229_n369#
+ a_n29_n369# VSUBS
X0 a_n29_n369# a_n229_n457# a_n287_n369# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=1
X1 a_229_n369# a_29_n457# a_n29_n369# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=1
C0 a_n287_n369# a_n29_n369# 0.219309f
C1 a_229_n369# a_n29_n369# 0.219309f
C2 a_229_n369# VSUBS 0.41069f
C3 a_n29_n369# VSUBS 0.138774f
C4 a_n287_n369# VSUBS 0.41069f
C5 a_29_n457# VSUBS 0.46679f
C6 a_n229_n457# VSUBS 0.46679f
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_TGDTCU a_n287_n431# a_29_n457# a_229_n431# a_n229_n457#
+ a_n29_n431# VSUBS
X0 a_n29_n431# a_n229_n457# a_n287_n431# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=1
X1 a_229_n431# a_29_n457# a_n29_n431# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=1
C0 a_n287_n431# a_n29_n431# 0.219309f
C1 a_229_n431# a_n29_n431# 0.219309f
C2 a_229_n431# VSUBS 0.41069f
C3 a_n29_n431# VSUBS 0.138774f
C4 a_n287_n431# VSUBS 0.41069f
C5 a_29_n457# VSUBS 0.46679f
C6 a_n229_n457# VSUBS 0.46679f
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_QJFS9J a_n73_n400# a_15_n400# a_n15_n426# VSUBS
X0 a_15_n400# a_n15_n426# a_n73_n400# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.15
C0 a_n73_n400# a_15_n400# 0.638918f
C1 a_15_n400# VSUBS 0.372089f
C2 a_n73_n400# VSUBS 0.372089f
.ends

.subckt trim S D DVSS G
Xsky130_fd_pr__nfet_01v8_lvt_UG4D4N_0 G D G D S DVSS sky130_fd_pr__nfet_01v8_lvt_UG4D4N
Xsky130_fd_pr__nfet_01v8_lvt_TGDTCU_0 D G D G S DVSS sky130_fd_pr__nfet_01v8_lvt_TGDTCU
Xsky130_fd_pr__nfet_01v8_lvt_QJFS9J_0 D D D DVSS sky130_fd_pr__nfet_01v8_lvt_QJFS9J
Xsky130_fd_pr__nfet_01v8_lvt_QJFS9J_1 D D D DVSS sky130_fd_pr__nfet_01v8_lvt_QJFS9J
Xsky130_fd_pr__nfet_01v8_lvt_QJFS9J_2 D D D DVSS sky130_fd_pr__nfet_01v8_lvt_QJFS9J
Xsky130_fd_pr__nfet_01v8_lvt_QJFS9J_3 D D D DVSS sky130_fd_pr__nfet_01v8_lvt_QJFS9J
C0 G S 0.15958f
C1 D S 0.145154f
C2 D G 0.403123f
C3 S DVSS 0.898422f
C4 D DVSS 2.777826f
C5 G DVSS 2.000921f
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_SJFSNB a_n73_n100# a_15_n100# a_n15_n126# VSUBS
X0 a_15_n100# a_n15_n126# a_n73_n100# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
C0 a_15_n100# a_n73_n100# 0.162113f
C1 a_15_n100# VSUBS 0.118371f
C2 a_n73_n100# VSUBS 0.118371f
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_U8VHVM a_n287_n131# a_29_n157# a_229_n131# a_n229_n157#
+ a_n29_n131# VSUBS
X0 a_229_n131# a_29_n157# a_n29_n131# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X1 a_n29_n131# a_n229_n157# a_n287_n131# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
C0 a_229_n131# VSUBS 0.127112f
C1 a_n287_n131# VSUBS 0.127112f
C2 a_29_n157# VSUBS 0.482705f
C3 a_n229_n157# VSUBS 0.482705f
.ends

.subckt vena G D S DVSS
Xsky130_fd_pr__nfet_01v8_lvt_SJFSNB_1 D D D DVSS sky130_fd_pr__nfet_01v8_lvt_SJFSNB
Xsky130_fd_pr__nfet_01v8_lvt_SJFSNB_2 D D D DVSS sky130_fd_pr__nfet_01v8_lvt_SJFSNB
Xsky130_fd_pr__nfet_01v8_lvt_U8VHVM_0 D G D G S DVSS sky130_fd_pr__nfet_01v8_lvt_U8VHVM
C0 D G 0.151015f
C1 D DVSS 0.982002f
C2 G DVSS 0.985505f
.ends

.subckt digital S3 D3 trim3 S2 trim2 trim1 trim0 S1 S0 VENA VBGTC SVBGSC SVBGTC AVDD
+ ENA DVDD DVSS VBGSC VDDE
Xpmos_ena_0 ENA AVDD DVDD VDDE pmos_ena
Xtrim_0 S3 D3 DVSS trim3 trim
Xtrim_1 S2 S3 DVSS trim2 trim
Xtrim_2 S1 S2 DVSS trim1 trim
Xtrim_3 S0 S1 DVSS trim0 trim
Xvena_0 VENA VBGTC SVBGTC DVSS vena
Xvena_1 VENA VBGSC SVBGSC DVSS vena
C0 S1 S2 0.651596f
C1 VBGSC S1 0.120014f
C2 S1 S0 0.104801f
C3 S3 S2 0.651595f
C4 DVDD trim3 0.146413f
C5 trim1 DVDD 0.139521f
C6 D3 DVDD 0.145467f
C7 DVDD ENA 0.121406f
C8 VENA ENA 0.147211f
C9 S1 VBGTC 0.120014f
C10 trim2 DVDD 0.139521f
C11 DVDD trim0 0.139521f
C12 D3 S3 0.546794f
C13 VENA DVDD 0.159829f
C14 VBGSC VSUBS 0.64886f
C15 VENA VSUBS 1.483952f
C16 VBGTC VSUBS 0.648859f
C17 S0 VSUBS 0.74708f
C18 S1 VSUBS 1.926616f
C19 trim0 VSUBS 1.504461f
C20 S2 VSUBS 1.850228f
C21 trim1 VSUBS 1.492518f
C22 S3 VSUBS 1.980663f
C23 trim2 VSUBS 1.49252f
C24 D3 VSUBS 1.269093f
C25 trim3 VSUBS 1.498829f
C26 AVDD VSUBS 0.490888f
C27 VDDE VSUBS 0.685901f
C28 ENA VSUBS 1.253672f
C29 DVDD VSUBS 90.219315f
.ends

.subckt pmos_startup D3 D4 VDDE D2
Xsky130_fd_pr__pfet_01v8_CVRJBD_1 D3 D2 D3 D3 VDDE VDDE VSUBS sky130_fd_pr__pfet_01v8_CVRJBD
Xsky130_fd_pr__pfet_01v8_8RMJP2_0 D2 D4 VDDE VDDE VDDE VDDE VSUBS sky130_fd_pr__pfet_01v8_8RMJP2
Xsky130_fd_pr__pfet_01v8_2XUZHN_0 D2 VDDE D2 D2 VSUBS sky130_fd_pr__pfet_01v8_2XUZHN
Xsky130_fd_pr__pfet_01v8_2XUZHN_1 VDDE VDDE VDDE VDDE VSUBS sky130_fd_pr__pfet_01v8_2XUZHN
Xsky130_fd_pr__pfet_01v8_2XUZHN_2 D3 VDDE D3 D3 VSUBS sky130_fd_pr__pfet_01v8_2XUZHN
Xsky130_fd_pr__pfet_01v8_2XUZHN_4 D4 VDDE D4 D4 VSUBS sky130_fd_pr__pfet_01v8_2XUZHN
C0 D2 VDDE 2.915652f
C1 VDDE D4 0.371001f
C2 D3 D2 2.154161f
C3 D3 VDDE 3.062172f
C4 D2 VSUBS 1.596815f
C5 D3 VSUBS 3.08946f
C6 VDDE VSUBS 18.958673f
.ends

.subckt sky130_fd_pr__res_high_po_0p35_KQ9YC9 a_n616_2132# a_n284_5284# a_380_n5716#
+ a_380_2668# a_214_2132# a_n284_n2564# a_n118_4748# a_48_n5180# a_n616_2668# a_n450_7364#
+ a_380_n484# a_48_n3100# a_n616_n2564# a_n118_5284# a_n616_n484# a_n450_n7796# a_214_2668#
+ a_214_n7796# a_n450_n5716# a_n284_7364# a_546_n5180# a_48_2132# a_214_n5716# a_380_4748#
+ a_214_n484# a_546_n3100# a_n746_n7926# a_n118_n2564# a_n616_4748# a_48_52# a_380_5284#
+ a_n616_52# a_48_2668# a_n284_n5180# a_n118_7364# a_n616_5284# a_546_52# a_n284_n3100#
+ a_214_4748# a_48_n7796# a_546_2132# a_n616_n5180# a_48_n484# a_48_n5716# a_n616_n3100#
+ a_214_5284# a_380_n2564# a_546_2668# a_380_7364# a_546_n7796# a_48_4748# a_n118_n5180#
+ a_546_n5716# a_n616_7364# a_546_n484# a_n450_2132# a_n118_n3100# a_48_5284# a_n284_n7796#
+ a_214_7364# a_n450_n2564# a_n450_52# a_214_n2564# a_n284_2132# a_n284_n5716# a_n450_2668#
+ a_546_4748# a_n616_n7796# a_380_52# a_n616_n5716# a_n284_52# a_380_n5180# a_214_52#
+ a_n450_n484# a_546_5284# a_380_n3100# a_n118_52# a_n284_2668# a_48_7364# a_n118_2132#
+ a_n118_n7796# a_n284_n484# a_48_n2564# a_n450_4748# a_n118_n5716# a_n450_n5180#
+ a_n118_2668# a_214_n5180# a_n450_n3100# a_n450_5284# a_546_7364# a_214_n3100# a_n284_4748#
+ a_380_2132# a_546_n2564# a_n118_n484# a_380_n7796#
X0 a_n616_n5716# a_n616_n7796# a_n746_n7926# sky130_fd_pr__res_high_po_0p35 l=8.4
X1 a_n616_n484# a_n616_n2564# a_n746_n7926# sky130_fd_pr__res_high_po_0p35 l=8.4
X2 a_214_7364# a_214_5284# a_n746_n7926# sky130_fd_pr__res_high_po_0p35 l=8.4
X3 a_546_4748# a_546_2668# a_n746_n7926# sky130_fd_pr__res_high_po_0p35 l=8.4
X4 a_380_n5716# a_380_n7796# a_n746_n7926# sky130_fd_pr__res_high_po_0p35 l=8.4
X5 a_546_n5716# a_546_n7796# a_n746_n7926# sky130_fd_pr__res_high_po_0p35 l=8.4
X6 a_n284_7364# a_n284_5284# a_n746_n7926# sky130_fd_pr__res_high_po_0p35 l=8.4
X7 a_380_n484# a_380_n2564# a_n746_n7926# sky130_fd_pr__res_high_po_0p35 l=8.4
X8 a_546_n484# a_546_n2564# a_n746_n7926# sky130_fd_pr__res_high_po_0p35 l=8.4
X9 a_n450_n3100# a_n450_n5180# a_n746_n7926# sky130_fd_pr__res_high_po_0p35 l=8.4
X10 a_n284_n3100# a_n284_n5180# a_n746_n7926# sky130_fd_pr__res_high_po_0p35 l=8.4
X11 a_n118_2132# a_n118_52# a_n746_n7926# sky130_fd_pr__res_high_po_0p35 l=8.4
X12 a_48_2132# a_48_52# a_n746_n7926# sky130_fd_pr__res_high_po_0p35 l=8.4
X13 a_48_n3100# a_48_n5180# a_n746_n7926# sky130_fd_pr__res_high_po_0p35 l=8.4
X14 a_214_4748# a_214_2668# a_n746_n7926# sky130_fd_pr__res_high_po_0p35 l=8.4
X15 a_214_2132# a_214_52# a_n746_n7926# sky130_fd_pr__res_high_po_0p35 l=8.4
X16 a_n450_7364# a_n450_5284# a_n746_n7926# sky130_fd_pr__res_high_po_0p35 l=8.4
X17 a_48_7364# a_48_5284# a_n746_n7926# sky130_fd_pr__res_high_po_0p35 l=8.4
X18 a_n450_n5716# a_n450_n7796# a_n746_n7926# sky130_fd_pr__res_high_po_0p35 l=8.4
X19 a_n284_n5716# a_n284_n7796# a_n746_n7926# sky130_fd_pr__res_high_po_0p35 l=8.4
X20 a_n284_4748# a_n284_2668# a_n746_n7926# sky130_fd_pr__res_high_po_0p35 l=8.4
X21 a_n616_2132# a_n616_52# a_n746_n7926# sky130_fd_pr__res_high_po_0p35 l=8.4
X22 a_n450_n484# a_n450_n2564# a_n746_n7926# sky130_fd_pr__res_high_po_0p35 l=8.4
X23 a_n284_n484# a_n284_n2564# a_n746_n7926# sky130_fd_pr__res_high_po_0p35 l=8.4
X24 a_48_n5716# a_48_n7796# a_n746_n7926# sky130_fd_pr__res_high_po_0p35 l=8.4
X25 a_n284_2132# a_n284_52# a_n746_n7926# sky130_fd_pr__res_high_po_0p35 l=8.4
X26 a_48_n484# a_48_n2564# a_n746_n7926# sky130_fd_pr__res_high_po_0p35 l=8.4
X27 a_n118_7364# a_n118_5284# a_n746_n7926# sky130_fd_pr__res_high_po_0p35 l=8.4
X28 a_380_2132# a_380_52# a_n746_n7926# sky130_fd_pr__res_high_po_0p35 l=8.4
X29 a_48_4748# a_48_2668# a_n746_n7926# sky130_fd_pr__res_high_po_0p35 l=8.4
X30 a_n450_4748# a_n450_2668# a_n746_n7926# sky130_fd_pr__res_high_po_0p35 l=8.4
X31 a_214_n3100# a_214_n5180# a_n746_n7926# sky130_fd_pr__res_high_po_0p35 l=8.4
X32 a_n118_4748# a_n118_2668# a_n746_n7926# sky130_fd_pr__res_high_po_0p35 l=8.4
X33 a_214_n5716# a_214_n7796# a_n746_n7926# sky130_fd_pr__res_high_po_0p35 l=8.4
X34 a_n616_7364# a_n616_5284# a_n746_n7926# sky130_fd_pr__res_high_po_0p35 l=8.4
X35 a_214_n484# a_214_n2564# a_n746_n7926# sky130_fd_pr__res_high_po_0p35 l=8.4
X36 a_n118_n3100# a_n118_n5180# a_n746_n7926# sky130_fd_pr__res_high_po_0p35 l=8.4
X37 a_380_7364# a_380_5284# a_n746_n7926# sky130_fd_pr__res_high_po_0p35 l=8.4
X38 a_n450_2132# a_n450_52# a_n746_n7926# sky130_fd_pr__res_high_po_0p35 l=8.4
X39 a_n616_n3100# a_n616_n5180# a_n746_n7926# sky130_fd_pr__res_high_po_0p35 l=8.4
X40 a_n118_n5716# a_n118_n7796# a_n746_n7926# sky130_fd_pr__res_high_po_0p35 l=8.4
X41 a_546_7364# a_546_5284# a_n746_n7926# sky130_fd_pr__res_high_po_0p35 l=8.4
X42 a_n118_n484# a_n118_n2564# a_n746_n7926# sky130_fd_pr__res_high_po_0p35 l=8.4
X43 a_n616_4748# a_n616_2668# a_n746_n7926# sky130_fd_pr__res_high_po_0p35 l=8.4
X44 a_380_4748# a_380_2668# a_n746_n7926# sky130_fd_pr__res_high_po_0p35 l=8.4
X45 a_546_2132# a_546_52# a_n746_n7926# sky130_fd_pr__res_high_po_0p35 l=8.4
X46 a_380_n3100# a_380_n5180# a_n746_n7926# sky130_fd_pr__res_high_po_0p35 l=8.4
X47 a_546_n3100# a_546_n5180# a_n746_n7926# sky130_fd_pr__res_high_po_0p35 l=8.4
C0 a_n118_n5716# a_48_n5716# 0.296258f
C1 a_n118_2668# a_48_2668# 0.296258f
C2 a_n118_n5180# a_48_n5180# 0.296258f
C3 a_n118_2132# a_n284_2132# 0.296258f
C4 a_n118_52# a_48_52# 0.296258f
C5 a_n284_n3100# a_n118_n3100# 0.296258f
C6 a_380_5284# a_214_5284# 0.296258f
C7 a_n450_n7796# a_n284_n7796# 0.296258f
C8 a_n616_7364# a_n450_7364# 0.296258f
C9 a_n118_n5716# a_n284_n5716# 0.296258f
C10 a_n284_2668# a_n450_2668# 0.296258f
C11 a_n616_n5180# a_n450_n5180# 0.296258f
C12 a_546_n5716# a_380_n5716# 0.296258f
C13 a_214_2668# a_380_2668# 0.296258f
C14 a_214_n5180# a_380_n5180# 0.296258f
C15 a_48_4748# a_214_4748# 0.296258f
C16 a_n118_n2564# a_48_n2564# 0.296258f
C17 a_n284_4748# a_n450_4748# 0.296258f
C18 a_380_n2564# a_546_n2564# 0.296258f
C19 a_48_2132# a_214_2132# 0.296258f
C20 a_n118_5284# a_48_5284# 0.296258f
C21 a_48_n3100# a_n118_n3100# 0.296258f
C22 a_n616_5284# a_n450_5284# 0.296258f
C23 a_48_2132# a_n118_2132# 0.296258f
C24 a_n450_n2564# a_n284_n2564# 0.296258f
C25 a_48_4748# a_n118_4748# 0.296258f
C26 a_n284_7364# a_n450_7364# 0.296258f
C27 a_546_7364# a_380_7364# 0.296258f
C28 a_48_n7796# a_n118_n7796# 0.296258f
C29 a_48_n7796# a_214_n7796# 0.296258f
C30 a_380_n2564# a_214_n2564# 0.296258f
C31 a_380_n484# a_546_n484# 0.296258f
C32 a_n616_52# a_n450_52# 0.296258f
C33 a_n450_2132# a_n616_2132# 0.296258f
C34 a_48_n5716# a_214_n5716# 0.296258f
C35 a_380_n7796# a_214_n7796# 0.296258f
C36 a_n118_5284# a_n284_5284# 0.296258f
C37 a_380_n7796# a_546_n7796# 0.296258f
C38 a_546_n5180# a_380_n5180# 0.296258f
C39 a_214_52# a_48_52# 0.296258f
C40 a_214_n5180# a_48_n5180# 0.296258f
C41 a_214_n3100# a_48_n3100# 0.296258f
C42 a_n616_2668# a_n450_2668# 0.296258f
C43 a_n118_n2564# a_n284_n2564# 0.296258f
C44 a_n284_7364# a_n118_7364# 0.296258f
C45 a_n284_n5180# a_n118_n5180# 0.296258f
C46 a_n284_52# a_n118_52# 0.296258f
C47 a_380_n484# a_214_n484# 0.296258f
C48 a_n118_7364# a_48_7364# 0.296258f
C49 a_n284_n5180# a_n450_n5180# 0.296258f
C50 a_n616_n5716# a_n450_n5716# 0.296258f
C51 a_n616_n484# a_n450_n484# 0.296258f
C52 a_546_2132# a_380_2132# 0.296258f
C53 a_n284_n484# a_n118_n484# 0.296258f
C54 a_n616_n3100# a_n450_n3100# 0.296258f
C55 a_48_5284# a_214_5284# 0.296258f
C56 a_380_n3100# a_546_n3100# 0.296258f
C57 a_214_n3100# a_380_n3100# 0.296258f
C58 a_546_52# a_380_52# 0.296258f
C59 a_214_2132# a_380_2132# 0.296258f
C60 a_214_2668# a_48_2668# 0.296258f
C61 a_n284_5284# a_n450_5284# 0.296258f
C62 a_n284_52# a_n450_52# 0.296258f
C63 a_n118_2668# a_n284_2668# 0.296258f
C64 a_n284_n3100# a_n450_n3100# 0.296258f
C65 a_n450_2132# a_n284_2132# 0.296258f
C66 a_n450_4748# a_n616_4748# 0.296258f
C67 a_n284_n484# a_n450_n484# 0.296258f
C68 a_n284_n5716# a_n450_n5716# 0.296258f
C69 a_48_n484# a_n118_n484# 0.296258f
C70 a_380_4748# a_546_4748# 0.296258f
C71 a_214_7364# a_380_7364# 0.296258f
C72 a_380_4748# a_214_4748# 0.296258f
C73 a_n450_n2564# a_n616_n2564# 0.296258f
C74 a_n284_n7796# a_n118_n7796# 0.296258f
C75 a_214_7364# a_48_7364# 0.296258f
C76 a_546_2668# a_380_2668# 0.296258f
C77 a_380_5284# a_546_5284# 0.296258f
C78 a_48_n484# a_214_n484# 0.296258f
C79 a_n450_n7796# a_n616_n7796# 0.296258f
C80 a_214_n5716# a_380_n5716# 0.296258f
C81 a_214_52# a_380_52# 0.296258f
C82 a_n284_4748# a_n118_4748# 0.296258f
C83 a_48_n2564# a_214_n2564# 0.296258f
C84 a_546_n7796# a_n746_n7926# 0.387223f
C85 a_546_n5716# a_n746_n7926# 0.356961f
C86 a_380_n7796# a_n746_n7926# 0.17691f
C87 a_380_n5716# a_n746_n7926# 0.146647f
C88 a_214_n7796# a_n746_n7926# 0.17691f
C89 a_214_n5716# a_n746_n7926# 0.146647f
C90 a_48_n7796# a_n746_n7926# 0.17691f
C91 a_48_n5716# a_n746_n7926# 0.146647f
C92 a_n118_n7796# a_n746_n7926# 0.17691f
C93 a_n118_n5716# a_n746_n7926# 0.146647f
C94 a_n284_n7796# a_n746_n7926# 0.17691f
C95 a_n284_n5716# a_n746_n7926# 0.146647f
C96 a_n450_n7796# a_n746_n7926# 0.17691f
C97 a_n450_n5716# a_n746_n7926# 0.146647f
C98 a_n616_n7796# a_n746_n7926# 0.387223f
C99 a_n616_n5716# a_n746_n7926# 0.356961f
C100 a_546_n5180# a_n746_n7926# 0.356961f
C101 a_546_n3100# a_n746_n7926# 0.356961f
C102 a_380_n5180# a_n746_n7926# 0.146647f
C103 a_380_n3100# a_n746_n7926# 0.146647f
C104 a_214_n5180# a_n746_n7926# 0.146647f
C105 a_214_n3100# a_n746_n7926# 0.146647f
C106 a_48_n5180# a_n746_n7926# 0.146647f
C107 a_48_n3100# a_n746_n7926# 0.146647f
C108 a_n118_n5180# a_n746_n7926# 0.146647f
C109 a_n118_n3100# a_n746_n7926# 0.146647f
C110 a_n284_n5180# a_n746_n7926# 0.146647f
C111 a_n284_n3100# a_n746_n7926# 0.146647f
C112 a_n450_n5180# a_n746_n7926# 0.146647f
C113 a_n450_n3100# a_n746_n7926# 0.146647f
C114 a_n616_n5180# a_n746_n7926# 0.356961f
C115 a_n616_n3100# a_n746_n7926# 0.356961f
C116 a_546_n2564# a_n746_n7926# 0.356961f
C117 a_546_n484# a_n746_n7926# 0.356961f
C118 a_380_n2564# a_n746_n7926# 0.146647f
C119 a_380_n484# a_n746_n7926# 0.146647f
C120 a_214_n2564# a_n746_n7926# 0.146647f
C121 a_214_n484# a_n746_n7926# 0.146647f
C122 a_48_n2564# a_n746_n7926# 0.146647f
C123 a_48_n484# a_n746_n7926# 0.146647f
C124 a_n118_n2564# a_n746_n7926# 0.146647f
C125 a_n118_n484# a_n746_n7926# 0.146647f
C126 a_n284_n2564# a_n746_n7926# 0.146647f
C127 a_n284_n484# a_n746_n7926# 0.146647f
C128 a_n450_n2564# a_n746_n7926# 0.146647f
C129 a_n450_n484# a_n746_n7926# 0.146647f
C130 a_n616_n2564# a_n746_n7926# 0.356961f
C131 a_n616_n484# a_n746_n7926# 0.356961f
C132 a_546_52# a_n746_n7926# 0.356961f
C133 a_546_2132# a_n746_n7926# 0.356961f
C134 a_380_52# a_n746_n7926# 0.146647f
C135 a_380_2132# a_n746_n7926# 0.146647f
C136 a_214_52# a_n746_n7926# 0.146647f
C137 a_214_2132# a_n746_n7926# 0.146647f
C138 a_48_52# a_n746_n7926# 0.146647f
C139 a_48_2132# a_n746_n7926# 0.146647f
C140 a_n118_52# a_n746_n7926# 0.146647f
C141 a_n118_2132# a_n746_n7926# 0.146647f
C142 a_n284_52# a_n746_n7926# 0.146647f
C143 a_n284_2132# a_n746_n7926# 0.146647f
C144 a_n450_52# a_n746_n7926# 0.146647f
C145 a_n450_2132# a_n746_n7926# 0.146647f
C146 a_n616_52# a_n746_n7926# 0.356961f
C147 a_n616_2132# a_n746_n7926# 0.356961f
C148 a_546_2668# a_n746_n7926# 0.356961f
C149 a_546_4748# a_n746_n7926# 0.356961f
C150 a_380_2668# a_n746_n7926# 0.146647f
C151 a_380_4748# a_n746_n7926# 0.146647f
C152 a_214_2668# a_n746_n7926# 0.146647f
C153 a_214_4748# a_n746_n7926# 0.146647f
C154 a_48_2668# a_n746_n7926# 0.146647f
C155 a_48_4748# a_n746_n7926# 0.146647f
C156 a_n118_2668# a_n746_n7926# 0.146647f
C157 a_n118_4748# a_n746_n7926# 0.146647f
C158 a_n284_2668# a_n746_n7926# 0.146647f
C159 a_n284_4748# a_n746_n7926# 0.146647f
C160 a_n450_2668# a_n746_n7926# 0.146647f
C161 a_n450_4748# a_n746_n7926# 0.146647f
C162 a_n616_2668# a_n746_n7926# 0.356961f
C163 a_n616_4748# a_n746_n7926# 0.356961f
C164 a_546_5284# a_n746_n7926# 0.356961f
C165 a_546_7364# a_n746_n7926# 0.387223f
C166 a_380_5284# a_n746_n7926# 0.146647f
C167 a_380_7364# a_n746_n7926# 0.17691f
C168 a_214_5284# a_n746_n7926# 0.146647f
C169 a_214_7364# a_n746_n7926# 0.17691f
C170 a_48_5284# a_n746_n7926# 0.146647f
C171 a_48_7364# a_n746_n7926# 0.17691f
C172 a_n118_5284# a_n746_n7926# 0.146647f
C173 a_n118_7364# a_n746_n7926# 0.17691f
C174 a_n284_5284# a_n746_n7926# 0.146647f
C175 a_n284_7364# a_n746_n7926# 0.17691f
C176 a_n450_5284# a_n746_n7926# 0.146647f
C177 a_n450_7364# a_n746_n7926# 0.17691f
C178 a_n616_5284# a_n746_n7926# 0.356961f
C179 a_n616_7364# a_n746_n7926# 0.387223f
.ends

.subckt res_trim AVSS A B 3 2 1
Xsky130_fd_pr__res_high_po_0p35_KQ9YC9_0 B 3 B 3 3 3 3 3 B 3 B 2 B B B B 1 2 B 2 3
+ 2 3 B 3 3 AVSS 2 B 3 3 B 3 2 3 2 3 1 2 3 3 B B B B 1 3 3 3 3 B B 3 2 3 3 3 2 A A
+ B B 2 2 1 B 3 B 3 B 3 3 B B 3 3 B 3 1 3 1 B 3 B 2 B 2 B 3 B 3 3 B 3 3 3 3 sky130_fd_pr__res_high_po_0p35_KQ9YC9
C0 A 3 0.18657f
C1 A 1 0.918452f
C2 1 3 2.919634f
C3 A 2 1.948186f
C4 A B 0.209476f
C5 2 3 1.850388f
C6 B 3 1.388352f
C7 1 2 1.329232f
C8 B 1 0.298952f
C9 B 2 3.728792f
C10 1 AVSS 9.578271f
C11 3 AVSS 19.373535f
C12 2 AVSS 11.816302f
C13 B AVSS 11.956904f
C14 A AVSS 2.781555f
.ends

.subckt sky130_fd_pr__pfet_01v8_C2SJBD a_n2029_n128# w_n4181_n164# a_2029_n64# a_n4145_n64#
+ a_2087_n128# a_4087_n64# a_n4087_n128# a_29_n128# a_n2087_n64# a_n29_n64# VSUBS
X0 a_n2087_n64# a_n4087_n128# a_n4145_n64# w_n4181_n164# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=10
X1 a_2029_n64# a_29_n128# a_n29_n64# w_n4181_n164# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=10
X2 a_n29_n64# a_n2029_n128# a_n2087_n64# w_n4181_n164# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=10
X3 a_4087_n64# a_2087_n128# a_2029_n64# w_n4181_n164# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=10
C0 a_29_n128# w_n4181_n164# 0.821111f
C1 a_n2029_n128# w_n4181_n164# 0.821111f
C2 w_n4181_n164# a_n4087_n128# 0.823465f
C3 a_2087_n128# w_n4181_n164# 0.823465f
C4 a_4087_n64# VSUBS 0.149664f
C5 a_2029_n64# VSUBS 0.112935f
C6 a_n29_n64# VSUBS 0.112935f
C7 a_n2087_n64# VSUBS 0.112935f
C8 a_n4145_n64# VSUBS 0.149664f
C9 a_2087_n128# VSUBS 2.76013f
C10 a_29_n128# VSUBS 2.74139f
C11 a_n2029_n128# VSUBS 2.74139f
C12 a_n4087_n128# VSUBS 2.76013f
C13 w_n4181_n164# VSUBS 9.08113f
.ends

.subckt sky130_fd_pr__pfet_01v8_8WJJP2 a_n2029_n162# a_2087_n162# a_4087_n136# a_n2087_n136#
+ a_n4087_n162# a_29_n162# w_n4181_n198# a_2029_n136# a_n29_n136# a_n4145_n136# VSUBS
X0 a_4087_n136# a_2087_n162# a_2029_n136# w_n4181_n198# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=10
X1 a_n2087_n136# a_n4087_n162# a_n4145_n136# w_n4181_n198# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=10
X2 a_2029_n136# a_29_n162# a_n29_n136# w_n4181_n198# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=10
X3 a_n29_n136# a_n2029_n162# a_n2087_n136# w_n4181_n198# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=10
C0 a_n4087_n162# w_n4181_n198# 0.823465f
C1 a_29_n162# w_n4181_n198# 0.821111f
C2 w_n4181_n198# a_n2029_n162# 0.821111f
C3 a_2087_n162# w_n4181_n198# 0.823465f
C4 a_4087_n136# VSUBS 0.149664f
C5 a_2029_n136# VSUBS 0.112935f
C6 a_n29_n136# VSUBS 0.112935f
C7 a_n2087_n136# VSUBS 0.112935f
C8 a_n4145_n136# VSUBS 0.149664f
C9 a_2087_n162# VSUBS 2.76013f
C10 a_29_n162# VSUBS 2.74139f
C11 a_n2029_n162# VSUBS 2.74139f
C12 a_n4087_n162# VSUBS 2.76013f
C13 w_n4181_n198# VSUBS 9.08113f
.ends

.subckt sky130_fd_pr__pfet_01v8_HVJJBB a_n29_n100# a_2029_n100# a_n4145_n100# a_n2029_n164#
+ a_2087_n164# w_n4181_n200# a_4087_n100# a_n4087_n164# a_n2087_n100# a_29_n164# VSUBS
X0 a_n2087_n100# a_n4087_n164# a_n4145_n100# w_n4181_n200# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=10
X1 a_2029_n100# a_29_n164# a_n29_n100# w_n4181_n200# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=10
X2 a_n29_n100# a_n2029_n164# a_n2087_n100# w_n4181_n200# sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=10
X3 a_4087_n100# a_2087_n164# a_2029_n100# w_n4181_n200# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=10
C0 a_29_n164# w_n4181_n200# 1.08317f
C1 w_n4181_n200# a_n4087_n164# 1.08575f
C2 w_n4181_n200# a_n2029_n164# 1.08317f
C3 a_2087_n164# w_n4181_n200# 1.08575f
C4 a_4087_n100# VSUBS 0.148535f
C5 a_2029_n100# VSUBS 0.111805f
C6 a_n29_n100# VSUBS 0.111805f
C7 a_n2087_n100# VSUBS 0.111805f
C8 a_n4145_n100# VSUBS 0.148535f
C9 a_2087_n164# VSUBS 3.08243f
C10 a_29_n164# VSUBS 3.05214f
C11 a_n2029_n164# VSUBS 3.05214f
C12 a_n4087_n164# VSUBS 3.08243f
C13 w_n4181_n200# VSUBS 10.0344f
.ends

.subckt pmos_current_bgr D2 D1 vdde G10 D10
Xsky130_fd_pr__pfet_01v8_C2SJBD_0 vdde vdde vdde D10 G10 D10 G10 vdde vdde vdde VSUBS
+ sky130_fd_pr__pfet_01v8_C2SJBD
Xsky130_fd_pr__pfet_01v8_8WJJP2_1 vdde G10 D10 vdde G10 vdde vdde vdde vdde D10 VSUBS
+ sky130_fd_pr__pfet_01v8_8WJJP2
Xsky130_fd_pr__pfet_01v8_HVJJBB_0 D1 vdde D2 D10 D10 vdde D2 D10 vdde D10 VSUBS sky130_fd_pr__pfet_01v8_HVJJBB
Xsky130_fd_pr__pfet_01v8_HVJJBB_1 D1 vdde D2 D10 D10 vdde D2 D10 vdde D10 VSUBS sky130_fd_pr__pfet_01v8_HVJJBB
Xsky130_fd_pr__pfet_01v8_2XUZHN_0 D2 vdde D2 D2 VSUBS sky130_fd_pr__pfet_01v8_2XUZHN
Xsky130_fd_pr__pfet_01v8_2XUZHN_1 D10 vdde D10 D10 VSUBS sky130_fd_pr__pfet_01v8_2XUZHN
Xsky130_fd_pr__pfet_01v8_2XUZHN_2 D2 vdde D2 D2 VSUBS sky130_fd_pr__pfet_01v8_2XUZHN
Xsky130_fd_pr__pfet_01v8_2XUZHN_3 D2 vdde D2 D2 VSUBS sky130_fd_pr__pfet_01v8_2XUZHN
Xsky130_fd_pr__pfet_01v8_2XUZHN_4 D10 vdde D10 D10 VSUBS sky130_fd_pr__pfet_01v8_2XUZHN
Xsky130_fd_pr__pfet_01v8_2XUZHN_5 D10 vdde D10 D10 VSUBS sky130_fd_pr__pfet_01v8_2XUZHN
Xsky130_fd_pr__pfet_01v8_2XUZHN_6 D2 vdde D2 D2 VSUBS sky130_fd_pr__pfet_01v8_2XUZHN
Xsky130_fd_pr__pfet_01v8_2XUZHN_8 D10 vdde D10 D10 VSUBS sky130_fd_pr__pfet_01v8_2XUZHN
C0 vdde G10 10.459311f
C1 D10 vdde 12.84378f
C2 D10 D1 0.291251f
C3 G10 D2 0.993985f
C4 D10 D2 4.023208f
C5 vdde D2 1.296424f
C6 D10 G10 14.075364f
C7 D10 VSUBS 13.69858f
C8 vdde VSUBS 70.53953f
C9 D2 VSUBS 0.787072f
C10 D1 VSUBS 0.330152f
C11 G10 VSUBS 5.778857f
.ends

.subckt sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 Emitter Collector Base m=1
X0 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
C0 Emitter Base 0.896583f
C1 Base Collector 1.10722f
.ends

.subckt bjt B A sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|0]/Collector sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|1]/Collector
+ sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3|0]/Collector sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Collector
+ sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3|1]/Collector sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|3]/Collector
+ sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3|2]/Collector sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|4]/Collector
+ sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3|3]/Collector sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3|4]/Collector
+ VSUBS AVSS
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[0|0] AVSS AVSS AVSS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[1|0] AVSS AVSS AVSS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[2|0] AVSS AVSS AVSS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3|0] AVSS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3|0]/Collector
+ AVSS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|0] AVSS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|0]/Collector
+ AVSS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[0|1] AVSS AVSS AVSS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[1|1] B AVSS AVSS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[2|1] B AVSS AVSS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3|1] B sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3|1]/Collector
+ AVSS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|1] AVSS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|1]/Collector
+ AVSS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[0|2] AVSS AVSS AVSS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[1|2] B AVSS AVSS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[2|2] A AVSS AVSS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3|2] B sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3|2]/Collector
+ AVSS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2] AVSS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2]/Collector
+ AVSS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[0|3] AVSS AVSS AVSS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[1|3] B AVSS AVSS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[2|3] B AVSS AVSS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3|3] B sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3|3]/Collector
+ AVSS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|3] AVSS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|3]/Collector
+ AVSS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[0|4] AVSS AVSS AVSS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[1|4] AVSS AVSS AVSS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[2|4] AVSS AVSS AVSS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3|4] AVSS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3|4]/Collector
+ AVSS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|4] AVSS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|4]/Collector
+ AVSS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
C0 B A 0.569863f
C1 AVSS A 2.60218f
C2 AVSS B 6.489541f
C3 B VSUBS -0.55543f
C4 AVSS VSUBS 0.154621p
.ends

.subckt pmos_current_bgr_2 D3 D8 vdde D9 D4
Xsky130_fd_pr__pfet_01v8_CVRJBD_0 D9 D9 D9 D8 vdde vdde VSUBS sky130_fd_pr__pfet_01v8_CVRJBD
Xsky130_fd_pr__pfet_01v8_CVRJBD_1 D4 D3 D4 D4 vdde vdde VSUBS sky130_fd_pr__pfet_01v8_CVRJBD
Xsky130_fd_pr__pfet_01v8_8RMJP2_0 D4 D3 vdde D4 D4 vdde VSUBS sky130_fd_pr__pfet_01v8_8RMJP2
Xsky130_fd_pr__pfet_01v8_8RMJP2_1 D9 D9 vdde D9 D8 vdde VSUBS sky130_fd_pr__pfet_01v8_8RMJP2
Xsky130_fd_pr__pfet_01v8_2XUZHN_0 D9 vdde D9 D9 VSUBS sky130_fd_pr__pfet_01v8_2XUZHN
Xsky130_fd_pr__pfet_01v8_2XUZHN_1 D4 vdde D4 D4 VSUBS sky130_fd_pr__pfet_01v8_2XUZHN
Xsky130_fd_pr__pfet_01v8_2XUZHN_2 D8 vdde D8 D8 VSUBS sky130_fd_pr__pfet_01v8_2XUZHN
Xsky130_fd_pr__pfet_01v8_2XUZHN_3 D9 vdde D9 D9 VSUBS sky130_fd_pr__pfet_01v8_2XUZHN
Xsky130_fd_pr__pfet_01v8_2XUZHN_4 D3 vdde D3 D3 VSUBS sky130_fd_pr__pfet_01v8_2XUZHN
Xsky130_fd_pr__pfet_01v8_2XUZHN_5 D4 vdde D4 D4 VSUBS sky130_fd_pr__pfet_01v8_2XUZHN
Xsky130_fd_pr__pfet_01v8_2XUZHN_6 D8 vdde D8 D8 VSUBS sky130_fd_pr__pfet_01v8_2XUZHN
Xsky130_fd_pr__pfet_01v8_2XUZHN_7 D3 vdde D3 D3 VSUBS sky130_fd_pr__pfet_01v8_2XUZHN
C0 vdde D3 1.176749f
C1 D4 vdde 6.652088f
C2 D8 D3 0.583947f
C3 D4 D8 0.759468f
C4 vdde D8 0.664206f
C5 D9 D3 1.157008f
C6 D4 D9 3.206212f
C7 D9 vdde 2.934962f
C8 D9 D8 2.129757f
C9 D4 D3 1.031305f
C10 D4 VSUBS 6.223401f
C11 D3 VSUBS 1.574039f
C12 vdde VSUBS 34.590233f
C13 D8 VSUBS 0.871461f
C14 D9 VSUBS 5.173591f
.ends

.subckt sky130_fd_pr__res_high_po_0p35_RXTQM4 a_380_1352# a_380_n484# a_n284_n1784#
+ a_214_1352# a_214_n484# a_48_52# a_48_1352# a_48_n484# a_n118_n1784# a_380_n1784#
+ a_n450_52# a_n450_1352# a_380_52# a_n284_52# a_n450_n1784# a_n450_n484# a_214_52#
+ a_214_n1784# a_n118_52# a_n284_1352# a_n284_n484# a_n118_1352# a_48_n1784# a_n118_n484#
+ VSUBS
X0 a_n450_n484# a_n450_n1784# VSUBS sky130_fd_pr__res_high_po_0p35 l=4.5
X1 a_n284_n484# a_n284_n1784# VSUBS sky130_fd_pr__res_high_po_0p35 l=4.5
X2 a_n118_1352# a_n118_52# VSUBS sky130_fd_pr__res_high_po_0p35 l=4.5
X3 a_48_1352# a_48_52# VSUBS sky130_fd_pr__res_high_po_0p35 l=4.5
X4 a_48_n484# a_48_n1784# VSUBS sky130_fd_pr__res_high_po_0p35 l=4.5
X5 a_214_1352# a_214_52# VSUBS sky130_fd_pr__res_high_po_0p35 l=4.5
X6 a_n284_1352# a_n284_52# VSUBS sky130_fd_pr__res_high_po_0p35 l=4.5
X7 a_380_1352# a_380_52# VSUBS sky130_fd_pr__res_high_po_0p35 l=4.5
X8 a_214_n484# a_214_n1784# VSUBS sky130_fd_pr__res_high_po_0p35 l=4.5
X9 a_n118_n484# a_n118_n1784# VSUBS sky130_fd_pr__res_high_po_0p35 l=4.5
X10 a_n450_1352# a_n450_52# VSUBS sky130_fd_pr__res_high_po_0p35 l=4.5
X11 a_380_n484# a_380_n1784# VSUBS sky130_fd_pr__res_high_po_0p35 l=4.5
C0 a_214_n1784# a_380_n1784# 0.296258f
C1 a_380_n484# a_214_n484# 0.296258f
C2 a_n118_1352# a_n284_1352# 0.296258f
C3 a_n284_1352# a_n450_1352# 0.296258f
C4 a_214_52# a_380_52# 0.296258f
C5 a_n450_52# a_n284_52# 0.296258f
C6 a_n284_n484# a_n450_n484# 0.296258f
C7 a_48_n1784# a_n118_n1784# 0.296258f
C8 a_48_52# a_n118_52# 0.296258f
C9 a_n118_n1784# a_n284_n1784# 0.296258f
C10 a_48_n1784# a_214_n1784# 0.296258f
C11 a_214_1352# a_48_1352# 0.296258f
C12 a_214_1352# a_380_1352# 0.296258f
C13 a_n118_n484# a_48_n484# 0.296258f
C14 a_n284_n484# a_n118_n484# 0.296258f
C15 a_n284_52# a_n118_52# 0.296258f
C16 a_n118_1352# a_48_1352# 0.296258f
C17 a_214_n484# a_48_n484# 0.296258f
C18 a_48_52# a_214_52# 0.296258f
C19 a_n284_n1784# a_n450_n1784# 0.296258f
C20 a_380_n1784# VSUBS 0.379926f
C21 a_380_n484# VSUBS 0.349738f
C22 a_214_n1784# VSUBS 0.171397f
C23 a_214_n484# VSUBS 0.141209f
C24 a_48_n1784# VSUBS 0.171397f
C25 a_48_n484# VSUBS 0.141209f
C26 a_n118_n1784# VSUBS 0.171397f
C27 a_n118_n484# VSUBS 0.141209f
C28 a_n284_n1784# VSUBS 0.171397f
C29 a_n284_n484# VSUBS 0.141209f
C30 a_n450_n1784# VSUBS 0.379926f
C31 a_n450_n484# VSUBS 0.349738f
C32 a_380_52# VSUBS 0.349738f
C33 a_380_1352# VSUBS 0.379926f
C34 a_214_52# VSUBS 0.141209f
C35 a_214_1352# VSUBS 0.171397f
C36 a_48_52# VSUBS 0.141209f
C37 a_48_1352# VSUBS 0.171397f
C38 a_n118_52# VSUBS 0.141209f
C39 a_n118_1352# VSUBS 0.171397f
C40 a_n284_52# VSUBS 0.141209f
C41 a_n284_1352# VSUBS 0.171397f
C42 a_n450_52# VSUBS 0.349738f
C43 a_n450_1352# VSUBS 0.379926f
.ends

.subckt resistor_op_tt A C B D AVSS m1_565_4092# m1_n99_4131# m1_n100_4024#
Xsky130_fd_pr__res_high_po_0p35_RXTQM4_0 AVSS m1_565_4092# A D m1_n100_4024# m1_n100_4024#
+ B m1_n99_4131# C AVSS m1_n265_4096# AVSS m1_565_4092# m1_n99_4131# AVSS m1_n265_4096#
+ m1_n99_4131# A m1_n100_4024# D m1_n100_4024# B C m1_n99_4131# AVSS sky130_fd_pr__res_high_po_0p35_RXTQM4
C0 AVSS m1_565_4092# 0.513483f
C1 C A 0.102033f
C2 B D 0.107281f
C3 m1_n100_4024# m1_n99_4131# 0.283262f
C4 AVSS m1_n265_4096# 0.51143f
C5 AVSS 0 -0.492796f
C6 C 0 0.464486f
C7 A 0 0.672239f
C8 m1_565_4092# 0 0.333004f
C9 m1_n100_4024# 0 0.831448f
C10 B 0 0.46606f
C11 m1_n99_4131# 0 0.714853f
C12 D 0 0.673631f
C13 m1_n265_4096# 0 0.335073f
.ends

.subckt sky130_fd_pr__nfet_01v8_3YKU97 a_n2058_n69# a_n2000_n124# a_2000_n69# VSUBS
X0 a_2000_n69# a_n2000_n124# a_n2058_n69# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=20
C0 a_2000_n69# VSUBS 0.157722f
C1 a_n2058_n69# VSUBS 0.157722f
C2 a_n2000_n124# VSUBS 7.01308f
.ends

.subckt sky130_fd_pr__nfet_01v8_P5G96Q a_n2000_n126# a_2000_n100# a_n2058_n100# VSUBS
X0 a_2000_n100# a_n2000_n126# a_n2058_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=20
C0 a_2000_n100# VSUBS 0.157722f
C1 a_n2058_n100# VSUBS 0.157722f
C2 a_n2000_n126# VSUBS 5.002221f
.ends

.subckt sky130_fd_pr__nfet_01v8_3KF9AC a_n2000_n157# a_2000_n131# a_n2058_n131# VSUBS
X0 a_2000_n131# a_n2000_n157# a_n2058_n131# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=20
C0 a_2000_n131# VSUBS 0.157722f
C1 a_n2058_n131# VSUBS 0.157722f
C2 a_n2000_n157# VSUBS 7.01308f
.ends

.subckt sky130_fd_pr__nfet_01v8_BSRS8Q a_n2000_n126# a_2000_n100# a_n2058_n100# VSUBS
X0 a_2000_n100# a_n2000_n126# a_n2058_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=20
C0 a_2000_n100# VSUBS 0.157722f
C1 a_n2058_n100# VSUBS 0.157722f
C2 a_n2000_n126# VSUBS 5.002221f
.ends

.subckt nmos_tail_current D4 S2 AVSS D1 D2 D3
Xsky130_fd_pr__nfet_01v8_3YKU97_0 AVSS D2 D2 AVSS sky130_fd_pr__nfet_01v8_3YKU97
Xsky130_fd_pr__nfet_01v8_P5G96Q_1 D2 S2 D1 AVSS sky130_fd_pr__nfet_01v8_P5G96Q
Xsky130_fd_pr__nfet_01v8_P5G96Q_4 D2 D3 AVSS AVSS sky130_fd_pr__nfet_01v8_P5G96Q
Xsky130_fd_pr__nfet_01v8_P5G96Q_6 D2 D4 AVSS AVSS sky130_fd_pr__nfet_01v8_P5G96Q
Xsky130_fd_pr__nfet_01v8_P5G96Q_5 D2 AVSS D4 AVSS sky130_fd_pr__nfet_01v8_P5G96Q
Xsky130_fd_pr__nfet_01v8_P5G96Q_7 D2 AVSS D3 AVSS sky130_fd_pr__nfet_01v8_P5G96Q
Xsky130_fd_pr__nfet_01v8_6H9P4D_0 D3 D3 D3 AVSS sky130_fd_pr__nfet_01v8_6H9P4D
Xsky130_fd_pr__nfet_01v8_6H9P4D_1 D2 D2 D2 AVSS sky130_fd_pr__nfet_01v8_6H9P4D
Xsky130_fd_pr__nfet_01v8_6H9P4D_2 D4 D4 D4 AVSS sky130_fd_pr__nfet_01v8_6H9P4D
Xsky130_fd_pr__nfet_01v8_6H9P4D_3 D1 D1 D1 AVSS sky130_fd_pr__nfet_01v8_6H9P4D
Xsky130_fd_pr__nfet_01v8_6H9P4D_4 D2 D2 D2 AVSS sky130_fd_pr__nfet_01v8_6H9P4D
Xsky130_fd_pr__nfet_01v8_6H9P4D_6 D4 D4 D4 AVSS sky130_fd_pr__nfet_01v8_6H9P4D
Xsky130_fd_pr__nfet_01v8_6H9P4D_5 D3 D3 D3 AVSS sky130_fd_pr__nfet_01v8_6H9P4D
Xsky130_fd_pr__nfet_01v8_6H9P4D_7 D1 D1 D1 AVSS sky130_fd_pr__nfet_01v8_6H9P4D
Xsky130_fd_pr__nfet_01v8_3KF9AC_0 D2 AVSS D2 AVSS sky130_fd_pr__nfet_01v8_3KF9AC
Xsky130_fd_pr__nfet_01v8_BSRS8Q_0 D2 D1 S2 AVSS sky130_fd_pr__nfet_01v8_BSRS8Q
C0 D4 D2 2.847725f
C1 D1 D4 0.749969f
C2 D1 D2 3.588877f
C3 D1 S2 0.12486f
C4 S2 D2 0.565761f
C5 D4 D3 1.267795f
C6 D1 D3 2.494244f
C7 D3 D2 1.957817f
C8 D1 AVSS 3.524498f
C9 D4 AVSS 2.129397f
C10 D3 AVSS 1.150177f
C11 S2 AVSS 1.074352f
C12 D2 AVSS 46.281666f
.ends

.subckt sky130_fd_pr__nfet_01v8_2A7GYR a_15_n90# a_n73_n90# a_n15_n116# VSUBS
X0 a_15_n90# a_n15_n116# a_n73_n90# VSUBS sky130_fd_pr__nfet_01v8 ad=0.261 pd=2.38 as=0.261 ps=2.38 w=0.9 l=0.15
C0 a_15_n90# a_n73_n90# 0.14622f
C1 a_15_n90# VSUBS 0.109913f
C2 a_n73_n90# VSUBS 0.109913f
.ends

.subckt sky130_fd_pr__nfet_01v8_G26DVX a_n2687_n90# a_n29_n90# a_n2629_n145# a_29_n145#
+ a_2629_n90# VSUBS
X0 a_n29_n90# a_n2629_n145# a_n2687_n90# VSUBS sky130_fd_pr__nfet_01v8 ad=0.1305 pd=1.19 as=0.261 ps=2.38 w=0.9 l=13
X1 a_2629_n90# a_29_n145# a_n29_n90# VSUBS sky130_fd_pr__nfet_01v8 ad=0.261 pd=2.38 as=0.1305 ps=1.19 w=0.9 l=13
C0 a_2629_n90# VSUBS 0.144951f
C1 a_n29_n90# VSUBS 0.108693f
C2 a_n2687_n90# VSUBS 0.144951f
C3 a_29_n145# VSUBS 5.227221f
C4 a_n2629_n145# VSUBS 5.227221f
.ends

.subckt sky130_fd_pr__nfet_01v8_7RJ44K a_n29_n121# a_n2687_n121# a_29_n147# a_n2629_n147#
+ a_2629_n121# VSUBS
X0 a_n29_n121# a_n2629_n147# a_n2687_n121# VSUBS sky130_fd_pr__nfet_01v8 ad=0.1305 pd=1.19 as=0.261 ps=2.38 w=0.9 l=13
X1 a_2629_n121# a_29_n147# a_n29_n121# VSUBS sky130_fd_pr__nfet_01v8 ad=0.261 pd=2.38 as=0.1305 ps=1.19 w=0.9 l=13
C0 a_2629_n121# VSUBS 0.144951f
C1 a_n29_n121# VSUBS 0.108693f
C2 a_n2687_n121# VSUBS 0.144951f
C3 a_29_n147# VSUBS 4.57928f
C4 a_n2629_n147# VSUBS 4.57928f
.ends

.subckt differential_pair AVSS S D3 D4 PLUS MINUS
Xsky130_fd_pr__nfet_01v8_2A7GYR_0 D3 D3 D3 AVSS sky130_fd_pr__nfet_01v8_2A7GYR
Xsky130_fd_pr__nfet_01v8_2A7GYR_1 D4 D4 D4 AVSS sky130_fd_pr__nfet_01v8_2A7GYR
Xsky130_fd_pr__nfet_01v8_2A7GYR_2 D4 D4 D4 AVSS sky130_fd_pr__nfet_01v8_2A7GYR
Xsky130_fd_pr__nfet_01v8_2A7GYR_4 D3 D3 D3 AVSS sky130_fd_pr__nfet_01v8_2A7GYR
Xsky130_fd_pr__nfet_01v8_G26DVX_0 D4 S MINUS PLUS D3 AVSS sky130_fd_pr__nfet_01v8_G26DVX
Xsky130_fd_pr__nfet_01v8_7RJ44K_0 S D3 MINUS PLUS D4 AVSS sky130_fd_pr__nfet_01v8_7RJ44K
C0 PLUS D4 0.239957f
C1 MINUS S 1.733783f
C2 MINUS D3 0.625456f
C3 D4 S 0.541965f
C4 D3 D4 0.945324f
C5 PLUS S 1.490222f
C6 MINUS D4 0.458755f
C7 PLUS D3 1.422312f
C8 MINUS PLUS 2.886209f
C9 D3 S 0.614386f
C10 D3 AVSS 2.60901f
C11 PLUS AVSS 9.041692f
C12 S AVSS 8.293343f
C13 D4 AVSS 2.61774f
C14 MINUS AVSS 7.922267f
.ends

.subckt sky130_fd_pr__res_high_po_0p35_SU58NF a_n616_3852# a_712_8188# a_n782_n484#
+ a_48_n8620# a_n284_n12956# a_48_4388# a_712_n12956# a_n284_12524# a_n284_n9156#
+ a_214_3852# a_n118_8724# a_380_n484# a_712_4388# a_546_8188# a_n616_12524# a_48_n4820#
+ a_n782_n8620# a_n616_n9156# a_n616_n484# a_380_n4284# a_546_n8620# a_n782_8724#
+ a_546_4388# a_712_n4284# a_n782_n4820# a_48_n12956# a_214_n484# a_48_3852# a_380_8724#
+ a_546_n4820# a_n118_12524# a_712_52# a_n782_52# a_n284_n8620# a_n118_n9156# a_n450_8188#
+ a_48_52# a_712_3852# a_n616_52# a_n616_8724# a_n450_n4284# a_n616_n8620# a_546_52#
+ a_214_n4284# a_214_n12956# a_n284_n4820# a_n284_8188# a_n450_4388# a_48_n484# a_214_8724#
+ a_546_3852# a_n616_n4820# a_n616_n12956# a_712_n484# a_380_12524# a_380_n9156# a_n284_4388#
+ a_n118_n8620# a_712_12524# a_546_n12956# a_712_n9156# a_n118_8188# a_48_8724# a_48_n4284#
+ a_546_n484# a_n118_n4820# a_n450_3852# a_n782_8188# a_712_8724# a_n450_n12956# a_n118_4388#
+ a_n450_12524# a_n450_52# a_n450_n9156# a_n782_n4284# a_214_12524# a_380_n8620# a_214_n9156#
+ a_n284_3852# a_380_8188# a_546_n4284# a_380_n12956# a_380_52# a_n782_4388# a_546_8724#
+ a_n284_52# a_712_n8620# a_214_52# a_n450_n484# a_n118_n12956# a_n616_8188# a_n782_n12956#
+ a_n118_52# a_380_n4820# a_380_4388# a_n284_n4284# a_712_n4820# a_n118_3852# a_214_8188#
+ a_n284_n484# a_n616_4388# a_48_12524# a_n450_n8620# a_n616_n4284# a_48_n9156# a_214_n8620#
+ a_n450_8724# a_n782_3852# a_214_4388# a_n450_n4820# a_n782_12524# a_n782_n9156#
+ a_214_n4820# a_48_8188# a_n118_n484# a_380_3852# a_546_12524# a_n284_8724# a_546_n9156#
+ VSUBS a_n118_n4284#
X0 a_214_n4820# a_214_n8620# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X1 a_n284_n9156# a_n284_n12956# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X2 a_712_n484# a_712_n4284# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X3 a_n118_n484# a_n118_n4284# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X4 a_n616_n9156# a_n616_n12956# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X5 a_n616_8188# a_n616_4388# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X6 a_380_8188# a_380_4388# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X7 a_n118_3852# a_n118_52# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X8 a_48_3852# a_48_52# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X9 a_712_n4820# a_712_n8620# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X10 a_48_n9156# a_48_n12956# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X11 a_n118_n4820# a_n118_n8620# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X12 a_n616_12524# a_n616_8724# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X13 a_380_12524# a_380_8724# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X14 a_214_3852# a_214_52# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X15 a_n616_n484# a_n616_n4284# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X16 a_546_8188# a_546_4388# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X17 a_214_n9156# a_214_n12956# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X18 a_n616_3852# a_n616_52# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X19 a_380_n484# a_380_n4284# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X20 a_546_n484# a_546_n4284# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X21 a_n284_3852# a_n284_52# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X22 a_n616_n4820# a_n616_n8620# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X23 a_546_12524# a_546_8724# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X24 a_712_3852# a_712_52# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X25 a_380_n4820# a_380_n8620# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X26 a_546_n4820# a_546_n8620# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X27 a_n782_n9156# a_n782_n12956# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X28 a_214_8188# a_214_4388# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X29 a_380_3852# a_380_52# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X30 a_546_n9156# a_546_n12956# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X31 a_n284_8188# a_n284_4388# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X32 a_n782_3852# a_n782_52# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X33 a_n450_n484# a_n450_n4284# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X34 a_n284_n484# a_n284_n4284# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X35 a_214_12524# a_214_8724# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X36 a_48_n484# a_48_n4284# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X37 a_n284_12524# a_n284_8724# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X38 a_n450_n4820# a_n450_n8620# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X39 a_n284_n4820# a_n284_n8620# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X40 a_380_n9156# a_380_n12956# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X41 a_48_n4820# a_48_n8620# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X42 a_48_8188# a_48_4388# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X43 a_n782_n484# a_n782_n4284# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X44 a_712_n9156# a_712_n12956# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X45 a_n450_8188# a_n450_4388# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X46 a_712_8188# a_712_4388# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X47 a_n118_n9156# a_n118_n12956# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X48 a_48_12524# a_48_8724# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X49 a_n782_n4820# a_n782_n8620# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X50 a_n450_12524# a_n450_8724# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X51 a_n782_8188# a_n782_4388# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X52 a_n118_8188# a_n118_4388# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X53 a_712_12524# a_712_8724# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X54 a_n450_3852# a_n450_52# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X55 a_n782_12524# a_n782_8724# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X56 a_n118_12524# a_n118_8724# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X57 a_214_n484# a_214_n4284# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X58 a_n450_n9156# a_n450_n12956# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
X59 a_546_3852# a_546_52# VSUBS sky130_fd_pr__res_high_po_0p35 l=17
C0 a_n450_n12956# a_n616_n12956# 0.296258f
C1 a_n284_n12956# a_n118_n12956# 0.296258f
C2 a_n616_n484# a_n450_n484# 0.296258f
C3 a_380_n12956# a_546_n12956# 0.296258f
C4 a_n118_n8620# a_48_n8620# 0.296258f
C5 a_48_12524# a_n118_12524# 0.296258f
C6 a_n284_n12956# a_n450_n12956# 0.296258f
C7 a_48_52# a_n118_52# 0.296258f
C8 a_n284_n484# a_n450_n484# 0.296258f
C9 a_n450_n9156# a_n616_n9156# 0.296258f
C10 a_712_n9156# a_546_n9156# 0.296258f
C11 a_214_n4284# a_48_n4284# 0.296258f
C12 a_n616_4388# a_n782_4388# 0.296258f
C13 a_380_8724# a_546_8724# 0.296258f
C14 a_n616_3852# a_n450_3852# 0.296258f
C15 a_n782_8724# a_n616_8724# 0.296258f
C16 a_n450_n4284# a_n616_n4284# 0.296258f
C17 a_n616_4388# a_n450_4388# 0.296258f
C18 a_n782_n9156# a_n616_n9156# 0.296258f
C19 a_214_n12956# a_48_n12956# 0.296258f
C20 a_380_n9156# a_214_n9156# 0.296258f
C21 a_380_n4820# a_214_n4820# 0.296258f
C22 a_48_8188# a_n118_8188# 0.296258f
C23 a_712_52# a_546_52# 0.296258f
C24 a_n616_n8620# a_n450_n8620# 0.296258f
C25 a_n284_n4820# a_n450_n4820# 0.296258f
C26 a_546_4388# a_712_4388# 0.296258f
C27 a_214_52# a_48_52# 0.296258f
C28 a_546_12524# a_712_12524# 0.296258f
C29 a_712_n12956# a_546_n12956# 0.296258f
C30 a_n450_n9156# a_n284_n9156# 0.296258f
C31 a_n616_n8620# a_n782_n8620# 0.296258f
C32 a_546_8188# a_712_8188# 0.296258f
C33 a_n782_n4284# a_n616_n4284# 0.296258f
C34 a_380_52# a_546_52# 0.296258f
C35 a_214_52# a_380_52# 0.296258f
C36 a_n118_3852# a_n284_3852# 0.296258f
C37 a_n118_n4284# a_48_n4284# 0.296258f
C38 a_546_8188# a_380_8188# 0.296258f
C39 a_214_8724# a_48_8724# 0.296258f
C40 a_n782_n484# a_n616_n484# 0.296258f
C41 a_n616_12524# a_n450_12524# 0.296258f
C42 a_380_n8620# a_214_n8620# 0.296258f
C43 a_n450_n4284# a_n284_n4284# 0.296258f
C44 a_n450_8188# a_n284_8188# 0.296258f
C45 a_214_12524# a_380_12524# 0.296258f
C46 a_712_3852# a_546_3852# 0.296258f
C47 a_n616_8188# a_n782_8188# 0.296258f
C48 a_n616_n4820# a_n450_n4820# 0.296258f
C49 a_n284_8724# a_n118_8724# 0.296258f
C50 a_n284_8724# a_n450_8724# 0.296258f
C51 a_214_8188# a_48_8188# 0.296258f
C52 a_48_n4820# a_214_n4820# 0.296258f
C53 a_n118_n4284# a_n284_n4284# 0.296258f
C54 a_n284_52# a_n118_52# 0.296258f
C55 a_380_n484# a_214_n484# 0.296258f
C56 a_712_n484# a_546_n484# 0.296258f
C57 a_n616_52# a_n450_52# 0.296258f
C58 a_n284_4388# a_n118_4388# 0.296258f
C59 a_546_n484# a_380_n484# 0.296258f
C60 a_48_n484# a_n118_n484# 0.296258f
C61 a_n118_n484# a_n284_n484# 0.296258f
C62 a_n118_3852# a_48_3852# 0.296258f
C63 a_380_4388# a_546_4388# 0.296258f
C64 a_546_8724# a_712_8724# 0.296258f
C65 a_380_n4284# a_214_n4284# 0.296258f
C66 a_n118_n9156# a_n284_n9156# 0.296258f
C67 a_n782_3852# a_n616_3852# 0.296258f
C68 a_n616_n12956# a_n782_n12956# 0.296258f
C69 a_380_n4284# a_546_n4284# 0.296258f
C70 a_214_n9156# a_48_n9156# 0.296258f
C71 a_n284_4388# a_n450_4388# 0.296258f
C72 a_n616_8724# a_n450_8724# 0.296258f
C73 a_712_n8620# a_546_n8620# 0.296258f
C74 a_48_n4820# a_n118_n4820# 0.296258f
C75 a_n284_n8620# a_n118_n8620# 0.296258f
C76 a_n284_12524# a_n450_12524# 0.296258f
C77 a_48_n484# a_214_n484# 0.296258f
C78 a_380_n8620# a_546_n8620# 0.296258f
C79 a_546_12524# a_380_12524# 0.296258f
C80 a_n118_8724# a_48_8724# 0.296258f
C81 a_n284_3852# a_n450_3852# 0.296258f
C82 a_214_8188# a_380_8188# 0.296258f
C83 a_n616_8188# a_n450_8188# 0.296258f
C84 a_380_n4820# a_546_n4820# 0.296258f
C85 a_214_3852# a_48_3852# 0.296258f
C86 a_546_n4284# a_712_n4284# 0.296258f
C87 a_380_n9156# a_546_n9156# 0.296258f
C88 a_214_3852# a_380_3852# 0.296258f
C89 a_n118_n12956# a_48_n12956# 0.296258f
C90 a_n616_12524# a_n782_12524# 0.296258f
C91 a_712_n4820# a_546_n4820# 0.296258f
C92 a_n616_52# a_n782_52# 0.296258f
C93 a_214_n8620# a_48_n8620# 0.296258f
C94 a_n284_n8620# a_n450_n8620# 0.296258f
C95 a_n284_8188# a_n118_8188# 0.296258f
C96 a_546_3852# a_380_3852# 0.296258f
C97 a_n782_n4820# a_n616_n4820# 0.296258f
C98 a_n284_12524# a_n118_12524# 0.296258f
C99 a_n284_52# a_n450_52# 0.296258f
C100 a_380_4388# a_214_4388# 0.296258f
C101 a_48_4388# a_214_4388# 0.296258f
C102 a_n284_n4820# a_n118_n4820# 0.296258f
C103 a_380_8724# a_214_8724# 0.296258f
C104 a_214_n12956# a_380_n12956# 0.296258f
C105 a_48_4388# a_n118_4388# 0.296258f
C106 a_n118_n9156# a_48_n9156# 0.296258f
C107 a_48_12524# a_214_12524# 0.296258f
C108 a_712_n12956# VSUBS 0.385365f
C109 a_712_n9156# VSUBS 0.355177f
C110 a_546_n12956# VSUBS 0.176835f
C111 a_546_n9156# VSUBS 0.146647f
C112 a_380_n12956# VSUBS 0.176835f
C113 a_380_n9156# VSUBS 0.146647f
C114 a_214_n12956# VSUBS 0.176835f
C115 a_214_n9156# VSUBS 0.146647f
C116 a_48_n12956# VSUBS 0.176835f
C117 a_48_n9156# VSUBS 0.146647f
C118 a_n118_n12956# VSUBS 0.176835f
C119 a_n118_n9156# VSUBS 0.146647f
C120 a_n284_n12956# VSUBS 0.176835f
C121 a_n284_n9156# VSUBS 0.146647f
C122 a_n450_n12956# VSUBS 0.176835f
C123 a_n450_n9156# VSUBS 0.146647f
C124 a_n616_n12956# VSUBS 0.176835f
C125 a_n616_n9156# VSUBS 0.146647f
C126 a_n782_n12956# VSUBS 0.385365f
C127 a_n782_n9156# VSUBS 0.355177f
C128 a_712_n8620# VSUBS 0.355177f
C129 a_712_n4820# VSUBS 0.355177f
C130 a_546_n8620# VSUBS 0.146647f
C131 a_546_n4820# VSUBS 0.146647f
C132 a_380_n8620# VSUBS 0.146647f
C133 a_380_n4820# VSUBS 0.146647f
C134 a_214_n8620# VSUBS 0.146647f
C135 a_214_n4820# VSUBS 0.146647f
C136 a_48_n8620# VSUBS 0.146647f
C137 a_48_n4820# VSUBS 0.146647f
C138 a_n118_n8620# VSUBS 0.146647f
C139 a_n118_n4820# VSUBS 0.146647f
C140 a_n284_n8620# VSUBS 0.146647f
C141 a_n284_n4820# VSUBS 0.146647f
C142 a_n450_n8620# VSUBS 0.146647f
C143 a_n450_n4820# VSUBS 0.146647f
C144 a_n616_n8620# VSUBS 0.146647f
C145 a_n616_n4820# VSUBS 0.146647f
C146 a_n782_n8620# VSUBS 0.355177f
C147 a_n782_n4820# VSUBS 0.355177f
C148 a_712_n4284# VSUBS 0.355177f
C149 a_712_n484# VSUBS 0.355177f
C150 a_546_n4284# VSUBS 0.146647f
C151 a_546_n484# VSUBS 0.146647f
C152 a_380_n4284# VSUBS 0.146647f
C153 a_380_n484# VSUBS 0.146647f
C154 a_214_n4284# VSUBS 0.146647f
C155 a_214_n484# VSUBS 0.146647f
C156 a_48_n4284# VSUBS 0.146647f
C157 a_48_n484# VSUBS 0.146647f
C158 a_n118_n4284# VSUBS 0.146647f
C159 a_n118_n484# VSUBS 0.146647f
C160 a_n284_n4284# VSUBS 0.146647f
C161 a_n284_n484# VSUBS 0.146647f
C162 a_n450_n4284# VSUBS 0.146647f
C163 a_n450_n484# VSUBS 0.146647f
C164 a_n616_n4284# VSUBS 0.146647f
C165 a_n616_n484# VSUBS 0.146647f
C166 a_n782_n4284# VSUBS 0.355177f
C167 a_n782_n484# VSUBS 0.355177f
C168 a_712_52# VSUBS 0.355177f
C169 a_712_3852# VSUBS 0.355177f
C170 a_546_52# VSUBS 0.146647f
C171 a_546_3852# VSUBS 0.146647f
C172 a_380_52# VSUBS 0.146647f
C173 a_380_3852# VSUBS 0.146647f
C174 a_214_52# VSUBS 0.146647f
C175 a_214_3852# VSUBS 0.146647f
C176 a_48_52# VSUBS 0.146647f
C177 a_48_3852# VSUBS 0.146647f
C178 a_n118_52# VSUBS 0.146647f
C179 a_n118_3852# VSUBS 0.146647f
C180 a_n284_52# VSUBS 0.146647f
C181 a_n284_3852# VSUBS 0.146647f
C182 a_n450_52# VSUBS 0.146647f
C183 a_n450_3852# VSUBS 0.146647f
C184 a_n616_52# VSUBS 0.146647f
C185 a_n616_3852# VSUBS 0.146647f
C186 a_n782_52# VSUBS 0.355177f
C187 a_n782_3852# VSUBS 0.355177f
C188 a_712_4388# VSUBS 0.355177f
C189 a_712_8188# VSUBS 0.355177f
C190 a_546_4388# VSUBS 0.146647f
C191 a_546_8188# VSUBS 0.146647f
C192 a_380_4388# VSUBS 0.146647f
C193 a_380_8188# VSUBS 0.146647f
C194 a_214_4388# VSUBS 0.146647f
C195 a_214_8188# VSUBS 0.146647f
C196 a_48_4388# VSUBS 0.146647f
C197 a_48_8188# VSUBS 0.146647f
C198 a_n118_4388# VSUBS 0.146647f
C199 a_n118_8188# VSUBS 0.146647f
C200 a_n284_4388# VSUBS 0.146647f
C201 a_n284_8188# VSUBS 0.146647f
C202 a_n450_4388# VSUBS 0.146647f
C203 a_n450_8188# VSUBS 0.146647f
C204 a_n616_4388# VSUBS 0.146647f
C205 a_n616_8188# VSUBS 0.146647f
C206 a_n782_4388# VSUBS 0.355177f
C207 a_n782_8188# VSUBS 0.355177f
C208 a_712_8724# VSUBS 0.355177f
C209 a_712_12524# VSUBS 0.385365f
C210 a_546_8724# VSUBS 0.146647f
C211 a_546_12524# VSUBS 0.176835f
C212 a_380_8724# VSUBS 0.146647f
C213 a_380_12524# VSUBS 0.176835f
C214 a_214_8724# VSUBS 0.146647f
C215 a_214_12524# VSUBS 0.176835f
C216 a_48_8724# VSUBS 0.146647f
C217 a_48_12524# VSUBS 0.176835f
C218 a_n118_8724# VSUBS 0.146647f
C219 a_n118_12524# VSUBS 0.176835f
C220 a_n284_8724# VSUBS 0.146647f
C221 a_n284_12524# VSUBS 0.176835f
C222 a_n450_8724# VSUBS 0.146647f
C223 a_n450_12524# VSUBS 0.176835f
C224 a_n616_8724# VSUBS 0.146647f
C225 a_n616_12524# VSUBS 0.176835f
C226 a_n782_8724# VSUBS 0.355177f
C227 a_n782_12524# VSUBS 0.385365f
.ends

.subckt resist_const A C E VBGTC D B AVSS F m1_28308_n3465# m1_6628_n3631# m1_19584_n3310#
+ m1_19584_n3642# m1_10964_n3465# m1_15300_n3631# m1_10964_n3133# m1_6628_n2469# m1_15248_n3476#
+ m1_10912_n3310# m1_10912_n3642# m1_6576_n3476# m1_10964_n2635# m1_15300_n3299# VBGSC
+ m1_6628_n3299# m1_10912_n2812# m1_15300_n2469# m1_28256_n3642#
Xsky130_fd_pr__res_high_po_0p35_SU58NF_0 m1_10964_n3465# m1_6628_n2303# m1_15300_n3797#
+ m1_23920_n2978# m1_28256_n3642# m1_10964_n2967# AVSS m1_2337_n3299# m1_23920_n3144#
+ m1_10964_n2967# m1_6576_n3144# m1_15300_n2469# m1_10964_n2303# m1_6576_n2646# B
+ m1_19584_n2812# m1_23972_n3797# m1_23920_n3476# m1_15248_n3476# m1_19636_n2635#
+ m1_23972_n2469# m1_6628_n3797# m1_10912_n2480# m1_19636_n2303# m1_19636_n3797# m1_28308_n2967#
+ m1_10912_n2812# m1_10912_n2812# m1_6576_n2646# m1_19636_n2635# m1_2420_n3133# m1_15300_n2303#
+ m1_15300_n3797# m1_23972_n3299# m1_23972_n3299# m1_6628_n3631# m1_10912_n2812# m1_10964_n2303#
+ m1_15300_n3631# m1_6628_n3631# m1_19636_n3465# m1_23972_n3631# m1_15300_n2469# m1_19584_n2812#
+ m1_28256_n2812# m1_15300_n3299# m1_6576_n3144# m1_10964_n3465# m1_15265_n3133# m1_6628_n2801#
+ m1_10964_n2635# m1_19636_n3465# m1_28256_n3642# m1_15300_n2303# C m1_23972_n2469#
+ m1_10912_n3310# m1_23920_n3144# AVSS m1_28256_n2812# m1_23972_n2303# m1_6628_n3299#
+ m1_6576_n2978# F m1_15248_n2646# m1_19584_n3310# m1_10912_n3642# m1_6628_n3797#
+ m1_6628_n2303# m1_28308_n3465# m1_10964_n3133# D m1_15248_n3476# m1_23972_n3631#
+ m1_19636_n3797# m1_2337_n3299# m1_23920_n2646# m1_23920_n2978# m1_10964_n3133# m1_6628_n2469#
+ m1_19584_n2480# m1_28308_n2967# m1_15248_n2646# m1_10964_n3797# m1_6628_n2469# m1_15300_n3299#
+ m1_23972_n2303# VBGSC m1_15300_n3631# m1_28308_n3465# m1_6576_n3476# AVSS m1_15265_n3133#
+ m1_19584_n2480# m1_10964_n2635# m1_19584_n3310# m1_19636_n2303# E m1_6576_n2978#
+ m1_10912_n3310# m1_10912_n3642# m1_2420_n3133# m1_23920_n3476# m1_19584_n3642# VBGTC
+ VBGTC m1_6576_n3476# m1_10964_n3797# m1_10912_n2812# m1_19584_n3642# AVSS m1_23972_n3797#
+ VBGSC m1_6628_n2801# m1_15300_n3299# m1_10912_n2480# A m1_6628_n3299# m1_23920_n2646#
+ AVSS m1_15300_n3299# sky130_fd_pr__res_high_po_0p35_SU58NF
C0 m1_6628_n2801# m1_6576_n2978# 0.123612f
C1 m1_10912_n2812# m1_10912_n3310# 0.682569f
C2 m1_23972_n3631# m1_23920_n3476# 0.123612f
C3 m1_19584_n2480# m1_19636_n2635# 0.123612f
C4 m1_23972_n3299# m1_23920_n3144# 0.123612f
C5 m1_10964_n2635# m1_10912_n2480# 0.123612f
C6 m1_2337_n3299# m1_2420_n3133# 0.12066f
C7 F VBGSC 0.217142f
C8 m1_15300_n3797# AVSS 0.463496f
C9 AVSS m1_6628_n3797# 0.463496f
C10 m1_10912_n3310# E 0.10571f
C11 m1_15300_n3631# m1_15248_n3476# 0.123612f
C12 AVSS m1_6628_n2303# 0.515465f
C13 VBGTC m1_23920_n2978# 0.123612f
C14 m1_10964_n3797# AVSS 0.463496f
C15 m1_23972_n3797# AVSS 0.463496f
C16 m1_6576_n3144# m1_6628_n3299# 0.123612f
C17 m1_28308_n2967# m1_28256_n2812# 0.128644f
C18 m1_23972_n2303# AVSS 0.515465f
C19 m1_28256_n3642# m1_28308_n3465# 0.128644f
C20 m1_15300_n3299# VBGSC 0.463805f
C21 m1_19636_n3797# AVSS 0.463496f
C22 m1_19584_n3642# m1_19636_n3465# 0.123612f
C23 m1_6628_n3631# m1_6576_n3476# 0.123612f
C24 m1_23920_n2646# m1_23972_n2469# 0.123612f
C25 VBGSC m1_15265_n3133# 0.243373f
C26 m1_10912_n2812# VBGSC 0.394952f
C27 m1_19584_n2812# VBGSC 0.310029f
C28 m1_19636_n2303# AVSS 0.515465f
C29 m1_10912_n2812# m1_10964_n2967# 0.210157f
C30 m1_10912_n3642# m1_10964_n3465# 0.123612f
C31 AVSS m1_15300_n2303# 0.515465f
C32 m1_10912_n3310# m1_10964_n3133# 0.163826f
C33 m1_10964_n2303# AVSS 0.515466f
C34 m1_15300_n3299# m1_10912_n3310# 0.284662f
C35 m1_15300_n2469# m1_15248_n2646# 0.123612f
C36 m1_6576_n2646# m1_6628_n2469# 0.123612f
C37 m1_15300_n3299# m1_19584_n3310# 0.245791f
C38 m1_28256_n2812# 0 0.542836f
C39 m1_23920_n2646# 0 0.412976f
C40 m1_28308_n2967# 0 0.589905f
C41 m1_23920_n2978# 0 0.364019f
C42 m1_23972_n3299# 0 0.351297f
C43 m1_28308_n3465# 0 0.589905f
C44 m1_23972_n3631# 0 0.350405f
C45 m1_28256_n3642# 0 0.541353f
C46 m1_23972_n2303# 0 0.341828f
C47 m1_23972_n2469# 0 0.350405f
C48 m1_19636_n2635# 0 0.349811f
C49 VBGTC 0 0.351297f
C50 m1_23920_n3144# 0 0.364018f
C51 m1_23920_n3476# 0 0.4124f
C52 m1_23972_n3797# 0 0.353369f
C53 m1_19636_n2303# 0 0.341828f
C54 m1_19584_n2480# 0 0.412973f
C55 m1_15248_n2646# 0 0.411441f
C56 m1_19584_n2812# 0 0.353548f
C57 F 0 0.137592f
C58 m1_15265_n3133# 0 0.336237f
C59 m1_19584_n3310# 0 0.347065f
C60 m1_19636_n3465# 0 0.349811f
C61 m1_19584_n3642# 0 0.412397f
C62 m1_19636_n3797# 0 0.353369f
C63 m1_15300_n2303# 0 0.341828f
C64 m1_15300_n2469# 0 0.349811f
C65 VBGSC 0 1.465823f
C66 m1_10964_n2967# 0 0.351297f
C67 E 0 0.152796f
C68 m1_15300_n3299# 0 1.783432f
C69 m1_15248_n3476# 0 0.410865f
C70 m1_15300_n3631# 0 0.349811f
C71 m1_15300_n3797# 0 0.353369f
C72 m1_10964_n2303# 0 0.341828f
C73 m1_10912_n2480# 0 0.411444f
C74 m1_10964_n2635# 0 0.350405f
C75 m1_10912_n2812# 0 1.711577f
C76 m1_10964_n3133# 0 0.351297f
C77 m1_10912_n3310# 0 1.398506f
C78 m1_10964_n3465# 0 0.350405f
C79 m1_10912_n3642# 0 0.410868f
C80 m1_10964_n3797# 0 0.353369f
C81 m1_6628_n2303# 0 0.341828f
C82 AVSS 0 -35.174644f
C83 m1_6628_n2469# 0 0.350405f
C84 A 0 0.167761f
C85 m1_6576_n2646# 0 0.412976f
C86 C 0 0.159785f
C87 m1_6628_n2801# 0 0.351297f
C88 m1_2337_n3299# 0 0.708589f
C89 m1_6576_n2978# 0 0.364019f
C90 m1_2420_n3133# 0 0.31019f
C91 m1_6576_n3144# 0 0.364018f
C92 m1_6628_n3299# 0 0.351297f
C93 m1_6576_n3476# 0 0.4124f
C94 D 0 0.16058f
C95 m1_6628_n3631# 0 0.350405f
C96 B 0 0.166411f
C97 m1_6628_n3797# 0 0.353369f
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_SXWHWZ c1_n3852_3880# c1_4172_n7280# c1_n7864_3880#
+ c1_n7864_n3560# m3_4132_n3600# m3_n3892_3840# m3_120_n3600# c1_n3852_n3560# c1_160_160#
+ m3_n7904_3840# c1_n3852_160# m3_n3892_n7320# c1_160_n3560# c1_n7864_n7280# m3_4132_n7320#
+ m3_120_n7320# c1_4172_160# m3_4132_3840# c1_n3852_n7280# m3_n7904_n3600# c1_4172_3880#
+ m3_4132_120# m3_n3892_120# m3_120_3840# c1_160_n7280# c1_160_3880# c1_4172_n3560#
+ m3_n7904_120# m3_n7904_n7320# m3_n3892_n3600# c1_n7864_160# m3_120_120# VSUBS
X0 c1_4172_160# m3_4132_120# sky130_fd_pr__cap_mim_m3_1 l=17 w=17
X1 c1_160_3880# m3_120_3840# sky130_fd_pr__cap_mim_m3_1 l=17 w=17
X2 c1_4172_3880# m3_4132_3840# sky130_fd_pr__cap_mim_m3_1 l=17 w=17
X3 c1_n7864_160# m3_n7904_120# sky130_fd_pr__cap_mim_m3_1 l=17 w=17
X4 c1_160_n7280# m3_120_n7320# sky130_fd_pr__cap_mim_m3_1 l=17 w=17
X5 c1_4172_n7280# m3_4132_n7320# sky130_fd_pr__cap_mim_m3_1 l=17 w=17
X6 c1_n3852_160# m3_n3892_120# sky130_fd_pr__cap_mim_m3_1 l=17 w=17
X7 c1_n3852_n3560# m3_n3892_n3600# sky130_fd_pr__cap_mim_m3_1 l=17 w=17
X8 c1_n3852_3880# m3_n3892_3840# sky130_fd_pr__cap_mim_m3_1 l=17 w=17
X9 c1_n7864_3880# m3_n7904_3840# sky130_fd_pr__cap_mim_m3_1 l=17 w=17
X10 c1_160_160# m3_120_120# sky130_fd_pr__cap_mim_m3_1 l=17 w=17
X11 c1_n3852_n7280# m3_n3892_n7320# sky130_fd_pr__cap_mim_m3_1 l=17 w=17
X12 c1_n7864_n3560# m3_n7904_n3600# sky130_fd_pr__cap_mim_m3_1 l=17 w=17
X13 c1_n7864_n7280# m3_n7904_n7320# sky130_fd_pr__cap_mim_m3_1 l=17 w=17
X14 c1_160_n3560# m3_120_n3600# sky130_fd_pr__cap_mim_m3_1 l=17 w=17
X15 c1_4172_n3560# m3_4132_n3600# sky130_fd_pr__cap_mim_m3_1 l=17 w=17
C0 c1_160_3880# m3_n3892_3840# 0.717601f
C1 m3_4132_n3600# c1_4172_n3560# 26.168001f
C2 m3_120_120# m3_120_3840# 0.896911f
C3 m3_n3892_n7320# m3_120_n7320# 0.891312f
C4 c1_4172_n7280# c1_4172_n3560# 0.609898f
C5 m3_120_3840# m3_n3892_3840# 0.891312f
C6 c1_160_3880# m3_120_3840# 26.168001f
C7 m3_n7904_n3600# m3_n7904_n7320# 0.896911f
C8 c1_n7864_3880# c1_n7864_160# 0.609898f
C9 c1_160_n3560# c1_160_160# 0.609898f
C10 m3_n3892_n3600# m3_n7904_n3600# 0.891312f
C11 c1_160_160# m3_n3892_120# 0.717601f
C12 m3_120_n7320# m3_4132_n7320# 0.891312f
C13 c1_n3852_3880# m3_n7904_3840# 0.717601f
C14 m3_120_n3600# m3_120_n7320# 0.896911f
C15 m3_n7904_120# c1_n3852_160# 0.717601f
C16 c1_4172_n3560# c1_4172_160# 0.609898f
C17 m3_120_n3600# c1_4172_n3560# 0.717601f
C18 m3_n7904_120# m3_n7904_n3600# 0.896911f
C19 c1_n3852_3880# m3_n3892_3840# 26.168001f
C20 m3_n7904_120# c1_n7864_160# 26.168001f
C21 c1_160_n7280# m3_120_n7320# 26.168001f
C22 m3_n3892_n3600# c1_160_n3560# 0.717601f
C23 m3_n3892_n3600# m3_n3892_120# 0.896911f
C24 c1_n3852_n3560# c1_n3852_n7280# 0.609898f
C25 m3_n3892_n3600# c1_n3852_n3560# 26.168001f
C26 c1_4172_3880# m3_4132_3840# 26.168001f
C27 m3_120_120# m3_n3892_120# 0.891312f
C28 m3_120_120# c1_160_160# 26.168001f
C29 m3_n3892_3840# m3_n3892_120# 0.896911f
C30 m3_120_n3600# c1_160_n3560# 26.168001f
C31 c1_n3852_3880# c1_n3852_160# 0.609898f
C32 m3_n7904_120# m3_n3892_120# 0.891312f
C33 c1_160_3880# c1_160_160# 0.609898f
C34 m3_n3892_n7320# m3_n7904_n7320# 0.891312f
C35 c1_n7864_3880# m3_n7904_3840# 26.168001f
C36 m3_4132_n3600# m3_4132_n7320# 0.896911f
C37 m3_n3892_n7320# c1_n3852_n7280# 26.168001f
C38 m3_n7904_n7320# c1_n3852_n7280# 0.717601f
C39 m3_n3892_n3600# m3_n3892_n7320# 0.896911f
C40 c1_4172_n7280# m3_4132_n7320# 26.168001f
C41 m3_4132_n3600# m3_120_n3600# 0.891312f
C42 m3_4132_120# m3_4132_3840# 0.896911f
C43 c1_160_n3560# c1_160_n7280# 0.609898f
C44 m3_4132_n3600# m3_4132_120# 0.896911f
C45 m3_120_3840# m3_4132_3840# 0.891312f
C46 c1_4172_3880# c1_4172_160# 0.609898f
C47 c1_n7864_n3560# c1_n7864_n7280# 0.609898f
C48 c1_n3852_160# m3_n3892_120# 26.168001f
C49 m3_n7904_3840# m3_n3892_3840# 0.891312f
C50 c1_n3852_160# c1_n3852_n3560# 0.609898f
C51 m3_n7904_120# m3_n7904_3840# 0.896911f
C52 m3_n3892_n3600# m3_120_n3600# 0.891312f
C53 c1_4172_3880# m3_120_3840# 0.717601f
C54 m3_120_120# c1_4172_160# 0.717601f
C55 c1_4172_n7280# m3_120_n7320# 0.717601f
C56 m3_n7904_n7320# c1_n7864_n7280# 26.168001f
C57 m3_n7904_n3600# c1_n3852_n3560# 0.717601f
C58 c1_160_n7280# m3_n3892_n7320# 0.717601f
C59 m3_4132_120# c1_4172_160# 26.168001f
C60 m3_120_120# m3_120_n3600# 0.896911f
C61 m3_n7904_n3600# c1_n7864_n3560# 26.168001f
C62 m3_120_120# m3_4132_120# 0.891312f
C63 c1_n7864_n3560# c1_n7864_160# 0.609898f
C64 c1_4172_n7280# VSUBS 0.735519f
C65 c1_160_n7280# VSUBS 0.735519f
C66 c1_n3852_n7280# VSUBS 0.735519f
C67 c1_n7864_n7280# VSUBS 1.243f
C68 c1_4172_n3560# VSUBS 0.228039f
C69 c1_160_n3560# VSUBS 0.228039f
C70 c1_n3852_n3560# VSUBS 0.228039f
C71 c1_n7864_n3560# VSUBS 0.735519f
C72 c1_4172_160# VSUBS 0.228039f
C73 c1_160_160# VSUBS 0.228039f
C74 c1_n3852_160# VSUBS 0.228039f
C75 c1_n7864_160# VSUBS 0.735519f
C76 c1_4172_3880# VSUBS 0.735519f
C77 c1_160_3880# VSUBS 0.735519f
C78 c1_n3852_3880# VSUBS 0.735519f
C79 c1_n7864_3880# VSUBS 1.243f
C80 m3_4132_n7320# VSUBS 6.48093f
C81 m3_120_n7320# VSUBS 5.35666f
C82 m3_n3892_n7320# VSUBS 5.35666f
C83 m3_n7904_n7320# VSUBS 5.93885f
C84 m3_4132_n3600# VSUBS 5.83462f
C85 m3_120_n3600# VSUBS 4.71035f
C86 m3_n3892_n3600# VSUBS 4.71035f
C87 m3_n7904_n3600# VSUBS 5.29254f
C88 m3_4132_120# VSUBS 5.83462f
C89 m3_120_120# VSUBS 4.71035f
C90 m3_n3892_120# VSUBS 4.71035f
C91 m3_n7904_120# VSUBS 5.29254f
C92 m3_4132_3840# VSUBS 6.48093f
C93 m3_120_3840# VSUBS 5.35666f
C94 m3_n3892_3840# VSUBS 5.35666f
C95 m3_n7904_3840# VSUBS 5.93885f
.ends

.subckt cap_op A B AVSS
Xsky130_fd_pr__cap_mim_m3_1_SXWHWZ_0 AVSS AVSS AVSS AVSS AVSS AVSS B A A AVSS A AVSS
+ A AVSS AVSS AVSS B AVSS AVSS AVSS AVSS B B AVSS AVSS AVSS AVSS AVSS AVSS B AVSS
+ B VSUBS sky130_fd_pr__cap_mim_m3_1_SXWHWZ
C0 A B 3.910106f
C1 B AVSS -0.727581f
C2 A AVSS 1.786197f
C3 A VSUBS 1.201286f
C4 AVSS VSUBS 72.348625f
C5 B VSUBS 24.467958f
.ends

.subckt bgr_op5_block_rev2 AVSS VREF TRIM3 TRIM2 TRIM1 TRIM0 VBGSC VENA VBGTC ENA
+ AVDD DVDD DVSS IPTAT VDDE
Xnmos_startup_0 AVSS pmos_startup_0/D3 pmos_startup_0/D4 nmos_startup
Xresistorstart_0 AVSS AVSS resistorstart_0/A resistorstart
Xpmos_iptat_0 VDDE IPTAT cap_op_0/A pmos_iptat
Xdigital_0 res_trim_0/1 res_trim_0/A TRIM3 res_trim_0/2 TRIM2 TRIM1 TRIM0 res_trim_0/3
+ bjt_0/B VENA VBGTC digital_0/SVBGSC digital_0/SVBGTC AVDD ENA DVDD DVSS VBGSC VDDE
+ digital
Xpmos_startup_0 pmos_startup_0/D3 pmos_startup_0/D4 VDDE resistorstart_0/A pmos_startup
Xres_trim_0 AVSS res_trim_0/A bjt_0/B res_trim_0/3 res_trim_0/2 res_trim_0/1 res_trim
Xpmos_current_bgr_0 VREF resist_const_0/C VDDE resistor_op_tt_0/C cap_op_0/A pmos_current_bgr
Xbjt_0 bjt_0/B bjt_0/A AVSS AVSS AVSS AVSS AVSS AVSS AVSS AVSS AVSS AVSS DVSS AVSS
+ bjt
Xpmos_current_bgr_2_0 nmos_tail_current_0/D2 resistor_op_tt_0/C VDDE differential_pair_0/D4
+ nmos_tail_current_0/D1 pmos_current_bgr_2
Xresistor_op_tt_0 resistor_op_tt_0/A resistor_op_tt_0/C AVSS cap_op_0/B AVSS resistor_op_tt_0/m1_565_4092#
+ resistor_op_tt_0/m1_n99_4131# resistor_op_tt_0/m1_n100_4024# resistor_op_tt
Xnmos_tail_current_0 differential_pair_0/S resistor_op_tt_0/A AVSS nmos_tail_current_0/D1
+ nmos_tail_current_0/D2 cap_op_0/A nmos_tail_current
Xdifferential_pair_0 AVSS differential_pair_0/S resistor_op_tt_0/C differential_pair_0/D4
+ resist_const_0/E bjt_0/A differential_pair
Xresist_const_0 VREF resist_const_0/C resist_const_0/E digital_0/SVBGTC bjt_0/A resist_const_0/E
+ AVSS res_trim_0/A resist_const_0/m1_28308_n3465# resist_const_0/m1_6628_n3631# resist_const_0/m1_19584_n3310#
+ resist_const_0/m1_19584_n3642# resist_const_0/m1_10964_n3465# resist_const_0/m1_15300_n3631#
+ resist_const_0/m1_10964_n3133# resist_const_0/m1_6628_n2469# resist_const_0/m1_15248_n3476#
+ resist_const_0/m1_10912_n3310# resist_const_0/m1_10912_n3642# resist_const_0/m1_6576_n3476#
+ resist_const_0/m1_10964_n2635# resist_const_0/m1_15300_n3299# digital_0/SVBGSC resist_const_0/m1_6628_n3299#
+ resist_const_0/m1_10912_n2812# resist_const_0/m1_15300_n2469# resist_const_0/m1_28256_n3642#
+ resist_const
Xcap_op_0 cap_op_0/A cap_op_0/B AVSS cap_op
C0 res_trim_0/2 bjt_0/B 0.498809f
C1 cap_op_0/A AVSS 7.171165f
C2 VDDE bjt_0/B 0.391695f
C3 TRIM0 VBGSC 0.288642f
C4 differential_pair_0/D4 resistor_op_tt_0/C 0.202707f
C5 resistor_op_tt_0/A AVSS 2.561098f
C6 cap_op_0/A VREF 0.518485f
C7 AVSS resist_const_0/m1_28308_n2967# 0.118204f
C8 cap_op_0/A pmos_startup_0/D3 0.621429f
C9 res_trim_0/2 res_trim_0/3 1.492988f
C10 VDDE res_trim_0/3 3.527917f
C11 TRIM0 ENA 0.187761f
C12 res_trim_0/2 AVSS 4.907239f
C13 VDDE AVSS 1.342642p
C14 bjt_0/A resistor_op_tt_0/C 2.405374f
C15 differential_pair_0/D4 bjt_0/A 1.442522f
C16 VDDE VREF 0.598308f
C17 res_trim_0/2 pmos_startup_0/D3 0.131403f
C18 VDDE pmos_startup_0/D3 0.570423f
C19 res_trim_0/1 resistor_op_tt_0/C 0.107236f
C20 differential_pair_0/D4 res_trim_0/1 0.190838f
C21 VDDE digital_0/SVBGSC 0.460149f
C22 resist_const_0/C AVSS 2.094939f
C23 resist_const_0/m1_28308_n3465# AVSS 0.118205f
C24 res_trim_0/A resistor_op_tt_0/C 0.642042f
C25 resist_const_0/C VREF 1.091755f
C26 res_trim_0/2 TRIM2 0.261291f
C27 resist_const_0/m1_6628_n2801# AVSS 0.108459f
C28 res_trim_0/A differential_pair_0/D4 0.235339f
C29 AVSS resist_const_0/m1_19636_n2635# 0.106973f
C30 bjt_0/A res_trim_0/1 0.995482f
C31 VDDE DVDD 0.218193f
C32 differential_pair_0/S resistor_op_tt_0/C 0.379939f
C33 AVDD AVSS 0.115133f
C34 VENA digital_0/SVBGSC 0.144957f
C35 resist_const_0/m1_10912_n2812# AVSS 0.641906f
C36 differential_pair_0/D4 resist_const_0/E 1.614079f
C37 cap_op_0/B cap_op_0/A 1.038589f
C38 res_trim_0/A bjt_0/A 0.226487f
C39 VBGSC digital_0/SVBGSC 0.179546f
C40 AVSS ENA 0.140855f
C41 res_trim_0/A resist_const_0/m1_15300_n3299# 0.127827f
C42 differential_pair_0/S bjt_0/A 0.341943f
C43 VBGTC digital_0/SVBGSC 0.280586f
C44 nmos_tail_current_0/D1 resistor_op_tt_0/C 0.581049f
C45 pmos_startup_0/D4 bjt_0/A 0.117727f
C46 res_trim_0/A res_trim_0/1 3.366679f
C47 resistor_op_tt_0/C nmos_tail_current_0/D2 0.352447f
C48 differential_pair_0/D4 nmos_tail_current_0/D2 1.421125f
C49 bjt_0/A resist_const_0/E 4.237452f
C50 VDDE digital_0/SVBGTC 0.296104f
C51 resistorstart_0/A bjt_0/A 0.76793f
C52 AVSS resist_const_0/m1_6628_n3631# 0.107567f
C53 bjt_0/B resistor_op_tt_0/C 0.124784f
C54 AVDD DVDD 0.133945f
C55 pmos_startup_0/D4 res_trim_0/1 0.407034f
C56 VBGTC DVDD 0.204855f
C57 AVSS resistor_op_tt_0/m1_n100_4024# 0.222488f
C58 AVSS resist_const_0/m1_10964_n3133# 0.108459f
C59 res_trim_0/1 resist_const_0/E 0.229111f
C60 bjt_0/A nmos_tail_current_0/D1 0.439226f
C61 resist_const_0/m1_15300_n3631# AVSS 0.106973f
C62 resist_const_0/m1_23972_n3631# AVSS 0.107567f
C63 bjt_0/A nmos_tail_current_0/D2 0.24978f
C64 resist_const_0/m1_10912_n3642# AVSS 0.106445f
C65 res_trim_0/A differential_pair_0/S 0.284266f
C66 cap_op_0/A res_trim_0/2 0.154947f
C67 cap_op_0/A VDDE 5.700596f
C68 ENA DVDD 0.145158f
C69 bjt_0/A bjt_0/B 4.985068f
C70 AVSS resistor_op_tt_0/C 2.64832f
C71 nmos_tail_current_0/D1 res_trim_0/1 0.242603f
C72 TRIM3 res_trim_0/1 0.255158f
C73 res_trim_0/A resist_const_0/E 0.349795f
C74 differential_pair_0/D4 AVSS 2.470804f
C75 VREF resistor_op_tt_0/C 0.194581f
C76 differential_pair_0/S resist_const_0/E 0.422873f
C77 resistor_op_tt_0/C pmos_startup_0/D3 0.271361f
C78 bjt_0/B res_trim_0/1 0.561608f
C79 bjt_0/A res_trim_0/3 0.647837f
C80 cap_op_0/A resist_const_0/C 0.243389f
C81 res_trim_0/A nmos_tail_current_0/D1 0.163561f
C82 res_trim_0/2 VDDE 0.366243f
C83 resist_const_0/m1_19636_n3465# AVSS 0.106973f
C84 resist_const_0/m1_23972_n3299# AVSS 0.108459f
C85 resistorstart_0/A resist_const_0/E 0.143558f
C86 res_trim_0/A nmos_tail_current_0/D2 0.840205f
C87 bjt_0/A AVSS 9.397478f
C88 AVSS resist_const_0/m1_6628_n2469# 0.107567f
C89 differential_pair_0/S nmos_tail_current_0/D1 0.111714f
C90 res_trim_0/1 res_trim_0/3 0.333964f
C91 AVSS resist_const_0/m1_15300_n3299# 0.728948f
C92 pmos_startup_0/D4 nmos_tail_current_0/D1 0.488571f
C93 res_trim_0/A resist_const_0/m1_19584_n3310# 0.117608f
C94 bjt_0/A VREF 0.200895f
C95 nmos_tail_current_0/D1 resist_const_0/E 1.193391f
C96 pmos_startup_0/D4 nmos_tail_current_0/D2 0.543903f
C97 bjt_0/A pmos_startup_0/D3 0.332112f
C98 AVSS res_trim_0/1 6.50791f
C99 resist_const_0/E nmos_tail_current_0/D2 1.554255f
C100 resistor_op_tt_0/m1_565_4092# resistor_op_tt_0/C 0.176467f
C101 pmos_startup_0/D4 bjt_0/B 0.531298f
C102 VDDE resist_const_0/C 0.399779f
C103 res_trim_0/A res_trim_0/3 0.614228f
C104 bjt_0/B resist_const_0/E 0.261906f
C105 res_trim_0/1 pmos_startup_0/D3 0.892383f
C106 AVSS resist_const_0/m1_6576_n3476# 0.108554f
C107 res_trim_0/A AVSS 4.935182f
C108 nmos_tail_current_0/D1 nmos_tail_current_0/D2 0.317675f
C109 res_trim_0/1 digital_0/SVBGSC 0.168167f
C110 pmos_startup_0/D4 res_trim_0/3 0.143357f
C111 differential_pair_0/S AVSS 1.708141f
C112 resist_const_0/E res_trim_0/3 0.149112f
C113 bjt_0/A resistor_op_tt_0/m1_565_4092# 0.195588f
C114 resistorstart_0/A res_trim_0/3 1.581278f
C115 VDDE VBGTC 0.151432f
C116 pmos_startup_0/D4 AVSS 1.219642f
C117 bjt_0/B nmos_tail_current_0/D2 0.121734f
C118 AVSS IPTAT 0.920267f
C119 resist_const_0/m1_15300_n2469# AVSS 0.106973f
C120 AVSS resist_const_0/E 9.163497f
C121 res_trim_0/A digital_0/SVBGSC 1.074798f
C122 resistorstart_0/A AVSS 2.419412f
C123 cap_op_0/B resistor_op_tt_0/C 0.154415f
C124 resist_const_0/m1_23972_n2469# AVSS 0.107567f
C125 nmos_tail_current_0/D1 res_trim_0/3 0.10491f
C126 pmos_startup_0/D4 pmos_startup_0/D3 0.144252f
C127 VREF resist_const_0/E 0.156823f
C128 resist_const_0/E pmos_startup_0/D3 0.12938f
C129 nmos_tail_current_0/D2 res_trim_0/3 0.333706f
C130 AVSS nmos_tail_current_0/D1 1.676919f
C131 VENA VBGSC 2.261153f
C132 resist_const_0/m1_15248_n3476# AVSS 0.106445f
C133 bjt_0/B res_trim_0/3 0.212717f
C134 AVSS nmos_tail_current_0/D2 20.311798f
C135 cap_op_0/A resistor_op_tt_0/C 0.87074f
C136 VENA VBGTC 2.684077f
C137 AVSS bjt_0/B 7.643015f
C138 differential_pair_0/D4 cap_op_0/A 0.78978f
C139 nmos_tail_current_0/D1 pmos_startup_0/D3 0.368843f
C140 TRIM0 DVDD 0.15761f
C141 cap_op_0/B bjt_0/A 1.984988f
C142 pmos_startup_0/D3 nmos_tail_current_0/D2 0.31894f
C143 resistor_op_tt_0/A resistor_op_tt_0/C 0.411298f
C144 AVDD VBGTC 0.331837f
C145 differential_pair_0/D4 resistor_op_tt_0/A 0.192912f
C146 digital_0/SVBGTC res_trim_0/1 0.106412f
C147 bjt_0/B pmos_startup_0/D3 0.17632f
C148 TRIM0 TRIM1 3.09903f
C149 cap_op_0/B res_trim_0/1 0.586744f
C150 AVSS res_trim_0/3 12.996652f
C151 bjt_0/B digital_0/SVBGSC 0.125306f
C152 AVDD ENA 0.3239f
C153 cap_op_0/A bjt_0/A 1.341538f
C154 TRIM3 TRIM2 4.093861f
C155 VDDE resistor_op_tt_0/C 0.502873f
C156 differential_pair_0/D4 res_trim_0/2 0.103746f
C157 differential_pair_0/D4 VDDE 0.149202f
C158 AVSS resist_const_0/m1_10964_n2967# 0.108459f
C159 ENA VBGTC 0.273684f
C160 TRIM3 DVDD 5.330606f
C161 res_trim_0/A digital_0/SVBGTC 7.039538f
C162 pmos_startup_0/D3 res_trim_0/3 0.141437f
C163 resistor_op_tt_0/A bjt_0/A 0.224331f
C164 AVSS resist_const_0/m1_10964_n2635# 0.107567f
C165 AVSS VREF 3.399339f
C166 cap_op_0/A res_trim_0/1 0.389119f
C167 res_trim_0/3 digital_0/SVBGSC 0.128463f
C168 AVSS pmos_startup_0/D3 1.208661f
C169 bjt_0/B DVDD 0.195361f
C170 AVSS digital_0/SVBGSC 2.869693f
C171 res_trim_0/2 bjt_0/A 0.292711f
C172 bjt_0/A VDDE 2.374622f
C173 resist_const_0/m1_28256_n3642# AVSS 0.132015f
C174 res_trim_0/A resist_const_0/m1_19584_n3642# 0.115908f
C175 res_trim_0/2 res_trim_0/1 1.047644f
C176 VDDE res_trim_0/1 0.33943f
C177 resist_const_0/m1_2337_n3299# AVSS 0.136252f
C178 AVSS DVDD 0.119514f
C179 pmos_startup_0/D4 cap_op_0/A 0.274708f
C180 cap_op_0/A IPTAT 0.372323f
C181 AVSS resist_const_0/m1_28256_n2812# 0.125005f
C182 bjt_0/A resist_const_0/C 3.262177f
C183 cap_op_0/A resist_const_0/E 0.361874f
C184 TRIM1 res_trim_0/3 0.26517f
C185 cap_op_0/A resistorstart_0/A 1.034035f
C186 res_trim_0/A VDDE 0.653722f
C187 resistor_op_tt_0/A resist_const_0/E 0.17816f
C188 resist_const_0/m1_6628_n3299# AVSS 0.108459f
C189 cap_op_0/B bjt_0/B 0.346223f
C190 differential_pair_0/S res_trim_0/2 0.424584f
C191 resistor_op_tt_0/m1_n99_4131# AVSS 0.247555f
C192 cap_op_0/A nmos_tail_current_0/D1 0.399153f
C193 TRIM0 VDDE 0.119374f
C194 resist_const_0/m1_10912_n3310# AVSS 0.647431f
C195 pmos_startup_0/D4 res_trim_0/2 0.195841f
C196 pmos_startup_0/D4 VDDE 0.108806f
C197 VDDE IPTAT 1.028307f
C198 cap_op_0/A nmos_tail_current_0/D2 0.335763f
C199 res_trim_0/2 resist_const_0/E 3.356485f
C200 VDDE resist_const_0/E 0.39882f
C201 resistorstart_0/A VDDE 0.693687f
C202 cap_op_0/A bjt_0/B 0.604849f
C203 TRIM2 DVDD 0.565581f
C204 AVSS digital_0/SVBGTC 1.154011f
C205 cap_op_0/B AVSS 25.666697f
C206 resistor_op_tt_0/C resistor_op_tt_0/m1_n100_4024# 0.185905f
C207 res_trim_0/2 nmos_tail_current_0/D1 0.860291f
C208 VDDE nmos_tail_current_0/D1 0.341044f
C209 TRIM1 TRIM2 3.594035f
C210 cap_op_0/A res_trim_0/3 0.410506f
C211 res_trim_0/2 nmos_tail_current_0/D2 1.174144f
C212 digital_0/SVBGTC digital_0/SVBGSC 6.821085f
C213 resist_const_0/C resist_const_0/E 0.486932f
C214 TRIM1 DVDD 0.218915f
C215 resistorstart_0/A resist_const_0/C 0.120526f
C216 resist_const_0/m1_10964_n3465# AVSS 0.107567f
C217 cap_op_0/B cap_op_0/VSUBS 21.465908f
C218 resist_const_0/m1_28256_n2812# cap_op_0/VSUBS 0.542836f
C219 resist_const_0/m1_23920_n2646# cap_op_0/VSUBS 0.412976f
C220 resist_const_0/m1_28308_n2967# cap_op_0/VSUBS 0.589905f
C221 resist_const_0/m1_23920_n2978# cap_op_0/VSUBS 0.364019f
C222 resist_const_0/m1_23972_n3299# cap_op_0/VSUBS 0.351297f
C223 resist_const_0/m1_28308_n3465# cap_op_0/VSUBS 0.589905f
C224 resist_const_0/m1_23972_n3631# cap_op_0/VSUBS 0.350405f
C225 resist_const_0/m1_28256_n3642# cap_op_0/VSUBS 0.541353f
C226 resist_const_0/m1_23972_n2303# cap_op_0/VSUBS 0.341828f
C227 resist_const_0/m1_23972_n2469# cap_op_0/VSUBS 0.350405f
C228 resist_const_0/m1_19636_n2635# cap_op_0/VSUBS 0.349811f
C229 resist_const_0/m1_23920_n3144# cap_op_0/VSUBS 0.364018f
C230 resist_const_0/m1_23920_n3476# cap_op_0/VSUBS 0.4124f
C231 resist_const_0/m1_23972_n3797# cap_op_0/VSUBS 0.353369f
C232 resist_const_0/m1_19636_n2303# cap_op_0/VSUBS 0.341828f
C233 resist_const_0/m1_19584_n2480# cap_op_0/VSUBS 0.412973f
C234 resist_const_0/m1_15248_n2646# cap_op_0/VSUBS 0.411441f
C235 resist_const_0/m1_19584_n2812# cap_op_0/VSUBS 0.353548f
C236 resist_const_0/m1_15265_n3133# cap_op_0/VSUBS 0.336237f
C237 resist_const_0/m1_19584_n3310# cap_op_0/VSUBS 0.347065f
C238 resist_const_0/m1_19636_n3465# cap_op_0/VSUBS 0.349811f
C239 resist_const_0/m1_19584_n3642# cap_op_0/VSUBS 0.412397f
C240 resist_const_0/m1_19636_n3797# cap_op_0/VSUBS 0.353369f
C241 resist_const_0/m1_15300_n2303# cap_op_0/VSUBS 0.341828f
C242 resist_const_0/m1_15300_n2469# cap_op_0/VSUBS 0.349811f
C243 digital_0/SVBGSC cap_op_0/VSUBS 2.030241f
C244 resist_const_0/m1_10964_n2967# cap_op_0/VSUBS 0.351297f
C245 resist_const_0/m1_15300_n3299# cap_op_0/VSUBS 1.783432f
C246 resist_const_0/m1_15248_n3476# cap_op_0/VSUBS 0.410865f
C247 resist_const_0/m1_15300_n3631# cap_op_0/VSUBS 0.349811f
C248 resist_const_0/m1_15300_n3797# cap_op_0/VSUBS 0.353369f
C249 resist_const_0/m1_10964_n2303# cap_op_0/VSUBS 0.341828f
C250 resist_const_0/m1_10912_n2480# cap_op_0/VSUBS 0.411444f
C251 resist_const_0/m1_10964_n2635# cap_op_0/VSUBS 0.350405f
C252 resist_const_0/m1_10912_n2812# cap_op_0/VSUBS 1.711577f
C253 resist_const_0/m1_10964_n3133# cap_op_0/VSUBS 0.351297f
C254 resist_const_0/m1_10912_n3310# cap_op_0/VSUBS 1.398506f
C255 resist_const_0/m1_10964_n3465# cap_op_0/VSUBS 0.350405f
C256 resist_const_0/m1_10912_n3642# cap_op_0/VSUBS 0.410868f
C257 resist_const_0/m1_10964_n3797# cap_op_0/VSUBS 0.353369f
C258 resist_const_0/m1_6628_n2303# cap_op_0/VSUBS 0.341828f
C259 resist_const_0/m1_6628_n2469# cap_op_0/VSUBS 0.350405f
C260 resist_const_0/m1_6576_n2646# cap_op_0/VSUBS 0.412976f
C261 resist_const_0/m1_6628_n2801# cap_op_0/VSUBS 0.351297f
C262 resist_const_0/m1_2337_n3299# cap_op_0/VSUBS 0.708589f
C263 resist_const_0/m1_6576_n2978# cap_op_0/VSUBS 0.364019f
C264 resist_const_0/m1_2420_n3133# cap_op_0/VSUBS 0.31019f
C265 resist_const_0/m1_6576_n3144# cap_op_0/VSUBS 0.364018f
C266 resist_const_0/m1_6628_n3299# cap_op_0/VSUBS 0.351297f
C267 resist_const_0/m1_6576_n3476# cap_op_0/VSUBS 0.4124f
C268 resist_const_0/m1_6628_n3631# cap_op_0/VSUBS 0.350405f
C269 resist_const_0/m1_6628_n3797# cap_op_0/VSUBS 0.353369f
C270 resistor_op_tt_0/C cap_op_0/VSUBS 7.696625f
C271 resist_const_0/E cap_op_0/VSUBS 7.064466f
C272 bjt_0/A cap_op_0/VSUBS 4.824366f
C273 differential_pair_0/S cap_op_0/VSUBS 8.474956f
C274 nmos_tail_current_0/D2 cap_op_0/VSUBS 35.11297f
C275 resistor_op_tt_0/A cap_op_0/VSUBS 1.007444f
C276 resistor_op_tt_0/m1_565_4092# cap_op_0/VSUBS 0.333004f
C277 resistor_op_tt_0/m1_n100_4024# cap_op_0/VSUBS 0.831448f
C278 resistor_op_tt_0/m1_n99_4131# cap_op_0/VSUBS 0.714853f
C279 resistor_op_tt_0/m1_n265_4096# cap_op_0/VSUBS 0.335073f
C280 nmos_tail_current_0/D1 cap_op_0/VSUBS 8.260718f
C281 differential_pair_0/D4 cap_op_0/VSUBS 7.176108f
C282 AVSS cap_op_0/VSUBS 0.116637p
C283 cap_op_0/A cap_op_0/VSUBS 19.137087f
C284 VREF cap_op_0/VSUBS 1.475629f
C285 resist_const_0/C cap_op_0/VSUBS 1.335326f
C286 res_trim_0/3 cap_op_0/VSUBS 18.880548f
C287 bjt_0/B cap_op_0/VSUBS 10.604116f
C288 pmos_startup_0/D4 cap_op_0/VSUBS 0.745713f
C289 resistorstart_0/A cap_op_0/VSUBS 2.082616f
C290 VDDE cap_op_0/VSUBS 0.981488p
C291 VBGSC cap_op_0/VSUBS 0.697994f
C292 VENA cap_op_0/VSUBS 0.71676f
C293 digital_0/SVBGTC cap_op_0/VSUBS 0.853344f
C294 VBGTC cap_op_0/VSUBS 0.471028f
C295 TRIM0 cap_op_0/VSUBS 1.031889f
C296 res_trim_0/2 cap_op_0/VSUBS 10.184617f
C297 TRIM1 cap_op_0/VSUBS 0.796594f
C298 res_trim_0/1 cap_op_0/VSUBS 9.457768f
C299 TRIM2 cap_op_0/VSUBS 0.774869f
C300 res_trim_0/A cap_op_0/VSUBS 3.713949f
C301 TRIM3 cap_op_0/VSUBS 0.814072f
C302 AVDD cap_op_0/VSUBS 0.916889f
C303 ENA cap_op_0/VSUBS 1.919369f
C304 DVDD cap_op_0/VSUBS 62.811504f
C305 IPTAT cap_op_0/VSUBS 0.341732f
C306 resistorstart_0/m1_21633_953# cap_op_0/VSUBS 0.358198f
C307 resistorstart_0/m1_21633_621# cap_op_0/VSUBS 0.358198f
C308 resistorstart_0/m1_21633_289# cap_op_0/VSUBS 0.358198f
C309 resistorstart_0/m1_17335_1285# cap_op_0/VSUBS 0.586944f
C310 resistorstart_0/m1_17335_1119# cap_op_0/VSUBS 0.301562f
C311 resistorstart_0/m1_17335_953# cap_op_0/VSUBS 0.301562f
C312 resistorstart_0/m1_17335_787# cap_op_0/VSUBS 0.301562f
C313 resistorstart_0/m1_17335_621# cap_op_0/VSUBS 0.301562f
C314 resistorstart_0/m1_17335_455# cap_op_0/VSUBS 0.301562f
C315 resistorstart_0/m1_17335_289# cap_op_0/VSUBS 0.301562f
C316 resistorstart_0/m1_17335_123# cap_op_0/VSUBS 0.586944f
C317 resistorstart_0/m1_12999_1285# cap_op_0/VSUBS 0.586944f
C318 resistorstart_0/m1_12999_1119# cap_op_0/VSUBS 0.301562f
C319 resistorstart_0/m1_12999_953# cap_op_0/VSUBS 0.301562f
C320 resistorstart_0/m1_12999_787# cap_op_0/VSUBS 0.301562f
C321 resistorstart_0/m1_12999_621# cap_op_0/VSUBS 0.301562f
C322 resistorstart_0/m1_12999_455# cap_op_0/VSUBS 0.301562f
C323 resistorstart_0/m1_12999_289# cap_op_0/VSUBS 0.301562f
C324 resistorstart_0/m1_12999_123# cap_op_0/VSUBS 0.586944f
C325 resistorstart_0/m1_8663_1285# cap_op_0/VSUBS 0.586944f
C326 resistorstart_0/m1_8663_1119# cap_op_0/VSUBS 0.301562f
C327 resistorstart_0/m1_8663_953# cap_op_0/VSUBS 0.301562f
C328 resistorstart_0/m1_8663_787# cap_op_0/VSUBS 0.301562f
C329 resistorstart_0/m1_8663_621# cap_op_0/VSUBS 0.301562f
C330 resistorstart_0/m1_8663_455# cap_op_0/VSUBS 0.301562f
C331 resistorstart_0/m1_8663_289# cap_op_0/VSUBS 0.301562f
C332 resistorstart_0/m1_8663_123# cap_op_0/VSUBS 0.586944f
C333 resistorstart_0/m1_4327_1285# cap_op_0/VSUBS 0.586944f
C334 resistorstart_0/m1_4327_1119# cap_op_0/VSUBS 0.301562f
C335 resistorstart_0/m1_4327_953# cap_op_0/VSUBS 0.301562f
C336 resistorstart_0/m1_119_788# cap_op_0/VSUBS 0.358214f
C337 resistorstart_0/m1_4327_787# cap_op_0/VSUBS 0.301562f
C338 resistorstart_0/m1_4327_621# cap_op_0/VSUBS 0.301562f
C339 resistorstart_0/m1_119_456# cap_op_0/VSUBS 0.358214f
C340 resistorstart_0/m1_4327_455# cap_op_0/VSUBS 0.301562f
C341 resistorstart_0/m1_4327_289# cap_op_0/VSUBS 0.301562f
C342 resistorstart_0/m1_4327_123# cap_op_0/VSUBS 0.586944f
C343 pmos_startup_0/D3 cap_op_0/VSUBS 3.917982f
.ends

