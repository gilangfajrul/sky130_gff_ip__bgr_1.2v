magic
tech sky130A
magscale 1 2
timestamp 1716351939
<< error_p >>
rect -450 552 -380 554
rect -284 552 -214 554
rect -118 552 -48 554
rect 48 552 118 554
rect 214 552 284 554
rect 380 552 450 554
rect -450 -484 -380 -482
rect -284 -484 -214 -482
rect -118 -484 -48 -482
rect 48 -484 118 -482
rect 214 -484 284 -482
rect 380 -484 450 -482
<< nwell >>
rect -643 -1159 643 1159
<< nsubdiff >>
rect -607 1089 -511 1123
rect 511 1089 607 1123
rect -607 1027 -573 1089
rect 573 1027 607 1089
rect -607 -1089 -573 -1027
rect 573 -1089 607 -1027
rect -607 -1123 -511 -1089
rect 511 -1123 607 -1089
<< nsubdiffcont >>
rect -511 1089 511 1123
rect -607 -1027 -573 1027
rect 573 -1027 607 1027
rect -511 -1123 511 -1089
<< xpolycontact >>
rect -450 552 -380 984
rect -450 52 -380 484
rect -284 552 -214 984
rect -284 52 -214 484
rect -118 552 -48 984
rect -118 52 -48 484
rect 48 552 118 984
rect 48 52 118 484
rect 214 552 284 984
rect 214 52 284 484
rect 380 552 450 984
rect 380 52 450 484
rect -450 -484 -380 -52
rect -450 -984 -380 -552
rect -284 -484 -214 -52
rect -284 -984 -214 -552
rect -118 -484 -48 -52
rect -118 -984 -48 -552
rect 48 -484 118 -52
rect 48 -984 118 -552
rect 214 -484 284 -52
rect 214 -984 284 -552
rect 380 -484 450 -52
rect 380 -984 450 -552
<< ppolyres >>
rect -450 484 -380 552
rect -284 484 -214 552
rect -118 484 -48 552
rect 48 484 118 552
rect 214 484 284 552
rect 380 484 450 552
rect -450 -552 -380 -484
rect -284 -552 -214 -484
rect -118 -552 -48 -484
rect 48 -552 118 -484
rect 214 -552 284 -484
rect 380 -552 450 -484
<< locali >>
rect -607 1089 -511 1123
rect 511 1089 607 1123
rect -607 1027 -573 1089
rect 573 1027 607 1089
rect -607 -1089 -573 -1027
rect 573 -1089 607 -1027
rect -607 -1123 -511 -1089
rect 511 -1123 607 -1089
<< viali >>
rect -434 569 -396 966
rect -268 569 -230 966
rect -102 569 -64 966
rect 64 569 102 966
rect 230 569 268 966
rect 396 569 434 966
rect -434 70 -396 467
rect -268 70 -230 467
rect -102 70 -64 467
rect 64 70 102 467
rect 230 70 268 467
rect 396 70 434 467
rect -434 -467 -396 -70
rect -268 -467 -230 -70
rect -102 -467 -64 -70
rect 64 -467 102 -70
rect 230 -467 268 -70
rect 396 -467 434 -70
rect -434 -966 -396 -569
rect -268 -966 -230 -569
rect -102 -966 -64 -569
rect 64 -966 102 -569
rect 230 -966 268 -569
rect 396 -966 434 -569
<< metal1 >>
rect -440 966 -390 978
rect -440 569 -434 966
rect -396 569 -390 966
rect -440 557 -390 569
rect -274 966 -224 978
rect -274 569 -268 966
rect -230 569 -224 966
rect -274 557 -224 569
rect -108 966 -58 978
rect -108 569 -102 966
rect -64 569 -58 966
rect -108 557 -58 569
rect 58 966 108 978
rect 58 569 64 966
rect 102 569 108 966
rect 58 557 108 569
rect 224 966 274 978
rect 224 569 230 966
rect 268 569 274 966
rect 224 557 274 569
rect 390 966 440 978
rect 390 569 396 966
rect 434 569 440 966
rect 390 557 440 569
rect -440 467 -390 479
rect -440 70 -434 467
rect -396 70 -390 467
rect -440 58 -390 70
rect -274 467 -224 479
rect -274 70 -268 467
rect -230 70 -224 467
rect -274 58 -224 70
rect -108 467 -58 479
rect -108 70 -102 467
rect -64 70 -58 467
rect -108 58 -58 70
rect 58 467 108 479
rect 58 70 64 467
rect 102 70 108 467
rect 58 58 108 70
rect 224 467 274 479
rect 224 70 230 467
rect 268 70 274 467
rect 224 58 274 70
rect 390 467 440 479
rect 390 70 396 467
rect 434 70 440 467
rect 390 58 440 70
rect -440 -70 -390 -58
rect -440 -467 -434 -70
rect -396 -467 -390 -70
rect -440 -479 -390 -467
rect -274 -70 -224 -58
rect -274 -467 -268 -70
rect -230 -467 -224 -70
rect -274 -479 -224 -467
rect -108 -70 -58 -58
rect -108 -467 -102 -70
rect -64 -467 -58 -70
rect -108 -479 -58 -467
rect 58 -70 108 -58
rect 58 -467 64 -70
rect 102 -467 108 -70
rect 58 -479 108 -467
rect 224 -70 274 -58
rect 224 -467 230 -70
rect 268 -467 274 -70
rect 224 -479 274 -467
rect 390 -70 440 -58
rect 390 -467 396 -70
rect 434 -467 440 -70
rect 390 -479 440 -467
rect -440 -569 -390 -557
rect -440 -966 -434 -569
rect -396 -966 -390 -569
rect -440 -978 -390 -966
rect -274 -569 -224 -557
rect -274 -966 -268 -569
rect -230 -966 -224 -569
rect -274 -978 -224 -966
rect -108 -569 -58 -557
rect -108 -966 -102 -569
rect -64 -966 -58 -569
rect -108 -978 -58 -966
rect 58 -569 108 -557
rect 58 -966 64 -569
rect 102 -966 108 -569
rect 58 -978 108 -966
rect 224 -569 274 -557
rect 224 -966 230 -569
rect 268 -966 274 -569
rect 224 -978 274 -966
rect 390 -569 440 -557
rect 390 -966 396 -569
rect 434 -966 440 -569
rect 390 -978 440 -966
<< properties >>
string FIXED_BBOX -590 -1106 590 1106
string gencell sky130_fd_pr__res_high_po_0p69
string library sky130
string parameters w 0.350 l 0.50 m 2 nx 6 wmin 0.350 lmin 0.50 rho 319.8 val 1.57k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.350 n_guard 1 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
