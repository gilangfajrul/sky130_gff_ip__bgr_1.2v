magic
tech sky130A
timestamp 1716212328
<< nmos >>
rect -2043 -50 -43 50
rect 43 -50 2043 50
<< ndiff >>
rect -2072 44 -2043 50
rect -2072 -44 -2066 44
rect -2049 -44 -2043 44
rect -2072 -50 -2043 -44
rect -43 44 -14 50
rect -43 -44 -37 44
rect -20 -44 -14 44
rect -43 -50 -14 -44
rect 14 44 43 50
rect 14 -44 20 44
rect 37 -44 43 44
rect 14 -50 43 -44
rect 2043 44 2072 50
rect 2043 -44 2049 44
rect 2066 -44 2072 44
rect 2043 -50 2072 -44
<< ndiffc >>
rect -2066 -44 -2049 44
rect -37 -44 -20 44
rect 20 -44 37 44
rect 2049 -44 2066 44
<< poly >>
rect -2043 50 -43 63
rect 43 50 2043 63
rect -2043 -63 -43 -50
rect 43 -63 2043 -50
<< locali >>
rect -2066 44 -2049 52
rect -2066 -52 -2049 -44
rect -37 44 -20 52
rect -37 -52 -20 -44
rect 20 44 37 52
rect 20 -52 37 -44
rect 2049 44 2066 52
rect 2049 -52 2066 -44
<< viali >>
rect -2066 -44 -2049 44
rect -37 -44 -20 44
rect 20 -44 37 44
rect 2049 -44 2066 44
<< metal1 >>
rect -2069 44 -2046 50
rect -2069 -44 -2066 44
rect -2049 -44 -2046 44
rect -2069 -50 -2046 -44
rect -40 44 -17 50
rect -40 -44 -37 44
rect -20 -44 -17 44
rect -40 -50 -17 -44
rect 17 44 40 50
rect 17 -44 20 44
rect 37 -44 40 44
rect 17 -50 40 -44
rect 2046 44 2069 50
rect 2046 -44 2049 44
rect 2066 -44 2069 44
rect 2046 -50 2069 -44
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 20 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
