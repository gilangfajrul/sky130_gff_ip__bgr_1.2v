magic
tech sky130A
magscale 1 2
timestamp 1716361751
<< metal1 >>
rect 128 3758 258 3808
rect 1164 3758 1304 3808
rect 2214 3758 2354 3808
rect -792 3591 -782 3643
rect -730 3591 -720 3643
rect 62 3584 72 3636
rect 124 3584 134 3636
rect 169 3592 252 3642
rect 169 3476 219 3592
rect 1182 3582 1298 3652
rect 2228 3592 2311 3642
rect 136 3426 219 3476
rect -794 3393 -744 3426
rect 254 3425 264 3477
rect 316 3425 326 3477
rect 1108 3425 1118 3477
rect 1170 3425 1180 3477
rect 1300 3425 1310 3477
rect 1362 3425 1372 3477
rect 2154 3425 2164 3477
rect 2216 3425 2226 3477
rect 2261 3476 2311 3592
rect 2346 3591 2356 3643
rect 2408 3591 2418 3643
rect 3200 3591 3210 3643
rect 3262 3591 3272 3643
rect 2261 3426 2344 3476
rect 3224 3393 3274 3432
rect -794 3343 3274 3393
rect 124 3260 254 3310
rect 1176 3260 1316 3310
rect 2216 3260 2356 3310
<< via1 >>
rect -782 3591 -730 3643
rect 72 3584 124 3636
rect 264 3425 316 3477
rect 1118 3425 1170 3477
rect 1310 3425 1362 3477
rect 2164 3425 2216 3477
rect 2356 3591 2408 3643
rect 3210 3591 3262 3643
<< metal2 >>
rect -782 3674 2408 3726
rect -782 3643 -730 3674
rect -782 3581 -730 3591
rect 70 3636 126 3646
rect 70 3570 126 3580
rect 168 3562 220 3674
rect 1214 3562 1266 3674
rect 2356 3643 2408 3674
rect 2356 3581 2408 3591
rect 3208 3645 3264 3655
rect 3208 3579 3264 3589
rect 168 3510 316 3562
rect 1214 3510 1362 3562
rect 264 3477 316 3510
rect 264 3415 316 3425
rect 1118 3477 1170 3487
rect 1118 3415 1170 3425
rect 1310 3477 1362 3510
rect 1310 3415 1362 3425
rect 2162 3479 2218 3489
rect 2162 3413 2218 3423
<< via2 >>
rect 70 3584 72 3636
rect 72 3584 124 3636
rect 124 3584 126 3636
rect 70 3580 126 3584
rect 3208 3643 3264 3645
rect 3208 3591 3210 3643
rect 3210 3591 3262 3643
rect 3262 3591 3264 3643
rect 3208 3589 3264 3591
rect 2162 3477 2218 3479
rect 2162 3425 2164 3477
rect 2164 3425 2216 3477
rect 2216 3425 2218 3477
rect 2162 3423 2218 3425
<< metal3 >>
rect 42 3636 142 3667
rect 42 3580 70 3636
rect 126 3580 142 3636
rect 42 3564 142 3580
rect 3180 3645 3280 3667
rect 3180 3589 3208 3645
rect 3264 3589 3280 3645
rect 3180 3564 3280 3589
rect 42 3504 3280 3564
rect 2134 3479 2234 3504
rect 2134 3423 2162 3479
rect 2218 3423 2234 3479
rect 2134 3401 2234 3423
use sky130_fd_pr__res_high_po_0p35_VSLXGP  sky130_fd_pr__res_high_po_0p35_VSLXGP_0
timestamp 1716351939
transform 0 1 1240 -1 0 3534
box -284 -2040 284 2040
<< end >>
