magic
tech sky130A
magscale 1 2
timestamp 1716188352
<< nwell >>
rect -2181 -162 2181 162
<< pmos >>
rect -2087 -100 -1087 100
rect -1029 -100 -29 100
rect 29 -100 1029 100
rect 1087 -100 2087 100
<< pdiff >>
rect -2145 88 -2087 100
rect -2145 -88 -2133 88
rect -2099 -88 -2087 88
rect -2145 -100 -2087 -88
rect -1087 88 -1029 100
rect -1087 -88 -1075 88
rect -1041 -88 -1029 88
rect -1087 -100 -1029 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 1029 88 1087 100
rect 1029 -88 1041 88
rect 1075 -88 1087 88
rect 1029 -100 1087 -88
rect 2087 88 2145 100
rect 2087 -88 2099 88
rect 2133 -88 2145 88
rect 2087 -100 2145 -88
<< pdiffc >>
rect -2133 -88 -2099 88
rect -1075 -88 -1041 88
rect -17 -88 17 88
rect 1041 -88 1075 88
rect 2099 -88 2133 88
<< poly >>
rect -2087 100 -1087 126
rect -1029 100 -29 126
rect 29 100 1029 126
rect 1087 100 2087 126
rect -2087 -126 -1087 -100
rect -1029 -126 -29 -100
rect 29 -126 1029 -100
rect 1087 -126 2087 -100
<< locali >>
rect -2133 88 -2099 104
rect -2133 -104 -2099 -88
rect -1075 88 -1041 104
rect -1075 -104 -1041 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 1041 88 1075 104
rect 1041 -104 1075 -88
rect 2099 88 2133 104
rect 2099 -104 2133 -88
<< viali >>
rect -2133 -88 -2099 88
rect -1075 -88 -1041 88
rect -17 -88 17 88
rect 1041 -88 1075 88
rect 2099 -88 2133 88
<< metal1 >>
rect -2139 88 -2093 100
rect -2139 -88 -2133 88
rect -2099 -88 -2093 88
rect -2139 -100 -2093 -88
rect -1081 88 -1035 100
rect -1081 -88 -1075 88
rect -1041 -88 -1035 88
rect -1081 -100 -1035 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 1035 88 1081 100
rect 1035 -88 1041 88
rect 1075 -88 1081 88
rect 1035 -100 1081 -88
rect 2093 88 2139 100
rect 2093 -88 2099 88
rect 2133 -88 2139 88
rect 2093 -100 2139 -88
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 5 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
