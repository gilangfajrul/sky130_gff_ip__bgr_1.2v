magic
tech sky130A
magscale 1 2
timestamp 1717694033
<< nwell >>
rect -2123 -164 2123 198
<< pmos >>
rect -2029 -64 -29 136
rect 29 -64 2029 136
<< pdiff >>
rect -2087 124 -2029 136
rect -2087 -52 -2075 124
rect -2041 -52 -2029 124
rect -2087 -64 -2029 -52
rect -29 124 29 136
rect -29 -52 -17 124
rect 17 -52 29 124
rect -29 -64 29 -52
rect 2029 124 2087 136
rect 2029 -52 2041 124
rect 2075 -52 2087 124
rect 2029 -64 2087 -52
<< pdiffc >>
rect -2075 -52 -2041 124
rect -17 -52 17 124
rect 2041 -52 2075 124
<< poly >>
rect -2029 136 -29 162
rect 29 136 2029 162
rect -2029 -111 -29 -64
rect -2029 -145 -2013 -111
rect -45 -145 -29 -111
rect -2029 -161 -29 -145
rect 29 -111 2029 -64
rect 29 -145 45 -111
rect 2013 -145 2029 -111
rect 29 -161 2029 -145
<< polycont >>
rect -2013 -145 -45 -111
rect 45 -145 2013 -111
<< locali >>
rect -2075 124 -2041 140
rect -2075 -68 -2041 -52
rect -17 124 17 140
rect -17 -68 17 -52
rect 2041 124 2075 140
rect 2041 -68 2075 -52
rect -2029 -145 -2013 -111
rect -45 -145 -29 -111
rect 29 -145 45 -111
rect 2013 -145 2029 -111
<< viali >>
rect -2075 -52 -2041 124
rect -17 -52 17 124
rect 2041 -52 2075 124
rect -1521 -145 -537 -111
rect 537 -145 1521 -111
<< metal1 >>
rect -2081 124 -2035 136
rect -2081 -52 -2075 124
rect -2041 -52 -2035 124
rect -2081 -64 -2035 -52
rect -23 124 23 136
rect -23 -52 -17 124
rect 17 -52 23 124
rect -23 -64 23 -52
rect 2035 124 2081 136
rect 2035 -52 2041 124
rect 2075 -52 2081 124
rect 2035 -64 2081 -52
rect -1533 -111 -525 -105
rect -1533 -145 -1521 -111
rect -537 -145 -525 -111
rect -1533 -151 -525 -145
rect 525 -111 1533 -105
rect 525 -145 537 -111
rect 1521 -145 1533 -111
rect 525 -151 1533 -145
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 10 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 50 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
