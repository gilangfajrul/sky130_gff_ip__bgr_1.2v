magic
tech sky130A
magscale 1 2
timestamp 1717768872
<< nwell >>
rect -323 -298 323 264
<< pmos >>
rect -229 -236 -29 164
rect 29 -236 229 164
<< pdiff >>
rect -287 152 -229 164
rect -287 -224 -275 152
rect -241 -224 -229 152
rect -287 -236 -229 -224
rect -29 152 29 164
rect -29 -224 -17 152
rect 17 -224 29 152
rect -29 -236 29 -224
rect 229 152 287 164
rect 229 -224 241 152
rect 275 -224 287 152
rect 229 -236 287 -224
<< pdiffc >>
rect -275 -224 -241 152
rect -17 -224 17 152
rect 241 -224 275 152
<< poly >>
rect -187 245 -71 261
rect -187 228 -171 245
rect -229 211 -171 228
rect -87 228 -71 245
rect 71 245 187 261
rect 71 228 87 245
rect -87 211 -29 228
rect -229 164 -29 211
rect 29 211 87 228
rect 171 228 187 245
rect 171 211 229 228
rect 29 164 229 211
rect -229 -262 -29 -236
rect 29 -262 229 -236
<< polycont >>
rect -171 211 -87 245
rect 87 211 171 245
<< locali >>
rect -187 211 -171 245
rect -87 211 -71 245
rect 71 211 87 245
rect 171 211 187 245
rect -275 152 -241 168
rect -275 -240 -241 -224
rect -17 152 17 168
rect -17 -240 17 -224
rect 241 152 275 168
rect 241 -240 275 -224
<< viali >>
rect -171 211 -87 245
rect 87 211 171 245
rect -275 -224 -241 152
rect -17 -224 17 152
rect 241 -224 275 152
<< metal1 >>
rect -183 245 -75 251
rect -183 211 -171 245
rect -87 211 -75 245
rect -183 205 -75 211
rect 75 245 183 251
rect 75 211 87 245
rect 171 211 183 245
rect 75 205 183 211
rect -281 152 -235 164
rect -281 -224 -275 152
rect -241 -224 -235 152
rect -281 -236 -235 -224
rect -23 152 23 164
rect -23 -224 -17 152
rect 17 -224 23 152
rect -23 -236 23 -224
rect 235 152 281 164
rect 235 -224 241 152
rect 275 -224 281 152
rect 235 -236 281 -224
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2 l 1 m 1 nf 2 diffcov 100 polycov 50 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
