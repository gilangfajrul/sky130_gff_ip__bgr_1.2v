magic
tech sky130A
magscale 1 2
timestamp 1717260083
<< psubdiff >>
rect -218 507 -158 541
rect 4316 507 4376 541
rect -218 481 -184 507
rect 4342 481 4376 507
rect -218 -627 -184 -601
rect 4342 -627 4376 -601
rect -218 -661 -158 -627
rect 4316 -661 4376 -627
<< psubdiffcont >>
rect -158 507 4316 541
rect -218 -601 -184 481
rect 4342 -601 4376 481
rect -158 -661 4316 -627
<< poly >>
rect -38 65 -8 87
rect -100 49 -8 65
rect -100 15 -84 49
rect -50 15 -8 49
rect -100 -1 -8 15
rect 4166 65 4196 87
rect 4166 49 4258 65
rect 4166 15 4208 49
rect 4242 15 4258 49
rect 4166 -1 4258 15
rect -100 -135 -8 -119
rect -100 -169 -84 -135
rect -50 -169 -8 -135
rect -100 -185 -8 -169
rect 4166 -135 4258 -119
rect 4166 -169 4208 -135
rect 4242 -169 4258 -135
rect 4166 -185 4258 -169
rect -38 -207 -8 -185
<< polycont >>
rect -84 15 -50 49
rect 4208 15 4242 49
rect -84 -169 -50 -135
rect 4208 -169 4242 -135
<< locali >>
rect -218 507 -158 541
rect 4316 507 4376 541
rect -218 481 -184 507
rect 4342 481 4376 507
rect -84 49 -50 87
rect -84 -1 -50 15
rect 4208 49 4242 87
rect 4208 -1 4242 15
rect -84 -135 -50 -119
rect -84 -207 -50 -169
rect 4208 -135 4242 -119
rect 4208 -244 4242 -169
rect -218 -627 -184 -601
rect 4342 -627 4376 -601
rect -218 -661 -158 -627
rect 4316 -661 4376 -627
<< viali >>
rect -218 3 -184 37
rect -84 15 -50 49
rect 4208 15 4242 49
rect 4342 15 4376 49
rect -218 -169 -184 -135
rect -84 -169 -50 -135
rect 4208 -169 4242 -135
rect 4342 -169 4376 -135
<< metal1 >>
rect -182 430 -172 482
rect -120 479 -110 482
rect 4268 479 4278 482
rect -120 433 4278 479
rect -120 430 -110 433
rect 2056 320 2102 433
rect 4268 430 4278 433
rect 4330 430 4340 482
rect -15 99 -5 315
rect 47 99 57 315
rect 2062 99 2096 320
rect -90 49 -44 87
rect -224 37 -84 49
rect -224 3 -218 37
rect -184 15 -84 37
rect -50 15 -44 49
rect -184 3 -44 15
rect 548 6 558 58
rect 1542 6 1552 58
rect 2606 6 2616 58
rect 3600 6 3610 58
rect -224 -9 -66 3
rect 4114 -37 4160 120
rect 4202 61 4248 87
rect 4202 49 4382 61
rect 4202 15 4208 49
rect 4242 15 4342 49
rect 4376 15 4382 49
rect 4202 3 4382 15
rect -2 -83 4160 -37
rect -224 -135 -44 -123
rect -224 -169 -218 -135
rect -184 -169 -84 -135
rect -50 -169 -44 -135
rect -224 -181 -44 -169
rect -90 -207 -44 -181
rect -2 -214 44 -83
rect 548 -178 558 -126
rect 1542 -178 1552 -126
rect 2606 -178 2616 -126
rect 3600 -178 3610 -126
rect 4202 -135 4382 -123
rect 4202 -169 4208 -135
rect 4242 -169 4342 -135
rect 4376 -169 4382 -135
rect 4202 -181 4382 -169
rect -182 -602 -172 -550
rect -120 -553 -110 -550
rect 2056 -553 2102 -207
rect 4101 -435 4111 -219
rect 4163 -435 4173 -219
rect 4202 -240 4248 -181
rect 4268 -553 4278 -550
rect -120 -599 4278 -553
rect -120 -602 -110 -599
rect 4268 -602 4278 -599
rect 4330 -602 4340 -550
<< via1 >>
rect -172 430 -120 482
rect 4278 430 4330 482
rect -5 99 47 315
rect 558 6 1542 58
rect 2616 6 3600 58
rect 558 -178 1542 -126
rect 2616 -178 3600 -126
rect -172 -602 -120 -550
rect 4111 -435 4163 -219
rect 4278 -602 4330 -550
<< metal2 >>
rect -172 482 -120 492
rect -172 -550 -120 430
rect 4278 482 4330 492
rect -5 315 47 325
rect -5 -34 47 99
rect 558 60 1542 70
rect 558 -6 1542 4
rect 2616 60 3600 70
rect 2616 -6 3600 4
rect -5 -86 4163 -34
rect 558 -124 1542 -114
rect 558 -190 1542 -180
rect 2616 -124 3600 -114
rect 2616 -190 3600 -180
rect 4111 -219 4163 -86
rect 4111 -445 4163 -435
rect -172 -612 -120 -602
rect 4278 -550 4330 430
rect 4278 -612 4330 -602
<< via2 >>
rect 558 58 1542 60
rect 558 6 1542 58
rect 558 4 1542 6
rect 2616 58 3600 60
rect 2616 6 3600 58
rect 2616 4 3600 6
rect 558 -126 1542 -124
rect 558 -178 1542 -126
rect 558 -180 1542 -178
rect 2616 -126 3600 -124
rect 2616 -178 3600 -126
rect 2616 -180 3600 -178
<< metal3 >>
rect 548 64 1552 65
rect 548 0 558 64
rect 1542 0 1552 64
rect 548 -1 1552 0
rect 2046 60 3610 65
rect 2046 4 2616 60
rect 3600 4 3610 60
rect 2046 -1 3610 4
rect 2046 -119 2112 -1
rect 548 -124 2112 -119
rect 548 -180 558 -124
rect 1542 -180 2112 -124
rect 548 -185 2112 -180
rect 2606 -120 3610 -119
rect 2606 -184 2616 -120
rect 3600 -184 3610 -120
rect 2606 -185 3610 -184
<< via3 >>
rect 558 60 1542 64
rect 558 4 1542 60
rect 558 0 1542 4
rect 2616 -124 3600 -120
rect 2616 -180 3600 -124
rect 2616 -184 3600 -180
<< metal4 >>
rect 557 64 1543 65
rect 557 0 558 64
rect 1542 0 2111 64
rect 557 -1 1543 0
rect 2047 -120 2111 0
rect 2615 -120 3601 -119
rect 2047 -184 2616 -120
rect 3600 -184 3601 -120
rect 2615 -185 3601 -184
use sky130_fd_pr__nfet_01v8_BHCXYW  sky130_fd_pr__nfet_01v8_BHCXYW_0
timestamp 1717258959
transform 1 0 2079 0 1 -327
box -2087 -208 2087 208
use sky130_fd_pr__nfet_01v8_BHCXYW  sky130_fd_pr__nfet_01v8_BHCXYW_1
timestamp 1717258959
transform 1 0 2079 0 1 207
box -2087 -208 2087 208
use sky130_fd_pr__nfet_01v8_HB7GG4  sky130_fd_pr__nfet_01v8_HB7GG4_1
timestamp 1717259999
transform 1 0 -23 0 1 -327
box -73 -146 73 146
use sky130_fd_pr__nfet_01v8_HB7GG4  sky130_fd_pr__nfet_01v8_HB7GG4_2
timestamp 1717259999
transform 1 0 -23 0 1 207
box -73 -146 73 146
use sky130_fd_pr__nfet_01v8_HB7GG4  sky130_fd_pr__nfet_01v8_HB7GG4_3
timestamp 1717259999
transform 1 0 4181 0 1 207
box -73 -146 73 146
use sky130_fd_pr__nfet_01v8_HB7GG4  sky130_fd_pr__nfet_01v8_HB7GG4_4
timestamp 1717259999
transform 1 0 4181 0 1 -327
box -73 -146 73 146
<< labels >>
flabel metal2 4130 -134 4130 -134 0 FreeSans 160 0 0 0 D3
port 1 nsew
flabel metal1 4136 25 4136 25 0 FreeSans 160 0 0 0 D4
port 2 nsew
flabel metal1 2081 -575 2081 -575 0 FreeSans 160 0 0 0 S
port 3 nsew
flabel psubdiffcont 2018 -642 2018 -642 0 FreeSans 160 0 0 0 GND
port 5 nsew
flabel metal4 2206 -137 2206 -137 0 FreeSans 160 0 0 0 plus
port 6 nsew
flabel metal3 2176 16 2176 16 0 FreeSans 160 0 0 0 minus
port 8 nsew
<< end >>
