** sch_path: /foss/pdks/ciel/sky130/versions/8afc8346a57fe1ab7934ba5a6056ea8b43078e71/sky130A/libs.tech/xschem/sky130_tests/test_nmos.sch
**.subckt test_nmos G1v8 D1v8 B
*.ipin G1v8
*.ipin D1v8
*.ipin B
Vd1 D1v8 net1 0
.save i(vd1)
Vd3 D3v3 net2 0
.save i(vd3)
Vd2 D1v8 net3 0
.save i(vd2)
Vd4 D5v0 net4 0
.save i(vd4)
E1 D5v0 0 D1v8 0 '5/1.8'
E2 D3v3 0 D1v8 0 '3.3/1.8'
E3 G5v0 0 G1v8 0 '5/1.8'
E4 G3v3 0 G1v8 0 '3.3/1.8'
Vd5 D10v5 net5 0
.save i(vd5)
E5 D10v5 0 D1v8 0 '10.5/1.8'
E6 D16v0 0 D1v8 0 '16.0/1.8'
Vd6 D16v0 net6 0
.save i(vd6)
Vd7 D1v8 net7 0
.save i(vd7)
E7 D20v0 0 D1v8 0 '20.0/1.8'
XM1 net1 G1v8 S B sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0
+ mult=1 m=1
XM2 net3 G1v8 S B sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0 mult=1
+ m=1
XM3 net2 G3v3 S B sky130_fd_pr__nfet_03v3_nvt L=0.5 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0
+ mult=1 m=1
XM4 net4 G5v0 S B sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0
+ mult=1 m=1
XM5 net5 G5v0 S B sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0
+ mult=1 m=1
XM6 net6 G5v0 S B sky130_fd_pr__nfet_g5v0d16v0 L=0.7 W=5.0 nf=1 ad=1.45 as=1.45 pd=10.58 ps=10.58 nrd=0.058 nrs=0.058 sa=0 sb=0
+ sd=0 mult=1 m=1
Vd8 D1v8 net8 0
.save i(vd8)
XM7 net7 G1v8 S B sky130_fd_pr__nfet_20v0 L=0.5 W=40 m=1
XM8 net8 G1v8 S B sky130_fd_pr__nfet_20v0_zvt W=60 L=0.5 m=1
Vd9 D1v8 net9 0
.save i(vd9)
XM9 net9 G1v8 S B sky130_fd_pr__nfet_01v8_lvt L=0.15 W='0.5 * 2 ' nf=2 ad=0.0725 as=0.145 pd=1.08 ps=2.16 nrd=0.58 nrs=0.58 sa=0 sb=0
+ sd=0 mult=1 m=1
Vd10 D1v8 net10 0
.save i(vd10)
Vd11 D1v8 net12 0
.save i(vd11)
Vd12 D3v3 net11 0
.save i(vd12)
Vd13 D5v0 net13 0
.save i(vd13)
Vd14 D10v5 net14 0
.save i(vd14)
Vd15 D16v0 net15 0
.save i(vd15)
Vd16 D1v8 net16 0
.save i(vd16)
XM10 net10 G1v8 S B sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0
+ mult=1 m=1
XM11 net12 G1v8 S B sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0
+ mult=1 m=1
XM12 net11 G3v3 S B sky130_fd_pr__nfet_03v3_nvt L=0.5 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0
+ mult=1 m=1
XM13 net13 G5v0 S B sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0
+ mult=1 m=1
XM14 net14 G5v0 S B sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0
+ mult=1 m=1
XM15 net15 G5v0 S B sky130_fd_pr__nfet_g5v0d16v0 L=0.7 W=5.0 nf=1 ad=1.45 as=1.45 pd=10.58 ps=10.58 nrd=0.058 nrs=0.058 sa=0 sb=0
+ sd=0 mult=1 m=1
XM16 net16 G1v8 S B sky130_fd_pr__nfet_20v0 L=0.5 W=40 m=1
XM32 net17 G5v0 S B sky130_fd_pr__esd_nfet_05v0_nvt L=2 W=10 nf=1 ad=2.9 as=2.9 pd=20.58 ps=20.58 nrd=0.029 nrs=0.029 sa=0 sb=0
+ sd=0 mult=1 m=1
Vd17 D5v0 net17 0
.save i(vd17)
**** begin user architecture code

* this option enables mos model bin
* selection based on W/NF instead of W
.option wnflag=1
.option savecurrents
vg G1v8 0 1.8
vs s 0 0
vd D1v8 0 1.8
vb b 0 0
.control
save all
save @m.xm9.msky130_fd_pr__nfet_01v8_lvt[gm]
save @m.xm8.m1[gm]
save @m.xm7.m1[gm]
save @m.xm6.xmain1.msky130_fd_pr__nfet_g5v0d16v0__base[gm]
save @m.xm6.xsky130_fd_pr__nfet_g5v0d16v0.msky130_fd_pr__nfet_g5v0d16v0_base[gm]
save @m.xm5.msky130_fd_pr__nfet_g5v0d10v5[gm]
save @m.xm4.msky130_fd_pr__nfet_05v0_nvt[gm]
save @m.xm3.msky130_fd_pr__nfet_03v3_nvt[gm]
save @m.xm2.msky130_fd_pr__nfet_01v8[gm]
save @m.xm1.msky130_fd_pr__nfet_01v8_lvt[gm]
save @m.xm16.m1[gm]
save @m.xm15.xsky130_fd_pr__nfet_g5v0d16v0.msky130_fd_pr__nfet_g5v0d16v0_base[gm]
save @m.xm14.msky130_fd_pr__nfet_g5v0d10v5[gm]
save @m.xm13.msky130_fd_pr__nfet_05v0_nvt[gm]
save @m.xm12.msky130_fd_pr__nfet_03v3_nvt[gm]
save @m.xm11.msky130_fd_pr__nfet_01v8[gm]
save @m.xm10.msky130_fd_pr__nfet_01v8_lvt[gm]
dc vd 0 1.8 0.005 vg 0 1.8 0.2
write test_nmos.raw
* dc vd 0 1.8 0.001 vg 0 1.2 0.1
plot all.vd1#branch vs D1v8
*plot all.vd2#branch vs D1v8
plot all.vd3#branch vs D3v3
*plot all.vd4#branch vs D5v0
plot all.vd5#branch vs D10v5
*plot all.vd6#branch vs D16v0
plot all.vd8#branch vs D1v8
plot all.vd7#branch vs D1v8
set appendwrite
op
write test_nmos.raw
quit 0
.endc


.lib /foss/pdks/sky130A/libs.tech/combined/sky130.lib.spice tt
**** end user architecture code
**.ends
.end
