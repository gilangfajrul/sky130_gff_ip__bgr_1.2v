magic
tech sky130A
magscale 1 2
timestamp 1717870769
<< viali >>
rect -259 5446 -221 5480
rect 571 5446 609 5480
rect -259 2252 -221 2286
rect 571 2252 609 2286
<< metal1 >>
rect -271 5480 -209 5486
rect -271 5446 -259 5480
rect -221 5446 -209 5480
rect -271 5440 -209 5446
rect 559 5480 621 5486
rect 559 5446 571 5480
rect 609 5446 621 5480
rect 559 5440 621 5446
rect -265 5334 -215 5440
rect -99 5377 449 5427
rect -99 5332 -49 5377
rect 56 5292 66 5344
rect 118 5292 128 5344
rect 222 5292 232 5344
rect 284 5292 294 5344
rect 399 5332 449 5377
rect 565 5339 615 5440
rect -265 3803 -215 3950
rect 56 3924 66 3976
rect 118 3924 128 3976
rect 222 3924 232 3976
rect 284 3924 294 3976
rect -99 3892 -49 3924
rect 399 3892 449 3927
rect -99 3842 449 3892
rect -110 3756 -100 3808
rect -48 3756 -38 3808
rect 67 3802 117 3842
rect 233 3798 283 3842
rect 388 3756 398 3808
rect 450 3756 460 3808
rect 565 3792 615 3939
rect -265 2292 -215 2399
rect -110 2388 -100 2440
rect -48 2388 -38 2440
rect 66 2355 116 2400
rect 233 2355 283 2400
rect 388 2388 398 2440
rect 450 2388 460 2440
rect 66 2305 283 2355
rect 565 2292 615 2425
rect -271 2286 -209 2292
rect -271 2252 -259 2286
rect -221 2252 -209 2286
rect -271 2246 -209 2252
rect 559 2286 621 2292
rect 559 2252 571 2286
rect 609 2252 621 2286
rect 559 2246 621 2252
<< via1 >>
rect 66 5292 118 5344
rect 232 5292 284 5344
rect 66 3924 118 3976
rect 232 3924 284 3976
rect -100 3756 -48 3808
rect 398 3756 450 3808
rect -100 2388 -48 2440
rect 398 2388 450 2440
<< metal2 >>
rect 66 5376 533 5428
rect 66 5344 118 5376
rect 66 5282 118 5292
rect 232 5344 284 5376
rect 232 5282 284 5292
rect 66 3976 118 3986
rect 66 3893 118 3924
rect 232 3976 284 3986
rect 232 3893 284 3924
rect -100 3841 450 3893
rect -100 3808 -48 3841
rect -100 3746 -48 3756
rect 398 3808 450 3841
rect 398 3746 450 3756
rect -100 2440 -48 2450
rect -100 2352 -48 2388
rect 398 2440 450 2450
rect 398 2352 450 2388
rect 481 2352 533 5376
rect -100 2300 533 2352
use sky130_fd_pr__res_high_po_0p35_4E8R5J  sky130_fd_pr__res_high_po_0p35_4E8R5J_0
timestamp 1717269017
transform 1 0 175 0 1 3866
box -616 -1650 616 1650
<< labels >>
flabel metal2 501 3866 501 3866 0 FreeSans 160 0 0 0 A
port 0 nsew
flabel metal2 259 3901 259 3901 0 FreeSans 160 0 0 0 B
port 1 nsew
flabel metal1 98 2361 98 2361 0 FreeSans 160 0 0 0 C
port 2 nsew
flabel metal1 -11 5410 -11 5410 0 FreeSans 160 0 0 0 D
port 4 nsew
flabel metal1 -244 5418 -244 5418 0 FreeSans 1600 0 0 0 AVSS
port 5 nsew
<< end >>
