magic
tech sky130A
magscale 1 2
timestamp 1762795171
<< metal1 >>
rect 16812 2790 16822 2842
rect 18106 2790 18116 2842
rect 9397 -1310 9407 -1238
rect 9479 -1310 19295 -1238
rect 19367 -1310 19377 -1238
rect 4529 -2291 4581 -2285
rect 4581 -2343 26555 -2291
rect 26607 -2343 26613 -2291
rect 4529 -2349 4581 -2343
rect 26778 -2544 26830 -2538
rect 8635 -2596 8645 -2544
rect 8697 -2596 26778 -2544
rect 26830 -2596 26840 -2544
rect 26778 -2602 26830 -2596
rect 9406 -2760 9416 -2704
rect 9472 -2760 9482 -2704
rect 19296 -4813 19368 -4807
rect 8985 -4885 8991 -4813
rect 9063 -4885 19296 -4813
rect 19296 -4891 19368 -4885
rect 26329 -4939 26339 -4938
rect 18892 -5012 18902 -4940
rect 18974 -5012 26339 -4939
rect 26411 -5010 26421 -4938
rect 17287 -5184 17297 -5108
rect 17373 -5184 25868 -5108
rect 25944 -5184 25954 -5108
rect 25626 -5645 25636 -5593
rect 26033 -5645 26043 -5593
rect 25626 -5811 25636 -5759
rect 26033 -5811 26043 -5759
rect 8819 -6309 8829 -6257
rect 9226 -6309 9236 -6257
rect 25626 -6641 25636 -6589
rect 26033 -6641 26043 -6589
rect 25626 -6807 25636 -6755
rect 26033 -6807 26043 -6755
<< via1 >>
rect 16822 2790 18106 2842
rect 9407 -1310 9479 -1238
rect 19295 -1310 19367 -1238
rect 4529 -2343 4581 -2291
rect 26555 -2343 26607 -2291
rect 8645 -2596 8697 -2544
rect 26778 -2596 26830 -2544
rect 9416 -2760 9472 -2704
rect 8991 -4885 9063 -4813
rect 19296 -4885 19368 -4813
rect 18902 -5012 18974 -4940
rect 26339 -5010 26411 -4938
rect 17297 -5184 17373 -5108
rect 25868 -5184 25944 -5108
rect 25636 -5645 26033 -5593
rect 25636 -5811 26033 -5759
rect 8829 -6309 9226 -6257
rect 25636 -6641 26033 -6589
rect 25636 -6807 26033 -6755
<< metal2 >>
rect 18084 2928 19374 2986
rect 16822 2845 18106 2852
rect 16822 2842 18978 2845
rect 18106 2790 18978 2842
rect 16822 2787 18978 2790
rect 16822 2780 18106 2787
rect 9034 1546 9095 1549
rect 9027 1490 9036 1546
rect 9092 1490 9101 1546
rect 9034 -1267 9095 1490
rect 8754 -1328 9095 -1267
rect 9407 -1238 9479 -1228
rect 4529 -2291 4581 -1340
rect 4523 -2343 4529 -2291
rect 4581 -2343 4587 -2291
rect 8645 -2544 8697 -1413
rect 8645 -2606 8697 -2596
rect 9407 -2704 9479 -1310
rect 9415 -2760 9416 -2704
rect 9472 -2760 9473 -2704
rect 9415 -2761 9473 -2760
rect 9416 -2770 9472 -2761
rect 8991 -4813 9063 -4807
rect 8991 -6247 9063 -4885
rect 18898 -4940 18978 2787
rect 19290 -1238 19374 2928
rect 19290 -1310 19295 -1238
rect 19367 -1310 19374 -1238
rect 19290 -4813 19374 -1310
rect 19290 -4885 19296 -4813
rect 19368 -4885 19374 -4813
rect 26555 -2291 26607 -2285
rect 18898 -5012 18902 -4940
rect 18974 -5012 18978 -4940
rect 18898 -5022 18978 -5012
rect 26339 -4938 26411 -4928
rect 17297 -5108 17373 -5098
rect 25868 -5108 25944 -5098
rect 17293 -5179 17297 -5113
rect 17373 -5179 17377 -5113
rect 17297 -5194 17373 -5184
rect 25868 -5194 25944 -5184
rect 25636 -5591 26033 -5581
rect 25636 -5657 26033 -5647
rect 26339 -5749 26411 -5010
rect 25636 -5759 26411 -5749
rect 26033 -5811 26411 -5759
rect 25636 -5821 26411 -5811
rect 17307 -6099 17363 -6089
rect 17307 -6165 17363 -6155
rect 8829 -6257 9226 -6247
rect 8829 -6319 9226 -6309
rect 25636 -6589 26033 -6579
rect 26555 -6589 26607 -2343
rect 26778 -2544 26830 -2534
rect 26772 -2596 26778 -2544
rect 26830 -2596 26836 -2544
rect 26033 -6641 26607 -6589
rect 25636 -6651 26033 -6641
rect 25636 -6755 26033 -6745
rect 26778 -6755 26830 -2596
rect 25634 -6807 25636 -6755
rect 26033 -6807 26830 -6755
rect 25636 -6817 26033 -6807
<< via2 >>
rect 9036 1490 9092 1546
rect 9416 -2760 9472 -2704
rect 17302 -5179 17368 -5113
rect 25868 -5184 25944 -5118
rect 25636 -5593 26033 -5591
rect 25636 -5645 26033 -5593
rect 25636 -5647 26033 -5645
rect 17307 -6155 17363 -6099
<< metal3 >>
rect 9031 1546 9097 1551
rect 9031 1490 9036 1546
rect 9092 1490 9097 1546
rect 9031 1485 9097 1490
rect 9396 -2700 9496 -2682
rect 9396 -2764 9412 -2700
rect 9476 -2764 9496 -2700
rect 9396 -2782 9496 -2764
rect 17297 -5113 17373 -5108
rect 17297 -5179 17302 -5113
rect 17368 -5179 17373 -5113
rect 17297 -6099 17373 -5179
rect 25858 -5118 25954 -5113
rect 25858 -5184 25868 -5118
rect 25944 -5184 25954 -5118
rect 25858 -5189 25954 -5184
rect 25868 -5586 25944 -5189
rect 25626 -5591 26043 -5586
rect 25626 -5647 25636 -5591
rect 26033 -5647 26043 -5591
rect 25626 -5652 26043 -5647
rect 17297 -6155 17307 -6099
rect 17363 -6155 17373 -6099
rect 17297 -6160 17373 -6155
<< via3 >>
rect 9412 -2704 9476 -2700
rect 9412 -2760 9416 -2704
rect 9416 -2760 9472 -2704
rect 9472 -2760 9476 -2704
rect 9412 -2764 9476 -2760
<< metal4 >>
rect 9411 -2700 9477 -2699
rect 9411 -2764 9412 -2700
rect 9476 -2764 9477 -2700
rect 9411 -3014 9477 -2764
use bjt  bjt_0
timestamp 1762795171
transform 1 0 -12427 0 1 -18123
box -53 -53 7324 6945
use digital  digital_0
timestamp 1720189102
transform 1 0 32771 0 1 -3754
box -397 -1200 2333 5008
use op5  op5_0
timestamp 1762786734
transform 1 0 9786 0 1 -6121
box -9786 6121 9272 13721
use pmos_current_bgr  pmos_current_bgr_0
timestamp 1762753955
transform 1 0 425 0 1 -1186
box -227 -676 8487 506
use res_trim  res_trim_0
timestamp 1720030020
transform 0 1 101 -1 0 -2857
box -31 -51 1533 15873
use resist_const  resist_const_0
timestamp 1720269525
transform -1 0 28465 0 -1 -9225
box 2257 -3964 28483 -2103
<< end >>
