magic
tech sky130A
magscale 1 2
timestamp 1717259999
<< error_p >>
rect -29 161 29 167
rect -29 127 -17 161
rect -29 121 29 127
<< nmos >>
rect -15 -151 15 89
<< ndiff >>
rect -73 77 -15 89
rect -73 -139 -61 77
rect -27 -139 -15 77
rect -73 -151 -15 -139
rect 15 77 73 89
rect 15 -139 27 77
rect 61 -139 73 77
rect 15 -151 73 -139
<< ndiffc >>
rect -61 -139 -27 77
rect 27 -139 61 77
<< poly >>
rect -33 161 33 177
rect -33 127 -17 161
rect 17 127 33 161
rect -33 111 33 127
rect -15 89 15 111
rect -15 -177 15 -151
<< polycont >>
rect -17 127 17 161
<< locali >>
rect -33 127 -17 161
rect 17 127 33 161
rect -61 77 -27 93
rect -61 -155 -27 -139
rect 27 77 61 93
rect 27 -155 61 -139
<< viali >>
rect -17 127 17 161
rect -61 -139 -27 77
rect 27 -139 61 77
<< metal1 >>
rect -29 161 29 167
rect -29 127 -17 161
rect 17 127 29 161
rect -29 121 29 127
rect -67 77 -21 89
rect -67 -139 -61 77
rect -27 -139 -21 77
rect -67 -151 -21 -139
rect 21 77 67 89
rect 21 -139 27 77
rect 61 -139 67 77
rect 21 -151 67 -139
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.2 l 0.150 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
