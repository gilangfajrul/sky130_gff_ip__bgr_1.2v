magic
tech sky130A
magscale 1 2
timestamp 1717913952
<< nmoslvt >>
rect -229 -431 -29 369
rect 29 -431 229 369
<< ndiff >>
rect -287 357 -229 369
rect -287 -419 -275 357
rect -241 -419 -229 357
rect -287 -431 -229 -419
rect -29 357 29 369
rect -29 -419 -17 357
rect 17 -419 29 357
rect -29 -431 29 -419
rect 229 357 287 369
rect 229 -419 241 357
rect 275 -419 287 357
rect 229 -431 287 -419
<< ndiffc >>
rect -275 -419 -241 357
rect -17 -419 17 357
rect 241 -419 275 357
<< poly >>
rect -229 441 -29 457
rect -229 407 -213 441
rect -45 407 -29 441
rect -229 369 -29 407
rect 29 441 229 457
rect 29 407 45 441
rect 213 407 229 441
rect 29 369 229 407
rect -229 -457 -29 -431
rect 29 -457 229 -431
<< polycont >>
rect -213 407 -45 441
rect 45 407 213 441
<< locali >>
rect -229 407 -213 441
rect -45 407 -29 441
rect 29 407 45 441
rect 213 407 229 441
rect -275 357 -241 373
rect -275 -435 -241 -419
rect -17 357 17 373
rect -17 -435 17 -419
rect 241 357 275 373
rect 241 -435 275 -419
<< viali >>
rect -213 407 -45 441
rect 45 407 213 441
rect -275 -419 -241 357
rect -17 -419 17 357
rect 241 -419 275 357
<< metal1 >>
rect -225 441 -33 447
rect -225 407 -213 441
rect -45 407 -33 441
rect -225 401 -33 407
rect 33 441 225 447
rect 33 407 45 441
rect 213 407 225 441
rect 33 401 225 407
rect -281 357 -235 369
rect -281 -419 -275 357
rect -241 -419 -235 357
rect -281 -431 -235 -419
rect -23 357 23 369
rect -23 -419 -17 357
rect 17 -419 23 357
rect -23 -431 23 -419
rect 235 357 281 369
rect 235 -419 241 357
rect 275 -419 281 357
rect 235 -431 281 -419
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 4 l 1 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
