magic
tech sky130A
magscale 1 2
timestamp 1716351939
<< error_p >>
rect -654 552 -516 554
rect -420 552 -282 554
rect -186 552 -48 554
rect 48 552 186 554
rect 282 552 420 554
rect 516 552 654 554
rect -654 -484 -516 -482
rect -420 -484 -282 -482
rect -186 -484 -48 -482
rect 48 -484 186 -482
rect 282 -484 420 -482
rect 516 -484 654 -482
<< nwell >>
rect -847 -1159 847 1159
<< nsubdiff >>
rect -811 1089 -715 1123
rect 715 1089 811 1123
rect -811 1027 -777 1089
rect 777 1027 811 1089
rect -811 -1089 -777 -1027
rect 777 -1089 811 -1027
rect -811 -1123 -715 -1089
rect 715 -1123 811 -1089
<< nsubdiffcont >>
rect -715 1089 715 1123
rect -811 -1027 -777 1027
rect 777 -1027 811 1027
rect -715 -1123 715 -1089
<< xpolycontact >>
rect -654 552 -516 984
rect -654 52 -516 484
rect -420 552 -282 984
rect -420 52 -282 484
rect -186 552 -48 984
rect -186 52 -48 484
rect 48 552 186 984
rect 48 52 186 484
rect 282 552 420 984
rect 282 52 420 484
rect 516 552 654 984
rect 516 52 654 484
rect -654 -484 -516 -52
rect -654 -984 -516 -552
rect -420 -484 -282 -52
rect -420 -984 -282 -552
rect -186 -484 -48 -52
rect -186 -984 -48 -552
rect 48 -484 186 -52
rect 48 -984 186 -552
rect 282 -484 420 -52
rect 282 -984 420 -552
rect 516 -484 654 -52
rect 516 -984 654 -552
<< ppolyres >>
rect -654 484 -516 552
rect -420 484 -282 552
rect -186 484 -48 552
rect 48 484 186 552
rect 282 484 420 552
rect 516 484 654 552
rect -654 -552 -516 -484
rect -420 -552 -282 -484
rect -186 -552 -48 -484
rect 48 -552 186 -484
rect 282 -552 420 -484
rect 516 -552 654 -484
<< locali >>
rect -811 1089 -715 1123
rect 715 1089 811 1123
rect -811 1027 -777 1089
rect 777 1027 811 1089
rect -811 -1089 -777 -1027
rect 777 -1089 811 -1027
rect -811 -1123 -715 -1089
rect 715 -1123 811 -1089
<< viali >>
rect -638 569 -532 966
rect -404 569 -298 966
rect -170 569 -64 966
rect 64 569 170 966
rect 298 569 404 966
rect 532 569 638 966
rect -638 70 -532 467
rect -404 70 -298 467
rect -170 70 -64 467
rect 64 70 170 467
rect 298 70 404 467
rect 532 70 638 467
rect -638 -467 -532 -70
rect -404 -467 -298 -70
rect -170 -467 -64 -70
rect 64 -467 170 -70
rect 298 -467 404 -70
rect 532 -467 638 -70
rect -638 -966 -532 -569
rect -404 -966 -298 -569
rect -170 -966 -64 -569
rect 64 -966 170 -569
rect 298 -966 404 -569
rect 532 -966 638 -569
<< metal1 >>
rect -644 966 -526 978
rect -644 569 -638 966
rect -532 569 -526 966
rect -644 557 -526 569
rect -410 966 -292 978
rect -410 569 -404 966
rect -298 569 -292 966
rect -410 557 -292 569
rect -176 966 -58 978
rect -176 569 -170 966
rect -64 569 -58 966
rect -176 557 -58 569
rect 58 966 176 978
rect 58 569 64 966
rect 170 569 176 966
rect 58 557 176 569
rect 292 966 410 978
rect 292 569 298 966
rect 404 569 410 966
rect 292 557 410 569
rect 526 966 644 978
rect 526 569 532 966
rect 638 569 644 966
rect 526 557 644 569
rect -644 467 -526 479
rect -644 70 -638 467
rect -532 70 -526 467
rect -644 58 -526 70
rect -410 467 -292 479
rect -410 70 -404 467
rect -298 70 -292 467
rect -410 58 -292 70
rect -176 467 -58 479
rect -176 70 -170 467
rect -64 70 -58 467
rect -176 58 -58 70
rect 58 467 176 479
rect 58 70 64 467
rect 170 70 176 467
rect 58 58 176 70
rect 292 467 410 479
rect 292 70 298 467
rect 404 70 410 467
rect 292 58 410 70
rect 526 467 644 479
rect 526 70 532 467
rect 638 70 644 467
rect 526 58 644 70
rect -644 -70 -526 -58
rect -644 -467 -638 -70
rect -532 -467 -526 -70
rect -644 -479 -526 -467
rect -410 -70 -292 -58
rect -410 -467 -404 -70
rect -298 -467 -292 -70
rect -410 -479 -292 -467
rect -176 -70 -58 -58
rect -176 -467 -170 -70
rect -64 -467 -58 -70
rect -176 -479 -58 -467
rect 58 -70 176 -58
rect 58 -467 64 -70
rect 170 -467 176 -70
rect 58 -479 176 -467
rect 292 -70 410 -58
rect 292 -467 298 -70
rect 404 -467 410 -70
rect 292 -479 410 -467
rect 526 -70 644 -58
rect 526 -467 532 -70
rect 638 -467 644 -70
rect 526 -479 644 -467
rect -644 -569 -526 -557
rect -644 -966 -638 -569
rect -532 -966 -526 -569
rect -644 -978 -526 -966
rect -410 -569 -292 -557
rect -410 -966 -404 -569
rect -298 -966 -292 -569
rect -410 -978 -292 -966
rect -176 -569 -58 -557
rect -176 -966 -170 -569
rect -64 -966 -58 -569
rect -176 -978 -58 -966
rect 58 -569 176 -557
rect 58 -966 64 -569
rect 170 -966 176 -569
rect 58 -978 176 -966
rect 292 -569 410 -557
rect 292 -966 298 -569
rect 404 -966 410 -569
rect 292 -978 410 -966
rect 526 -569 644 -557
rect 526 -966 532 -569
rect 638 -966 644 -569
rect 526 -978 644 -966
<< properties >>
string FIXED_BBOX -794 -1106 794 1106
string gencell sky130_fd_pr__res_high_po_0p69
string library sky130
string parameters w 0.690 l 0.50 m 2 nx 6 wmin 0.690 lmin 0.50 rho 319.8 val 796.434 dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.690 n_guard 1 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
