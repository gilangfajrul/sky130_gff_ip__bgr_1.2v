magic
tech sky130A
magscale 1 2
timestamp 1718385342
<< psubdiff >>
rect -176 410 -116 444
rect 690 410 750 444
rect -176 384 -142 410
rect 716 384 750 410
rect -176 -34 -142 -8
rect 716 -34 750 -8
rect -176 -68 -116 -34
rect 690 -68 750 -34
<< psubdiffcont >>
rect -116 410 690 444
rect -176 -8 -142 384
rect 716 -8 750 384
rect -116 -68 690 -34
<< poly >>
rect -92 360 0 376
rect -92 326 -76 360
rect -42 326 0 360
rect -92 310 0 326
rect -30 288 0 310
rect 574 50 666 66
rect 574 16 616 50
rect 650 16 666 50
rect 574 0 666 16
<< polycont >>
rect -76 326 -42 360
rect 616 16 650 50
<< locali >>
rect -176 410 -116 444
rect 690 410 750 444
rect -176 384 -142 410
rect 716 384 750 410
rect -76 360 -42 376
rect -76 288 -42 326
rect 616 50 650 99
rect 616 0 650 16
rect -176 -34 -142 -8
rect 716 -34 750 -8
rect -176 -68 -116 -34
rect 690 -68 750 -34
<< viali >>
rect -176 326 -142 360
rect -76 326 -42 360
rect 616 16 650 50
rect 716 16 750 50
<< metal1 >>
rect -182 360 -36 372
rect -182 326 -176 360
rect -142 326 -76 360
rect -42 326 -36 360
rect -182 314 -36 326
rect 254 320 320 366
rect -82 288 -36 314
rect 264 266 310 288
rect 6 52 52 90
rect 522 52 568 95
rect 6 6 568 52
rect 610 62 656 97
rect 610 50 756 62
rect 610 16 616 50
rect 650 16 716 50
rect 750 16 756 50
rect 610 4 756 16
use sky130_fd_pr__nfet_01v8_lvt_SJFSNB  sky130_fd_pr__nfet_01v8_lvt_SJFSNB_1
timestamp 1717911345
transform 1 0 -15 0 1 188
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_lvt_SJFSNB  sky130_fd_pr__nfet_01v8_lvt_SJFSNB_2
timestamp 1717911345
transform 1 0 589 0 1 188
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_lvt_U8VHVM  sky130_fd_pr__nfet_01v8_lvt_U8VHVM_0
timestamp 1717912059
transform 1 0 287 0 1 219
box -287 -157 287 157
<< labels >>
flabel metal1 284 354 284 354 0 FreeSans 160 0 0 0 G
port 0 nsew
flabel metal1 282 32 282 32 0 FreeSans 160 0 0 0 D
port 1 nsew
flabel metal1 288 280 288 280 0 FreeSans 160 0 0 0 S
port 2 nsew
flabel metal1 702 30 702 30 0 FreeSans 160 0 0 0 DVSS
port 3 nsew
<< end >>
