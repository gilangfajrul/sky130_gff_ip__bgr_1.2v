magic
tech sky130A
magscale 1 2
timestamp 1762795171
<< dnwell >>
rect -53 -53 6945 6945
<< locali >>
rect 6108 5760 6142 5794
rect 1481 5644 1482 5741
rect 2869 5644 2870 5741
rect 4257 5644 4258 5741
rect 5645 5644 5646 5741
rect 1151 5409 1247 5412
rect 1151 4021 1247 4024
rect 1151 2633 1247 2636
rect 1481 1151 1482 1245
rect 2635 1151 2646 1238
rect 4257 1151 4258 1245
rect 5645 1154 5646 1231
<< viali >>
rect 1079 5741 1151 5813
rect 1215 5741 1314 5813
rect 1414 5741 1513 5813
rect 1577 5741 1649 5813
rect 2467 5741 2539 5813
rect 2603 5741 2702 5813
rect 2802 5741 2901 5813
rect 2965 5741 3037 5813
rect 3855 5741 3927 5813
rect 3991 5741 4090 5813
rect 4190 5741 4289 5813
rect 4353 5741 4425 5813
rect 5243 5741 5315 5813
rect 5379 5741 5478 5813
rect 5578 5741 5677 5813
rect 5741 5741 5813 5813
rect 1079 5578 1151 5677
rect 5741 5578 5813 5677
rect 1079 5379 1151 5478
rect 1079 5243 1151 5315
rect 1079 4353 1151 4425
rect 2467 4353 2539 4425
rect 2603 4353 2702 4425
rect 2802 4353 2901 4425
rect 2965 4353 3037 4425
rect 3855 4353 3927 4425
rect 3991 4353 4090 4425
rect 4190 4353 4289 4425
rect 4353 4353 4425 4425
rect 5741 4353 5813 4425
rect 1079 4190 1151 4289
rect 2467 4190 2539 4289
rect 4353 4190 4425 4289
rect 5741 4190 5813 4289
rect 1079 3991 1151 4090
rect 2467 3991 2539 4090
rect 2965 3991 3037 4090
rect 3855 3991 3927 4090
rect 4353 3991 4425 4090
rect 5741 3991 5813 4090
rect 1079 3855 1151 3927
rect 2467 3855 2539 3927
rect 2802 3855 2901 3927
rect 2965 3855 3037 3927
rect 3855 3855 3927 3927
rect 3991 3855 4090 3927
rect 4353 3855 4425 3927
rect 5741 3855 5813 3927
rect 1079 2965 1151 3037
rect 2467 2965 2539 3037
rect 2802 2965 2901 3037
rect 2965 2965 3037 3037
rect 3855 2965 3927 3037
rect 3991 2965 4090 3037
rect 4353 2965 4425 3037
rect 5741 2965 5813 3037
rect 1079 2802 1151 2901
rect 2467 2802 2539 2901
rect 2965 2802 3037 2901
rect 3855 2802 3927 2901
rect 4353 2802 4425 2901
rect 5741 2802 5813 2901
rect 1079 2603 1151 2702
rect 2467 2603 2539 2702
rect 4353 2603 4425 2702
rect 5741 2603 5813 2702
rect 1079 2467 1151 2539
rect 2467 2467 2539 2539
rect 2603 2467 2702 2539
rect 2802 2467 2901 2539
rect 2965 2467 3037 2539
rect 3855 2467 3927 2539
rect 3991 2467 4090 2539
rect 4190 2467 4289 2539
rect 4353 2467 4425 2539
rect 5741 2467 5813 2539
rect 1079 1577 1151 1649
rect 5741 1577 5813 1649
rect 1079 1414 1151 1513
rect 5741 1414 5813 1513
rect 1079 1216 1151 1315
rect 1079 1080 1151 1152
rect 1215 1080 1314 1152
rect 5741 1215 5813 1314
rect 1414 1079 1513 1151
rect 1577 1079 1649 1151
rect 2467 1079 2539 1151
rect 2603 1079 2702 1151
rect 2802 1079 2901 1151
rect 2965 1079 3037 1151
rect 3855 1079 3927 1151
rect 3991 1079 4090 1151
rect 4190 1079 4289 1151
rect 4353 1079 4425 1151
rect 5243 1079 5315 1151
rect 5379 1079 5478 1151
rect 5578 1079 5677 1151
rect 5741 1079 5813 1151
<< metal1 >>
rect 876 6372 6232 6528
rect 364 5552 520 5988
rect 1340 5826 1388 6372
rect 2728 5826 2776 6372
rect 4116 5826 4164 6372
rect 5504 5826 5552 6372
rect 1066 5813 5826 5826
rect 1066 5741 1079 5813
rect 1151 5741 1215 5813
rect 1314 5741 1414 5813
rect 1513 5741 1577 5813
rect 1649 5741 2467 5813
rect 2539 5741 2603 5813
rect 2702 5780 2802 5813
rect 2702 5741 2726 5780
rect 1066 5728 2726 5741
rect 2778 5741 2802 5780
rect 2901 5741 2965 5813
rect 3037 5741 3855 5813
rect 3927 5741 3991 5813
rect 4090 5780 4190 5813
rect 4090 5741 4114 5780
rect 2778 5728 4114 5741
rect 4166 5741 4190 5780
rect 4289 5741 4353 5813
rect 4425 5741 5243 5813
rect 5315 5741 5379 5813
rect 5478 5741 5578 5813
rect 5677 5741 5741 5813
rect 5813 5741 5826 5813
rect 4166 5728 5826 5741
rect 1066 5677 1164 5728
rect 1066 5578 1079 5677
rect 1151 5578 1164 5677
rect 1066 5552 1164 5578
rect 364 5504 1164 5552
rect 364 4164 520 5504
rect 1066 5478 1164 5504
rect 1066 5379 1079 5478
rect 1151 5379 1164 5478
rect 1066 5315 1164 5379
rect 1066 5243 1079 5315
rect 1151 5243 1164 5315
rect 1066 4425 1164 5243
rect 5728 5677 5826 5728
rect 5728 5578 5741 5677
rect 5813 5578 5826 5677
rect 5728 5552 5826 5578
rect 6371 5552 6527 6028
rect 5728 5504 6527 5552
rect 1066 4353 1079 4425
rect 1151 4353 1164 4425
rect 1066 4289 1164 4353
rect 1066 4190 1079 4289
rect 1151 4190 1164 4289
rect 1066 4164 1164 4190
rect 364 4116 1164 4164
rect 364 2776 520 4116
rect 1066 4090 1164 4116
rect 1066 3991 1079 4090
rect 1151 3991 1164 4090
rect 1066 3927 1164 3991
rect 1066 3855 1079 3927
rect 1151 3855 1164 3927
rect 1066 3037 1164 3855
rect 1066 2965 1079 3037
rect 1151 2965 1164 3037
rect 1066 2901 1164 2965
rect 1066 2802 1079 2901
rect 1151 2802 1164 2901
rect 1066 2776 1164 2802
rect 364 2728 1164 2776
rect 364 1388 520 2728
rect 1066 2702 1164 2728
rect 1066 2603 1079 2702
rect 1151 2603 1164 2702
rect 1066 2539 1164 2603
rect 1066 2467 1079 2539
rect 1151 2467 1164 2539
rect 1066 1649 1164 2467
rect 1753 5007 5139 5139
rect 1753 1885 1885 5007
rect 2455 4425 2726 4437
rect 2455 4353 2467 4425
rect 2539 4353 2603 4425
rect 2702 4385 2726 4425
rect 2778 4425 4114 4437
rect 2778 4385 2802 4425
rect 2702 4353 2802 4385
rect 2901 4353 2965 4425
rect 3037 4353 3855 4425
rect 3927 4353 3991 4425
rect 4090 4385 4114 4425
rect 4166 4425 4437 4437
rect 4166 4385 4190 4425
rect 4090 4353 4190 4385
rect 4289 4353 4353 4425
rect 4425 4353 4437 4425
rect 2455 4341 4437 4353
rect 2455 4289 2551 4341
rect 2455 4190 2467 4289
rect 2539 4190 2551 4289
rect 2455 4090 2551 4190
rect 4341 4289 4437 4341
rect 4341 4190 4353 4289
rect 4425 4190 4437 4289
rect 2455 3991 2467 4090
rect 2539 3991 2551 4090
rect 2455 3932 2551 3991
rect 2959 4090 3043 4102
rect 2959 3991 2965 4090
rect 3037 3991 3043 4090
rect 2959 3933 3043 3991
rect 3849 4090 3933 4102
rect 3849 3991 3855 4090
rect 3927 3991 3933 4090
rect 3849 3933 3933 3991
rect 4341 4090 4437 4190
rect 4341 3991 4353 4090
rect 4425 3991 4437 4090
rect 4341 3933 4437 3991
rect 2790 3932 4437 3933
rect 2455 3927 4437 3932
rect 2455 3855 2467 3927
rect 2539 3855 2802 3927
rect 2901 3855 2965 3927
rect 3037 3855 3855 3927
rect 3927 3855 3991 3927
rect 4090 3855 4353 3927
rect 4425 3855 4437 3927
rect 2455 3849 4437 3855
rect 2455 3848 2895 3849
rect 2455 3043 2551 3848
rect 2959 3043 3043 3849
rect 3320 3402 3330 3506
rect 3578 3402 3588 3506
rect 3849 3043 3933 3849
rect 4341 3043 4437 3849
rect 2455 3037 4437 3043
rect 2455 2965 2467 3037
rect 2539 2965 2802 3037
rect 2901 2965 2965 3037
rect 3037 2965 3855 3037
rect 3927 2965 3991 3037
rect 4090 2965 4353 3037
rect 4425 2965 4437 3037
rect 2455 2959 4437 2965
rect 2455 2901 2551 2959
rect 2455 2802 2467 2901
rect 2539 2802 2551 2901
rect 2455 2702 2551 2802
rect 2959 2901 3043 2959
rect 2959 2802 2965 2901
rect 3037 2802 3043 2901
rect 2959 2790 3043 2802
rect 3849 2901 3933 2959
rect 3849 2802 3855 2901
rect 3927 2802 3933 2901
rect 3849 2790 3933 2802
rect 4341 2901 4437 2959
rect 4341 2802 4353 2901
rect 4425 2802 4437 2901
rect 2455 2603 2467 2702
rect 2539 2603 2551 2702
rect 2455 2551 2551 2603
rect 4341 2702 4437 2802
rect 4341 2603 4353 2702
rect 4425 2603 4437 2702
rect 4341 2551 4437 2603
rect 2455 2539 4437 2551
rect 2455 2467 2467 2539
rect 2539 2467 2603 2539
rect 2702 2507 2802 2539
rect 2702 2467 2726 2507
rect 2455 2455 2726 2467
rect 2778 2467 2802 2507
rect 2901 2467 2965 2539
rect 3037 2467 3855 2539
rect 3927 2467 3991 2539
rect 4090 2507 4190 2539
rect 4090 2467 4114 2507
rect 2778 2455 4114 2467
rect 4166 2467 4190 2507
rect 4289 2467 4353 2539
rect 4425 2467 4437 2539
rect 4166 2455 4437 2467
rect 5007 1885 5139 5007
rect 1753 1753 5139 1885
rect 5728 4425 5826 5504
rect 5728 4353 5741 4425
rect 5813 4353 5826 4425
rect 5728 4289 5826 4353
rect 5728 4190 5741 4289
rect 5813 4190 5826 4289
rect 5728 4164 5826 4190
rect 6371 4164 6527 5504
rect 5728 4116 6527 4164
rect 5728 4090 5826 4116
rect 5728 3991 5741 4090
rect 5813 3991 5826 4090
rect 5728 3927 5826 3991
rect 5728 3855 5741 3927
rect 5813 3855 5826 3927
rect 5728 3037 5826 3855
rect 5728 2965 5741 3037
rect 5813 2965 5826 3037
rect 5728 2901 5826 2965
rect 5728 2802 5741 2901
rect 5813 2802 5826 2901
rect 5728 2776 5826 2802
rect 6371 2776 6527 4116
rect 5728 2728 6527 2776
rect 5728 2702 5826 2728
rect 5728 2603 5741 2702
rect 5813 2603 5826 2702
rect 5728 2539 5826 2603
rect 5728 2467 5741 2539
rect 5813 2467 5826 2539
rect 1066 1577 1079 1649
rect 1151 1577 1164 1649
rect 1066 1513 1164 1577
rect 1066 1414 1079 1513
rect 1151 1414 1164 1513
rect 1066 1388 1164 1414
rect 364 1340 1164 1388
rect 364 629 520 1340
rect 1066 1315 1164 1340
rect 1066 1216 1079 1315
rect 1151 1216 1164 1315
rect 1066 1165 1164 1216
rect 5728 1649 5826 2467
rect 5728 1577 5741 1649
rect 5813 1577 5826 1649
rect 5728 1513 5826 1577
rect 5728 1414 5741 1513
rect 5813 1414 5826 1513
rect 5728 1388 5826 1414
rect 6371 1388 6527 2728
rect 5728 1340 6527 1388
rect 5728 1314 5826 1340
rect 5728 1215 5741 1314
rect 5813 1215 5826 1314
rect 5728 1165 5826 1215
rect 1066 1152 2726 1165
rect 1066 1080 1079 1152
rect 1151 1080 1215 1152
rect 1314 1151 2726 1152
rect 1314 1080 1414 1151
rect 1066 1079 1414 1080
rect 1513 1079 1577 1151
rect 1649 1079 2467 1151
rect 2539 1079 2603 1151
rect 2702 1113 2726 1151
rect 2778 1151 4114 1165
rect 2778 1113 2802 1151
rect 2702 1079 2802 1113
rect 2901 1079 2965 1151
rect 3037 1079 3855 1151
rect 3927 1079 3991 1151
rect 4090 1113 4114 1151
rect 4166 1151 5826 1165
rect 4166 1113 4190 1151
rect 4090 1079 4190 1113
rect 4289 1079 4353 1151
rect 4425 1079 5243 1151
rect 5315 1079 5379 1151
rect 5478 1079 5578 1151
rect 5677 1079 5741 1151
rect 5813 1079 5826 1151
rect 1066 1067 5826 1079
rect 1340 520 1388 1067
rect 2728 520 2776 1067
rect 4116 520 4164 1067
rect 5504 520 5552 1067
rect 6371 672 6527 1340
rect 877 364 6233 520
<< via1 >>
rect 2726 5728 2778 5780
rect 4114 5728 4166 5780
rect 2726 4385 2778 4437
rect 4114 4385 4166 4437
rect 3330 3402 3578 3506
rect 2726 2455 2778 2507
rect 4114 2455 4166 2507
rect 2726 1113 2778 1165
rect 4114 1113 4166 1165
<< metal2 >>
rect 2726 5780 2778 5790
rect 2726 4437 2778 5728
rect 2726 4375 2778 4385
rect 4114 5780 4166 5790
rect 4114 4437 4166 5728
rect 4114 4375 4166 4385
rect 3330 3506 7324 3516
rect 3578 3402 7324 3506
rect 3330 3392 7324 3402
rect 2726 2507 2778 2517
rect 2726 1165 2778 2455
rect 2726 1103 2778 1113
rect 4114 2507 4166 2517
rect 4114 1165 4166 2455
rect 4114 1103 4166 1113
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
array 0 4 1388 0 4 1388
timestamp 1759091000
transform 1 0 0 0 1 0
box 0 0 1340 1340
<< labels >>
flabel metal2 7097 3423 7097 3423 0 FreeSans 1600 0 0 0 A
port 14 nsew
flabel metal1 5064 4136 5064 4136 0 FreeSans 1600 0 0 0 B
port 9 nsew
flabel metal1 5785 2755 5785 2755 0 FreeSans 1600 0 0 0 AVSS
port 5 nsew
<< end >>
