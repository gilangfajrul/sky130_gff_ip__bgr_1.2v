magic
tech sky130A
magscale 1 2
timestamp 1762707440
<< nwell >>
rect 0 0 8362 836
<< metal1 >>
rect 2087 548 2097 724
rect 2149 548 2159 724
rect 6203 548 6213 724
rect 6265 548 6275 724
rect 29 112 39 288
rect 91 112 101 288
rect 2087 112 2097 288
rect 2149 112 2159 288
rect 6203 112 6213 288
rect 6265 112 6275 288
<< via1 >>
rect 2097 548 2149 724
rect 6213 548 6265 724
rect 39 112 91 288
rect 2097 112 2149 288
rect 6213 112 6265 288
<< metal2 >>
rect 2097 724 2149 734
rect 39 288 91 298
rect 39 102 91 112
rect 2097 288 2149 548
rect 2097 102 2149 112
rect 6213 724 6265 734
rect 6213 288 6265 548
rect 6213 102 6265 112
use sky130_fd_pr__pfet_01v8_NDVM6J  sky130_fd_pr__pfet_01v8_NDVM6J_0
timestamp 1762707440
transform 1 0 4181 0 1 418
box -4181 -418 4181 418
<< end >>
