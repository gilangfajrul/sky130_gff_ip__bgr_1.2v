magic
tech sky130A
magscale 1 2
timestamp 1762704772
<< error_p >>
rect -2123 18 2123 236
<< nwell >>
rect -2123 18 2123 418
rect -2123 -418 2123 -18
<< pmos >>
rect -2029 118 -29 318
rect 29 118 2029 318
rect -2029 -318 -29 -118
rect 29 -318 2029 -118
<< pdiff >>
rect -2087 306 -2029 318
rect -2087 130 -2075 306
rect -2041 130 -2029 306
rect -2087 118 -2029 130
rect -29 306 29 318
rect -29 130 -17 306
rect 17 130 29 306
rect -29 118 29 130
rect 2029 306 2087 318
rect 2029 130 2041 306
rect 2075 130 2087 306
rect 2029 118 2087 130
rect -2087 -130 -2029 -118
rect -2087 -306 -2075 -130
rect -2041 -306 -2029 -130
rect -2087 -318 -2029 -306
rect -29 -130 29 -118
rect -29 -306 -17 -130
rect 17 -306 29 -130
rect -29 -318 29 -306
rect 2029 -130 2087 -118
rect 2029 -306 2041 -130
rect 2075 -306 2087 -130
rect 2029 -318 2087 -306
<< pdiffc >>
rect -2075 130 -2041 306
rect -17 130 17 306
rect 2041 130 2075 306
rect -2075 -306 -2041 -130
rect -17 -306 17 -130
rect 2041 -306 2075 -130
<< poly >>
rect -2029 399 -29 415
rect -2029 365 -2013 399
rect -45 365 -29 399
rect -2029 318 -29 365
rect 29 399 2029 415
rect 29 365 45 399
rect 2013 365 2029 399
rect 29 318 2029 365
rect -2029 71 -29 118
rect -2029 37 -2013 71
rect -45 37 -29 71
rect -2029 21 -29 37
rect 29 71 2029 118
rect 29 37 45 71
rect 2013 37 2029 71
rect 29 21 2029 37
rect -2029 -37 -29 -21
rect -2029 -71 -2013 -37
rect -45 -71 -29 -37
rect -2029 -118 -29 -71
rect 29 -37 2029 -21
rect 29 -71 45 -37
rect 2013 -71 2029 -37
rect 29 -118 2029 -71
rect -2029 -365 -29 -318
rect -2029 -399 -2013 -365
rect -45 -399 -29 -365
rect -2029 -415 -29 -399
rect 29 -365 2029 -318
rect 29 -399 45 -365
rect 2013 -399 2029 -365
rect 29 -415 2029 -399
<< polycont >>
rect -2013 365 -45 399
rect 45 365 2013 399
rect -2013 37 -45 71
rect 45 37 2013 71
rect -2013 -71 -45 -37
rect 45 -71 2013 -37
rect -2013 -399 -45 -365
rect 45 -399 2013 -365
<< locali >>
rect -2029 365 -2013 399
rect -45 365 -29 399
rect 29 365 45 399
rect 2013 365 2029 399
rect -2075 306 -2041 322
rect -2075 114 -2041 130
rect -17 306 17 322
rect -17 114 17 130
rect 2041 306 2075 322
rect 2041 114 2075 130
rect -2029 37 -2013 71
rect -45 37 -29 71
rect 29 37 45 71
rect 2013 37 2029 71
rect -2029 -71 -2013 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 2013 -71 2029 -37
rect -2075 -130 -2041 -114
rect -2075 -322 -2041 -306
rect -17 -130 17 -114
rect -17 -322 17 -306
rect 2041 -130 2075 -114
rect 2041 -322 2075 -306
rect -2029 -399 -2013 -365
rect -45 -399 -29 -365
rect 29 -399 45 -365
rect 2013 -399 2029 -365
<< viali >>
rect -2013 365 -45 399
rect 45 365 2013 399
rect -2075 130 -2041 306
rect -17 130 17 306
rect 2041 130 2075 306
rect -2013 37 -45 71
rect 45 37 2013 71
rect -2013 -71 -45 -37
rect 45 -71 2013 -37
rect -2075 -306 -2041 -130
rect -17 -306 17 -130
rect 2041 -306 2075 -130
rect -2013 -399 -45 -365
rect 45 -399 2013 -365
<< metal1 >>
rect -2025 399 -33 405
rect -2025 365 -2013 399
rect -45 365 -33 399
rect -2025 359 -33 365
rect 33 399 2025 405
rect 33 365 45 399
rect 2013 365 2025 399
rect 33 359 2025 365
rect -2081 306 -2035 318
rect -2081 130 -2075 306
rect -2041 130 -2035 306
rect -2081 118 -2035 130
rect -23 306 23 318
rect -23 130 -17 306
rect 17 130 23 306
rect -23 118 23 130
rect 2035 306 2081 318
rect 2035 130 2041 306
rect 2075 130 2081 306
rect 2035 118 2081 130
rect -2025 71 -33 77
rect -2025 37 -2013 71
rect -45 37 -33 71
rect -2025 31 -33 37
rect 33 71 2025 77
rect 33 37 45 71
rect 2013 37 2025 71
rect 33 31 2025 37
rect -2025 -37 -33 -31
rect -2025 -71 -2013 -37
rect -45 -71 -33 -37
rect -2025 -77 -33 -71
rect 33 -37 2025 -31
rect 33 -71 45 -37
rect 2013 -71 2025 -37
rect 33 -77 2025 -71
rect -2081 -130 -2035 -118
rect -2081 -306 -2075 -130
rect -2041 -306 -2035 -130
rect -2081 -318 -2035 -306
rect -23 -130 23 -118
rect -23 -306 -17 -130
rect 17 -306 23 -130
rect -23 -318 23 -306
rect 2035 -130 2081 -118
rect 2035 -306 2041 -130
rect 2075 -306 2081 -130
rect 2035 -318 2081 -306
rect -2025 -365 -33 -359
rect -2025 -399 -2013 -365
rect -45 -399 -33 -365
rect -2025 -405 -33 -399
rect 33 -365 2025 -359
rect 33 -399 45 -365
rect 2013 -399 2025 -365
rect 33 -405 2025 -399
<< labels >>
rlabel pdiffc -2058 -218 -2058 -218 0 D0_0
port 1 nsew
rlabel polycont -1029 -54 -1029 -54 0 G0_0
port 2 nsew
rlabel pdiffc -2058 218 -2058 218 0 D0_1
port 3 nsew
rlabel polycont -1029 382 -1029 382 0 G0_1
port 4 nsew
rlabel pdiffc 0 -218 0 -218 0 S1_0
port 5 nsew
rlabel polycont 1029 -54 1029 -54 0 G1_0
port 6 nsew
rlabel pdiffc 0 218 0 218 0 S1_1
port 7 nsew
rlabel polycont 1029 382 1029 382 0 G1_1
port 8 nsew
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 10 m 2 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 conn_gates 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 doports 1
<< end >>
