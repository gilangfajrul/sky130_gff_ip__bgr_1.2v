magic
tech sky130A
magscale 1 2
timestamp 1720425981
<< dnwell >>
rect -17914 13826 9178 22978
rect -17914 226 -1066 13826
rect 8559 226 9178 13826
rect -17914 -412 9178 226
<< nwell >>
rect -17994 22772 9258 23058
rect -17994 -206 -17708 22772
rect -16736 14678 -2960 17678
rect -16736 14626 -3776 14678
rect 8972 -206 9258 22772
rect -17994 -492 9258 -206
<< pwell >>
rect -17561 20831 8723 22741
rect -413 20788 8402 20831
rect 8584 17910 8723 18355
rect -1328 17868 8723 17910
rect 8584 17858 8723 17868
rect -1328 14640 8723 17858
<< nsubdiff >>
rect -17957 23001 9221 23021
rect -17957 22967 -17877 23001
rect 9141 22967 9221 23001
rect -17957 22947 9221 22967
rect -17957 22941 -17883 22947
rect -17957 -375 -17937 22941
rect -17903 -375 -17883 22941
rect -17957 -381 -17883 -375
rect 9147 22941 9221 22947
rect 9147 -375 9167 22941
rect 9201 -375 9221 22941
rect 9147 -381 9221 -375
rect -17957 -401 9221 -381
rect -17957 -435 -17877 -401
rect 9141 -435 9221 -401
rect -17957 -455 9221 -435
<< nsubdiffcont >>
rect -17877 22967 9141 23001
rect -17937 -375 -17903 22941
rect 9167 -375 9201 22941
rect -17877 -435 9141 -401
<< locali >>
rect -17937 22967 -17877 23001
rect 9141 22967 9201 23001
rect -17937 22941 -17903 22967
rect 9167 22941 9201 22967
rect -17937 -401 -17903 -375
rect 9167 -401 9201 -375
rect -17937 -435 -17877 -401
rect 9141 -435 9201 -401
<< viali >>
rect 604 10291 638 10471
rect 757 9973 937 10007
<< metal1 >>
rect -17365 22325 -17355 22395
rect -16923 22325 -16913 22395
rect -17365 22159 -17355 22229
rect -16923 22159 -16913 22229
rect 342 22002 352 22054
rect 404 22002 414 22054
rect -540 21836 -530 21888
rect -133 21836 -123 21888
rect 4678 21836 4688 21888
rect 4740 21836 4750 21888
rect -17074 21338 -17064 21390
rect -16940 21338 -16930 21390
rect -17336 21162 -17326 21234
rect -17254 21162 -17244 21234
rect -17402 20218 -16759 20880
rect -13038 20772 -12065 20878
rect -13013 20441 -12955 20732
rect -17412 20077 -17402 20218
rect -16759 20077 -16749 20218
rect -13011 19608 -13001 19660
rect -12604 19608 -12594 19660
rect -7744 18369 -7734 18435
rect -7668 18369 -6604 18435
rect -2178 17409 -2044 17928
rect -2188 17275 -2178 17409
rect -2044 17275 -2034 17409
rect -16527 16799 -16517 16975
rect -16395 16799 -16385 16975
rect -988 16861 -978 16913
rect -894 16861 -884 16913
rect -8030 16391 -7978 16397
rect -8030 16333 -7978 16339
rect -3302 16282 -3292 16458
rect -3240 16282 -3230 16458
rect -102 16094 -92 16270
rect -40 16094 -30 16270
rect 856 15845 1662 15948
rect 2709 15821 4264 15885
rect 4328 15821 4338 15885
rect -12144 15579 -11338 15682
rect -11736 15462 -11726 15514
rect -10742 15462 -10732 15514
rect -9678 15462 -9668 15514
rect -8684 15462 -8674 15514
rect -7949 15494 -7540 15685
rect -6595 15563 -5789 15666
rect -12387 15101 -12377 15153
rect -12325 15101 -12315 15153
rect -7847 14457 -7631 15494
rect -7472 15301 -7462 15477
rect -7410 15301 -7400 15477
rect -3189 15351 -3179 15423
rect -3127 15351 -3117 15423
rect -1198 15341 -862 15391
rect -1198 15225 -1120 15341
rect 2063 15340 2073 15392
rect 2193 15340 2203 15392
rect 2709 15310 2773 15821
rect 4659 15762 5632 15940
rect 8369 15650 8379 15710
rect 8439 15650 8449 15710
rect 3795 15575 3805 15627
rect 5089 15575 5099 15627
rect 6453 15573 6463 15629
rect 7747 15573 7757 15629
rect 2709 15240 2773 15246
rect -1198 15175 -863 15225
rect 2063 15174 2073 15226
rect 2193 15174 2203 15226
rect -3190 14882 -3180 14942
rect -3128 14882 -3118 14942
rect -7847 14456 5584 14457
rect -7847 14240 5594 14456
rect 773 11390 783 12166
rect 835 11390 845 12166
rect 4418 11812 4428 11864
rect 4604 11812 4614 11864
rect 5378 11791 5594 14240
rect 4989 11707 5983 11791
rect 4418 11466 4428 11518
rect 4604 11466 4614 11518
rect 4635 11255 4645 11307
rect 4697 11255 4707 11307
rect 6025 10917 9119 10966
rect 4418 10698 4428 10750
rect 4604 10698 4614 10750
rect 594 10471 647 10483
rect 594 10291 604 10471
rect 638 10291 647 10471
rect 4418 10352 4428 10404
rect 4604 10352 4614 10404
rect 594 9818 647 10291
rect 745 10007 949 10013
rect 745 9973 757 10007
rect 937 9973 949 10007
rect 745 9967 949 9973
rect 1041 9979 1093 10351
rect 1933 10059 1985 10347
rect 2825 10139 2877 10348
rect 3717 10219 3769 10346
rect 3717 10167 9119 10219
rect 2825 10087 9119 10139
rect 1933 10007 9119 10059
rect 821 9899 874 9967
rect 1041 9927 9119 9979
rect 821 9846 9119 9899
rect 594 9765 9119 9818
rect 2225 6234 2235 6500
rect 2501 6234 2511 6500
rect 658 1904 668 2515
rect 1278 1904 1288 2515
<< via1 >>
rect -17355 22325 -16923 22395
rect -17355 22159 -16923 22229
rect 352 22002 404 22054
rect -530 21836 -133 21888
rect 4688 21836 4740 21888
rect -17064 21338 -16940 21390
rect -17326 21162 -17254 21234
rect -17402 20077 -16759 20218
rect -13001 19608 -12604 19660
rect -7734 18369 -7668 18435
rect -2178 17275 -2044 17409
rect -16517 16799 -16395 16975
rect -978 16861 -894 16913
rect -8030 16339 -7978 16391
rect -3292 16282 -3240 16458
rect -92 16094 -40 16270
rect 4264 15821 4328 15885
rect -11726 15462 -10742 15514
rect -9668 15462 -8684 15514
rect -12377 15101 -12325 15153
rect -7462 15301 -7410 15477
rect -3179 15351 -3127 15423
rect 2073 15340 2193 15392
rect 8379 15650 8439 15710
rect 3805 15575 5089 15627
rect 6463 15573 7747 15629
rect 2709 15246 2773 15310
rect 2073 15174 2193 15226
rect -3180 14882 -3128 14942
rect 783 11390 835 12166
rect 4428 11812 4604 11864
rect 4428 11466 4604 11518
rect 4645 11255 4697 11307
rect 4428 10698 4604 10750
rect 4428 10352 4604 10404
rect 2235 6234 2501 6500
rect 668 1904 1278 2515
<< metal2 >>
rect -17355 22404 -16923 22405
rect -17610 22395 -16923 22404
rect -17610 22394 -17355 22395
rect -17611 22325 -17355 22394
rect -17611 22315 -16923 22325
rect -17611 22314 -17268 22315
rect -17611 20658 -17487 22314
rect -17355 22229 -16923 22239
rect -17355 22149 -16923 22159
rect 352 22054 404 22064
rect -530 21888 -133 21898
rect -530 21826 -133 21836
rect -8684 21733 -8675 21805
rect -8603 21733 -8594 21805
rect -8675 21670 -8603 21733
rect -17064 21390 -16940 21400
rect -17326 21234 -17254 21244
rect -17326 21152 -17254 21162
rect -17064 20811 -16940 21338
rect -17064 20697 -17059 20811
rect -16945 20697 -16940 20811
rect -364 20808 -298 21826
rect 352 21154 404 22002
rect 4688 21888 4740 21898
rect 348 21145 408 21154
rect 348 21076 408 21085
rect 4688 20938 4740 21836
rect 4675 20878 4684 20938
rect 4744 20878 4753 20938
rect -364 20752 -359 20808
rect -303 20752 -298 20808
rect -364 20747 -298 20752
rect -359 20743 -303 20747
rect -17064 20692 -16940 20697
rect -17059 20688 -16945 20692
rect -17611 20534 -16542 20658
rect -17402 20218 -16759 20228
rect -17402 20067 -16759 20077
rect -16666 17149 -16542 20534
rect -13001 19660 -12604 19670
rect -13001 19598 -12604 19608
rect -12694 18926 -12634 19598
rect -8763 19438 -8703 19447
rect -8763 19260 -8703 19378
rect -8763 19200 -7242 19260
rect -7626 19128 -7502 19138
rect -7378 19004 -7369 19128
rect -7626 18994 -7502 19004
rect -7878 18926 -7822 18933
rect -12694 18924 -7820 18926
rect -12694 18868 -7878 18924
rect -7822 18868 -7820 18924
rect -12694 18866 -7820 18868
rect -7878 18859 -7822 18866
rect -7734 18435 -7668 18445
rect -7734 18359 -7668 18369
rect -7502 17594 -7378 18880
rect -7302 17711 -7242 19200
rect -159 17711 -103 17719
rect -7302 17709 -101 17711
rect -7302 17653 -159 17709
rect -103 17653 -94 17709
rect -7302 17651 -101 17653
rect -159 17643 -103 17651
rect -1777 17594 -1549 17599
rect -7502 17589 -1544 17594
rect -7502 17475 -1777 17589
rect -1549 17475 -1540 17589
rect -7502 17470 -1663 17475
rect -1777 17465 -1663 17470
rect -2178 17409 -2044 17419
rect -2182 17280 -2178 17404
rect -2044 17280 -2040 17404
rect -1549 17470 -1544 17475
rect -1663 17351 -1549 17361
rect -2178 17265 -2044 17275
rect -2842 17233 -2770 17242
rect -2770 17161 -967 17233
rect -2842 17152 -2770 17161
rect -16666 17025 -16394 17149
rect -16518 16975 -16394 17025
rect -16518 16800 -16517 16975
rect -16395 16800 -16394 16975
rect -12324 16974 -12268 16985
rect -16517 16789 -16395 16799
rect -1120 16857 -1111 16917
rect -1051 16913 -1042 16917
rect -978 16913 -894 16923
rect -1051 16861 -978 16913
rect -1051 16857 -1042 16861
rect -12324 16789 -12268 16799
rect -3281 16855 -1364 16857
rect -3281 16799 -1422 16855
rect -1366 16799 -1357 16855
rect -978 16851 -894 16861
rect -1281 16803 -1221 16812
rect -3281 16797 -1364 16799
rect -1281 16734 -1221 16743
rect 41 16664 97 16674
rect -3123 16582 -136 16628
rect 41 16478 97 16488
rect -3292 16458 -3240 16468
rect -8036 16339 -8030 16391
rect -7978 16339 -7398 16391
rect -2426 16453 -2366 16462
rect -1109 16453 -1053 16460
rect -2366 16451 -1051 16453
rect -2366 16395 -1109 16451
rect -1053 16395 -1051 16451
rect -2366 16393 -1051 16395
rect -2426 16384 -2366 16393
rect -1109 16386 -1053 16393
rect -3128 16312 -3072 16319
rect -3292 16173 -3240 16282
rect -3130 16310 -40 16312
rect -3130 16254 -3128 16310
rect -3072 16270 -40 16310
rect -3072 16254 -92 16270
rect -3130 16252 -92 16254
rect -3128 16245 -3072 16252
rect -3292 16121 -236 16173
rect -288 15929 -236 16121
rect -92 16084 -40 16094
rect -161 16034 -101 16044
rect 6458 16030 6467 16034
rect -101 15978 6467 16030
rect 6458 15974 6467 15978
rect 6527 15974 6536 16034
rect -161 15964 -101 15974
rect 3079 15929 3088 15933
rect -1971 15916 -1875 15926
rect -375 15916 -319 15917
rect -2977 15856 -2968 15916
rect -2908 15856 -1971 15916
rect -2977 15849 -1971 15856
rect -1875 15914 -318 15916
rect -1875 15858 -1279 15914
rect -1223 15909 -318 15914
rect -1223 15907 -317 15909
rect -1223 15858 -375 15907
rect -1875 15851 -375 15858
rect -319 15851 -317 15907
rect -288 15877 3088 15929
rect 3079 15873 3088 15877
rect 3148 15873 3157 15933
rect 4264 15885 4328 15895
rect -1875 15849 -317 15851
rect -1971 15839 -1875 15849
rect -375 15841 -319 15849
rect 4259 15825 4264 15881
rect 4328 15825 4333 15881
rect 4264 15811 4328 15821
rect -10820 15658 -10742 15798
rect -9668 15658 -9590 15800
rect -1668 15791 -1544 15801
rect -1544 15737 3857 15789
rect -1668 15725 -1544 15735
rect -10820 15656 -2908 15658
rect -10820 15600 -2966 15656
rect -2910 15600 -2901 15656
rect -1424 15653 -1364 15663
rect 2888 15653 2944 15661
rect -10820 15598 -2908 15600
rect -10820 15524 -10742 15598
rect -11726 15514 -10742 15524
rect -11726 15452 -10742 15462
rect -9668 15524 -9590 15598
rect 2879 15651 2944 15653
rect 2879 15649 2888 15651
rect -1364 15597 2888 15649
rect -1424 15583 -1364 15593
rect -9668 15514 -8684 15524
rect -9668 15452 -8684 15462
rect -7889 15431 -7880 15491
rect -7820 15487 -7811 15491
rect -7820 15477 -7410 15487
rect -7820 15435 -7462 15477
rect -7820 15431 -7811 15435
rect -3179 15423 -3127 15433
rect -3127 15418 -2770 15423
rect -3127 15356 -2837 15418
rect -2775 15356 -2766 15418
rect -2675 15413 -1322 15418
rect -2679 15357 -2670 15413
rect -2614 15357 -1322 15413
rect -3127 15351 -2770 15356
rect -2675 15352 -1322 15357
rect -1256 15352 -1247 15418
rect 2073 15392 2193 15597
rect 2879 15595 2888 15597
rect 2944 15595 2953 15651
rect 3805 15637 3857 15737
rect 8379 15710 8439 15720
rect 8372 15652 8379 15708
rect 8439 15652 8446 15708
rect 6463 15639 6532 15649
rect 8379 15640 8439 15650
rect 3805 15627 5089 15637
rect 2888 15585 2944 15595
rect 3805 15565 5089 15575
rect 6532 15629 7747 15639
rect 6532 15563 7747 15573
rect 6463 15553 6532 15563
rect -3179 15341 -3127 15351
rect -7462 15291 -7410 15301
rect 2073 15226 2193 15340
rect 2531 15246 2709 15310
rect 2773 15246 2779 15310
rect 2073 15164 2193 15174
rect -12377 15153 -12325 15163
rect -17788 15101 -12377 15153
rect 2886 15115 2946 15125
rect -12377 15091 -12325 15101
rect -1155 15079 -1065 15088
rect -1065 15008 -898 15060
rect 2877 15055 2886 15115
rect 2946 15111 2955 15115
rect 2946 15059 3147 15111
rect 2946 15055 2955 15059
rect 2886 15045 2946 15055
rect -1155 14980 -1065 14989
rect -3180 14942 -3128 14952
rect -3128 14940 -2366 14942
rect -3128 14884 -2424 14940
rect -2368 14884 -2359 14940
rect -3128 14882 -2366 14884
rect -3180 14872 -3128 14882
rect -2187 14813 -2178 14947
rect -2044 14942 -582 14947
rect -2044 14818 -711 14942
rect -587 14818 -578 14942
rect -2044 14813 -582 14818
rect -1668 14715 -1544 14725
rect -7743 14573 -7734 14639
rect -7668 14573 -1739 14639
rect -1805 14306 -1739 14573
rect -1544 14591 -1420 14601
rect -913 14591 -799 14596
rect -1420 14586 -794 14591
rect -1420 14467 -913 14586
rect -1668 14457 -1420 14467
rect -799 14467 -794 14586
rect 776 14582 842 14587
rect 772 14526 781 14582
rect 837 14526 846 14582
rect -913 14348 -799 14358
rect -266 14306 -210 14310
rect -1805 14301 -205 14306
rect -1805 14245 -266 14301
rect -210 14245 -205 14301
rect -1805 14240 -205 14245
rect -266 14236 -210 14240
rect -1322 14020 -415 14025
rect -1326 13964 -1317 14020
rect -1261 13964 -415 14020
rect -1322 13959 -415 13964
rect -349 13959 -340 14025
rect 776 12166 842 14526
rect 4724 14430 4784 14439
rect 4724 14361 4784 14370
rect 2817 14306 2884 14316
rect 4326 14275 4382 14282
rect 2817 14230 2884 14240
rect 4324 14273 4384 14275
rect 1926 14175 1992 14184
rect 1034 14020 1100 14025
rect 1030 13964 1039 14020
rect 1095 13964 1104 14020
rect 776 11390 783 12166
rect 835 11390 842 12166
rect 776 11380 842 11390
rect 1034 10386 1100 13964
rect 1926 10388 1992 14109
rect 2817 10386 2883 14230
rect 4324 14217 4326 14273
rect 4382 14217 4384 14273
rect 4324 10750 4384 14217
rect 4428 11864 4604 11874
rect 4728 11864 4780 14361
rect 4604 11812 4780 11864
rect 4428 11802 4604 11812
rect 4428 11518 4604 11528
rect 4604 11466 4863 11518
rect 4428 11456 4604 11466
rect 4645 11307 4697 11317
rect 4697 11255 4783 11307
rect 4645 11245 4697 11255
rect 4428 10750 4604 10760
rect 4324 10698 4428 10750
rect 4428 10688 4604 10698
rect 4731 10495 4783 11255
rect 4811 10589 4863 11466
rect 4991 11076 9119 11422
rect 4811 10537 9119 10589
rect 4731 10443 9119 10495
rect -1158 9162 -1062 9171
rect -1715 9068 -1629 9072
rect -1720 9066 -1158 9068
rect 3717 9123 3769 10408
rect 4428 10404 4604 10414
rect 4604 10352 9119 10404
rect 4428 10342 4604 10352
rect -1720 9063 -1062 9066
rect -1720 8977 -1715 9063
rect -1629 8977 -1062 9063
rect -1720 8972 -1062 8977
rect -918 8988 -794 8998
rect -725 8989 -716 9123
rect -582 9118 3769 9123
rect -582 8994 2291 9118
rect 2415 8994 3769 9118
rect -582 8989 3769 8994
rect -1715 8968 -1629 8972
rect -794 8864 -670 8874
rect -927 8740 -918 8864
rect -670 8740 3803 8864
rect -918 8730 -670 8740
rect 2235 6500 2501 6510
rect 2235 6224 2501 6234
rect 668 2515 1278 2525
rect 668 1894 1278 1904
<< via2 >>
rect -17355 22159 -16923 22229
rect -8675 21733 -8603 21805
rect -17321 21167 -17259 21229
rect -17059 20697 -16945 20811
rect 348 21085 408 21145
rect 4684 20878 4744 20938
rect -359 20752 -303 20808
rect -17402 20077 -16759 20218
rect -8763 19378 -8703 19438
rect -7626 19004 -7378 19128
rect -7878 18868 -7822 18924
rect -7502 18880 -7378 19004
rect -7734 18369 -7668 18435
rect -159 17653 -103 17709
rect -1777 17475 -1549 17589
rect -2173 17280 -2049 17404
rect -1663 17361 -1549 17475
rect -2842 17161 -2770 17233
rect -12324 16799 -12268 16974
rect -1111 16857 -1051 16917
rect -1422 16799 -1366 16855
rect -1281 16743 -1221 16803
rect 41 16488 97 16664
rect -2426 16393 -2366 16453
rect -1109 16395 -1053 16451
rect -3128 16254 -3072 16310
rect -161 15974 -101 16034
rect 6467 15974 6527 16034
rect -2968 15856 -2908 15916
rect -1971 15849 -1875 15916
rect -1279 15858 -1223 15914
rect -375 15851 -319 15907
rect 3088 15873 3148 15933
rect 4264 15821 4328 15885
rect -1668 15735 -1544 15791
rect -2966 15600 -2910 15656
rect -1424 15593 -1364 15653
rect -7880 15431 -7820 15491
rect -2837 15356 -2775 15418
rect -2670 15357 -2614 15413
rect -1322 15352 -1256 15418
rect 2888 15595 2944 15651
rect 8381 15652 8437 15708
rect 6463 15629 6532 15639
rect 6463 15573 6532 15629
rect 6463 15563 6532 15573
rect -1155 14989 -1065 15079
rect 2886 15055 2946 15115
rect -2424 14884 -2368 14940
rect -2178 14813 -2044 14947
rect -711 14818 -587 14942
rect -7734 14573 -7668 14639
rect -1668 14591 -1544 14715
rect -1668 14467 -1420 14591
rect -913 14358 -799 14586
rect 781 14526 837 14582
rect -266 14245 -210 14301
rect -1317 13964 -1261 14020
rect -415 13959 -349 14025
rect 4724 14370 4784 14430
rect 2817 14240 2884 14306
rect 1926 14109 1992 14175
rect 1039 13964 1095 14020
rect 4326 14217 4382 14273
rect -1158 9066 -1062 9162
rect -1715 8977 -1629 9063
rect -716 8989 -582 9123
rect 2291 8994 2415 9118
rect -918 8864 -794 8988
rect -918 8740 -670 8864
rect 2235 6234 2501 6500
rect 668 1904 1278 2515
<< metal3 >>
rect -17365 22232 -16913 22234
rect -17617 22229 -16913 22232
rect -17617 22159 -17355 22229
rect -16923 22159 -16913 22229
rect -17617 22156 -16913 22159
rect -17617 20629 -17541 22156
rect -17365 22154 -16913 22156
rect -8680 21805 -8598 21810
rect -17481 21733 -8675 21805
rect -8603 21733 -8598 21805
rect -17481 21234 -17409 21733
rect -8763 21668 -8598 21733
rect -17481 21229 -17254 21234
rect -17481 21167 -17321 21229
rect -17259 21167 -17254 21229
rect -17481 21162 -17254 21167
rect -17064 20811 -13191 20816
rect -17064 20697 -17059 20811
rect -16945 20697 -13191 20811
rect -17064 20692 -13191 20697
rect -17617 20553 -13377 20629
rect -17412 20218 -16749 20223
rect -17412 20077 -17402 20218
rect -16759 20077 -16749 20218
rect -17412 20072 -16749 20077
rect -13453 18920 -13377 20553
rect -13315 19128 -13191 20692
rect -8763 19443 -8703 21668
rect 343 21145 413 21150
rect 8570 21147 8634 21153
rect 343 21085 348 21145
rect 408 21085 8570 21145
rect 343 21080 413 21085
rect 8570 21077 8634 21083
rect 4679 20938 4749 20943
rect 8427 20938 8433 20940
rect 4679 20878 4684 20938
rect 4744 20878 8433 20938
rect 4679 20873 4749 20878
rect 8427 20876 8433 20878
rect 8497 20876 8503 20940
rect 8309 20813 8373 20818
rect -364 20812 8374 20813
rect -364 20808 8309 20812
rect -364 20752 -359 20808
rect -303 20752 8309 20808
rect -364 20748 8309 20752
rect 8373 20748 8374 20812
rect -364 20747 8374 20748
rect 8309 20742 8373 20747
rect -8768 19438 -8698 19443
rect -8768 19378 -8763 19438
rect -8703 19378 -8698 19438
rect -8768 19373 -8698 19378
rect -7636 19128 -7368 19133
rect -13315 19004 -7626 19128
rect -7636 18999 -7502 19004
rect -7883 18924 -7817 18929
rect -13453 18844 -12258 18920
rect -7883 18868 -7878 18924
rect -7822 18868 -7817 18924
rect -7512 18880 -7502 18999
rect -7378 18880 -7368 19128
rect -7512 18875 -7368 18880
rect -7883 18863 -7817 18868
rect -12334 16974 -12258 18844
rect -12334 16799 -12324 16974
rect -12268 16799 -12258 16974
rect -12334 16794 -12258 16799
rect -7880 15496 -7820 18863
rect -7744 18435 -7658 18440
rect -7744 18369 -7734 18435
rect -7668 18369 -7658 18435
rect -7744 18364 -7658 18369
rect -7885 15491 -7815 15496
rect -7885 15431 -7880 15491
rect -7820 15431 -7815 15491
rect -7885 15426 -7815 15431
rect -7734 14644 -7668 18364
rect -2674 17640 -2610 17645
rect -2675 17639 -2609 17640
rect -2675 17575 -2674 17639
rect -2610 17575 -2609 17639
rect -2847 17233 -2765 17238
rect -2847 17161 -2842 17233
rect -2770 17161 -2765 17233
rect -2847 17156 -2765 17161
rect -3133 16310 -3067 16315
rect -3133 16254 -3128 16310
rect -3072 16254 -3067 16310
rect -3133 16249 -3067 16254
rect -2973 15916 -2903 15921
rect -2973 15856 -2968 15916
rect -2908 15856 -2903 15916
rect -2973 15851 -2903 15856
rect -2968 15661 -2908 15851
rect -2971 15656 -2905 15661
rect -2971 15600 -2966 15656
rect -2910 15600 -2905 15656
rect -2971 15595 -2905 15600
rect -2842 15418 -2770 17156
rect -2842 15356 -2837 15418
rect -2775 15356 -2770 15418
rect -2842 15351 -2770 15356
rect -2675 15413 -2609 17575
rect -1787 17589 -1539 17594
rect -1787 17475 -1777 17589
rect -1787 17470 -1663 17475
rect -2178 17404 -2044 17409
rect -2178 17280 -2173 17404
rect -2049 17280 -2044 17404
rect -1673 17361 -1663 17470
rect -1549 17361 -1539 17589
rect -1673 17356 -1539 17361
rect -2431 16453 -2361 16458
rect -2431 16393 -2426 16453
rect -2366 16393 -2361 16453
rect -2431 16388 -2361 16393
rect -2675 15357 -2670 15413
rect -2614 15357 -2609 15413
rect -2675 15352 -2609 15357
rect -2426 14945 -2366 16388
rect -2178 14952 -2044 17280
rect -1981 15916 -1865 15921
rect -1981 15849 -1971 15916
rect -1875 15849 -1865 15916
rect -1981 15844 -1865 15849
rect -1971 15205 -1875 15844
rect -1668 15796 -1544 17356
rect -1116 16917 -1046 16922
rect -1427 16855 -1361 16860
rect -1427 16799 -1422 16855
rect -1366 16799 -1361 16855
rect -1116 16857 -1111 16917
rect -1051 16857 -1046 16917
rect -1116 16852 -1046 16857
rect -1427 16794 -1361 16799
rect -1286 16803 -1216 16808
rect -1678 15791 -1534 15796
rect -1678 15735 -1668 15791
rect -1544 15735 -1534 15791
rect -1678 15730 -1534 15735
rect -1980 15111 -1970 15205
rect -1876 15111 -1866 15205
rect -1971 15110 -1875 15111
rect -2183 14947 -2039 14952
rect -2429 14940 -2363 14945
rect -2429 14884 -2424 14940
rect -2368 14884 -2363 14940
rect -2429 14879 -2363 14884
rect -2183 14813 -2178 14947
rect -2044 14813 -2039 14947
rect -2183 14808 -2039 14813
rect -1668 14720 -1544 15730
rect -1424 15658 -1364 16794
rect -1286 16743 -1281 16803
rect -1221 16743 -1216 16803
rect -1286 16738 -1216 16743
rect -1281 15919 -1221 16738
rect -1111 16456 -1051 16852
rect -1114 16451 -1048 16456
rect -1114 16395 -1109 16451
rect -1053 16395 -1048 16451
rect -1114 16390 -1048 16395
rect -1284 15914 -1218 15919
rect -1284 15858 -1279 15914
rect -1223 15858 -1218 15914
rect -1284 15853 -1218 15858
rect -1434 15653 -1354 15658
rect -1434 15593 -1424 15653
rect -1364 15593 -1354 15653
rect -1434 15588 -1354 15593
rect -1327 15418 -1251 15423
rect -1327 15352 -1322 15418
rect -1256 15352 -1251 15418
rect -1327 15347 -1251 15352
rect -1678 14715 -1534 14720
rect -7739 14639 -7663 14644
rect -7739 14573 -7734 14639
rect -7668 14573 -7663 14639
rect -7739 14568 -7663 14573
rect -1678 14467 -1668 14715
rect -1544 14596 -1534 14715
rect -1544 14591 -1410 14596
rect -1420 14467 -1410 14591
rect -1678 14462 -1410 14467
rect -1322 14020 -1256 15347
rect -1160 15079 -1060 15084
rect -1160 14989 -1155 15079
rect -1065 14989 -1060 15079
rect -1160 14984 -1060 14989
rect -1322 13964 -1317 14020
rect -1261 13964 -1256 14020
rect -1322 13959 -1256 13964
rect -1158 9167 -1062 14984
rect -716 14942 -582 14947
rect -716 14818 -711 14942
rect -587 14818 -582 14942
rect -923 14586 -789 14591
rect -923 14358 -913 14586
rect -799 14358 -789 14586
rect -923 14353 -789 14358
rect -1163 9162 -1057 9167
rect -1719 9068 -1625 9073
rect -1720 9067 -1624 9068
rect -1720 8973 -1719 9067
rect -1625 8973 -1624 9067
rect -1163 9066 -1158 9162
rect -1062 9066 -1057 9162
rect -1163 9061 -1057 9066
rect -918 8993 -794 14353
rect -716 9128 -582 14818
rect -511 14175 -445 17819
rect -169 17709 -93 17714
rect -169 17653 -159 17709
rect -103 17653 -93 17709
rect -169 17648 -93 17653
rect -161 16039 -101 17648
rect 31 16664 107 16669
rect 31 16488 41 16664
rect 97 16488 107 16664
rect 31 16483 107 16488
rect -171 16034 -91 16039
rect -171 15974 -161 16034
rect -101 15974 -91 16034
rect -171 15969 -91 15974
rect -385 15909 -309 15912
rect 39 15909 99 16483
rect -385 15907 99 15909
rect -385 15851 -375 15907
rect -319 15851 99 15907
rect 3083 15933 3153 15938
rect 3083 15873 3088 15933
rect 3148 15873 3153 15933
rect 4264 15890 4328 16144
rect 6462 16034 6532 16039
rect 6462 15974 6467 16034
rect 6527 15974 6532 16034
rect 3083 15868 3153 15873
rect 4254 15885 4338 15890
rect -385 15849 99 15851
rect -385 15846 -309 15849
rect 2878 15651 2954 15656
rect 2878 15595 2888 15651
rect 2944 15595 2954 15651
rect 2878 15590 2954 15595
rect 2886 15120 2946 15590
rect 3088 15418 3148 15868
rect 4254 15821 4264 15885
rect 4328 15821 4338 15885
rect 4254 15816 4338 15821
rect 6462 15644 6532 15974
rect 8379 15713 8439 16734
rect 8376 15708 8442 15713
rect 8376 15652 8381 15708
rect 8437 15652 8442 15708
rect 8376 15647 8442 15652
rect 6453 15639 6542 15644
rect 6453 15563 6463 15639
rect 6532 15563 6542 15639
rect 6453 15558 6542 15563
rect 2876 15115 2956 15120
rect 2876 15055 2886 15115
rect 2946 15055 2956 15115
rect 2876 15050 2956 15055
rect 776 14586 8593 14587
rect 776 14582 8528 14586
rect 776 14526 781 14582
rect 837 14526 8528 14582
rect 776 14522 8528 14526
rect 8592 14522 8598 14586
rect 776 14521 8593 14522
rect 4719 14430 4789 14435
rect 8646 14430 8652 14432
rect 4719 14370 4724 14430
rect 4784 14370 8652 14430
rect 4719 14365 4789 14370
rect 8646 14368 8652 14370
rect 8716 14368 8722 14432
rect 2807 14306 2894 14311
rect -271 14301 2817 14306
rect -271 14245 -266 14301
rect -210 14245 2817 14301
rect -271 14240 2817 14245
rect 2884 14240 2894 14306
rect 2807 14235 2894 14240
rect 4321 14275 4387 14278
rect 8769 14275 8775 14277
rect 4321 14273 8775 14275
rect 4321 14217 4326 14273
rect 4382 14217 8775 14273
rect 4321 14215 8775 14217
rect 4321 14212 4387 14215
rect 8769 14213 8775 14215
rect 8839 14213 8845 14277
rect 1921 14175 1997 14180
rect -511 14109 1926 14175
rect 1992 14109 1997 14175
rect 1921 14104 1997 14109
rect -420 14025 -344 14030
rect -420 13959 -415 14025
rect -349 14020 1100 14025
rect -349 13964 1039 14020
rect 1095 13964 1100 14020
rect -349 13959 1100 13964
rect -420 13954 -344 13959
rect -721 9123 -577 9128
rect -1720 8972 -1624 8973
rect -928 8988 -784 8993
rect -1719 8967 -1625 8972
rect -928 8740 -918 8988
rect -794 8869 -784 8988
rect -721 8989 -716 9123
rect -582 8989 -577 9123
rect -721 8984 -577 8989
rect 2286 9118 2420 9123
rect 2286 8994 2291 9118
rect 2415 8994 2420 9118
rect -794 8864 -660 8869
rect -670 8740 -660 8864
rect -928 8735 -660 8740
rect 2286 7516 2420 8994
rect 2300 6505 2406 7516
rect 2225 6500 2511 6505
rect 2225 6234 2235 6500
rect 2501 6234 2511 6500
rect 2225 6229 2511 6234
rect 658 2515 1288 2520
rect 658 1904 668 2515
rect 1278 1904 1288 2515
rect 658 1899 1288 1904
<< via3 >>
rect -17402 20077 -16759 20218
rect 8570 21083 8634 21147
rect 8433 20876 8497 20940
rect 8309 20748 8373 20812
rect -2674 17575 -2610 17639
rect -1970 15111 -1876 15205
rect -1719 9063 -1625 9067
rect -1719 8977 -1715 9063
rect -1715 8977 -1629 9063
rect -1629 8977 -1625 9063
rect -1719 8973 -1625 8977
rect 8528 14522 8592 14586
rect 8652 14368 8716 14432
rect 8775 14213 8839 14277
rect 668 1904 1278 2515
<< metal4 >>
rect 8569 21147 8635 21148
rect 8569 21083 8570 21147
rect 8634 21083 8635 21147
rect 8569 21082 8635 21083
rect 8432 20940 8498 20941
rect 8432 20876 8433 20940
rect 8497 20876 8498 20940
rect 8432 20875 8498 20876
rect 8308 20812 8374 20813
rect 8308 20748 8309 20812
rect 8373 20748 8374 20812
rect -17403 20218 -16758 20219
rect -17403 20077 -17402 20218
rect -16759 20077 -16758 20218
rect -17403 20076 -16758 20077
rect -17402 13968 -16759 20076
rect -6977 19116 -4706 19182
rect -6977 17640 -6911 19116
rect 8308 17675 8374 20748
rect 8435 17808 8495 20875
rect 8572 17957 8632 21082
rect 8572 17897 8837 17957
rect 8435 17748 8714 17808
rect -6977 17639 -2609 17640
rect -6977 17575 -2674 17639
rect -2610 17575 -2609 17639
rect 8308 17609 8593 17675
rect -6977 17574 -2609 17575
rect -1971 15205 -1410 15206
rect -1971 15111 -1970 15205
rect -1876 15111 -1410 15205
rect -1971 15110 -1410 15111
rect -16227 13968 -15584 13970
rect -17402 13325 -15583 13968
rect -16227 1904 -15584 13325
rect -1857 9067 -1624 9068
rect -1857 8973 -1719 9067
rect -1625 8973 -1624 9067
rect -1857 8972 -1624 8973
rect -1506 7210 -1410 15110
rect 8527 14586 8593 17609
rect 8527 14522 8528 14586
rect 8592 14522 8593 14586
rect 8527 14521 8593 14522
rect 8654 14433 8714 17748
rect 8651 14432 8717 14433
rect 8651 14368 8652 14432
rect 8716 14368 8717 14432
rect 8651 14367 8717 14368
rect 8777 14278 8837 17897
rect 8774 14277 8840 14278
rect 8774 14213 8775 14277
rect 8839 14213 8840 14277
rect 8774 14212 8840 14213
rect -1790 7114 -1410 7210
rect 667 2515 1279 2516
rect 667 2487 668 2515
rect -2370 1904 668 2487
rect 1278 1904 1279 2515
rect -16227 1903 1279 1904
rect -16227 1873 1208 1903
rect -16227 1846 668 1873
rect -16227 1261 -1874 1846
rect -16227 163 -15584 1261
use bjt  bjt_0
timestamp 1720190288
transform 0 -1 7195 1 0 1540
box -53 -53 7324 6945
use cap_op  cap_op_0
timestamp 1718554435
transform 1 0 -5617 0 1 11002
box -12037 -11160 3906 3480
use differential_pair  differential_pair_0
timestamp 1720116957
transform 1 0 3459 0 1 14898
box -606 -124 5240 892
use digital  digital_0
timestamp 1720189102
transform 0 1 1450 -1 0 12249
box -397 -1200 2333 5008
use nmos_startup  nmos_startup_0
timestamp 1720119402
transform 1 0 -1078 0 1 16928
box -204 -154 746 692
use nmos_tail_current  nmos_tail_current_0
timestamp 1720118050
transform -1 0 8378 0 1 16054
box -321 -141 8599 1579
use pmos_current_bgr  pmos_current_bgr_0
timestamp 1720110902
transform 1 0 -16475 0 1 17121
box -260 -1493 8610 556
use pmos_current_bgr_2  pmos_current_bgr_2_0
timestamp 1720112176
transform -1 0 -3210 0 1 17072
box -250 -1450 4496 516
use pmos_iptat  pmos_iptat_0
timestamp 1720112315
transform 1 0 -12328 0 1 14730
box -191 -104 4438 898
use pmos_startup  pmos_startup_0
timestamp 1720267898
transform -1 0 -3176 0 1 15183
box -176 -494 4422 430
use res_trim  res_trim_0
timestamp 1720030020
transform 0 -1 8672 1 0 17734
box -31 -51 1533 15873
use resist_const  resist_const_0
timestamp 1720269525
transform 1 0 -19769 0 1 24804
box 2257 -3964 28483 -2103
use resistor_op_tt  resistor_op_tt_0
timestamp 1720284839
transform 0 -1 4860 1 0 15108
box -417 2220 767 6092
use resistorstart  resistorstart_0
timestamp 1718868641
transform 1 0 -13132 0 -1 20778
box -53 -53 21855 1511
<< labels >>
flabel metal4 -17203 19230 -17203 19230 0 FreeSans 1600 0 0 0 AVSS
port 2 nsew
flabel metal2 -16596 19440 -16596 19440 0 FreeSans 1600 0 0 0 VREF
port 3 nsew
flabel metal1 9111 9954 9111 9954 0 FreeSans 160 0 0 0 TRIM3
port 4 nsew
flabel metal1 9111 10033 9111 10033 0 FreeSans 160 0 0 0 TRIM2
port 5 nsew
flabel metal1 9111 10113 9111 10113 0 FreeSans 160 0 0 0 TRIM1
port 6 nsew
flabel metal1 9111 10193 9111 10193 0 FreeSans 160 0 0 0 TRIM0
port 7 nsew
flabel metal2 9111 10379 9111 10379 0 FreeSans 160 0 0 0 VBGSC
port 8 nsew
flabel metal2 9111 10471 9111 10471 0 FreeSans 160 0 0 0 VENA
port 9 nsew
flabel metal2 9111 10564 9111 10564 0 FreeSans 160 0 0 0 VBGTC
port 10 nsew
flabel metal1 9111 10941 9111 10941 0 FreeSans 160 0 0 0 ENA
port 11 nsew
flabel metal1 9110 9871 9110 9871 0 FreeSans 160 0 0 0 DVDD
port 13 nsew
flabel metal1 9110 9790 9110 9790 0 FreeSans 160 0 0 0 DVSS
port 14 nsew
flabel metal2 -17769 15128 -17769 15128 0 FreeSans 160 0 0 0 IPTAT
port 15 nsew
flabel metal2 9111 11252 9111 11252 0 FreeSans 160 0 0 0 AVDD
port 12 nsew
flabel metal1 -7792 15260 -7792 15260 0 FreeSans 160 0 0 0 VDDE
port 16 nsew
<< end >>
