magic
tech sky130A
magscale 1 2
timestamp 1764413320
<< dnwell >>
rect -5408 -8432 -2510 10622
rect -1012 -8432 27624 10622
rect 28904 -8432 37567 10622
<< nwell >>
rect -5488 10416 -2430 10702
rect -5488 -8226 -5202 10416
rect -2716 -8226 -2430 10416
rect -5488 -8512 -2430 -8226
rect -1092 10416 27704 10702
rect -1092 -8226 -806 10416
rect 27418 -8226 27704 10416
rect -1092 -8512 27704 -8226
rect 28824 10416 37647 10702
rect 28824 -8226 29110 10416
rect 37361 -8226 37647 10416
rect 28824 -8512 37647 -8226
<< pwell >>
rect 352 -3415 494 -3301
rect 8543 -4591 8902 -4356
<< psubdiff >>
rect 8661 -4441 8785 -4417
rect 8661 -4505 8686 -4441
rect 8761 -4505 8785 -4441
rect 8661 -4528 8785 -4505
<< nsubdiff >>
rect -5451 10645 -2467 10665
rect -5451 10611 -5371 10645
rect -2547 10611 -2467 10645
rect -5451 10591 -2467 10611
rect -5451 10585 -5377 10591
rect -5451 -8395 -5431 10585
rect -5397 -8395 -5377 10585
rect -5451 -8401 -5377 -8395
rect -2541 10585 -2467 10591
rect -2541 -8395 -2521 10585
rect -2487 -8395 -2467 10585
rect -2541 -8401 -2467 -8395
rect -5451 -8421 -2467 -8401
rect -5451 -8455 -5371 -8421
rect -2547 -8455 -2467 -8421
rect -5451 -8475 -2467 -8455
rect -1055 10645 27667 10665
rect -1055 10611 -975 10645
rect 27587 10611 27667 10645
rect -1055 10591 27667 10611
rect -1055 10585 -981 10591
rect -1055 -8395 -1035 10585
rect -1001 -8395 -981 10585
rect 27593 10585 27667 10591
rect -1055 -8401 -981 -8395
rect 27593 -8395 27613 10585
rect 27647 -8395 27667 10585
rect 27593 -8401 27667 -8395
rect -1055 -8421 27667 -8401
rect -1055 -8455 -975 -8421
rect 27587 -8455 27667 -8421
rect -1055 -8475 27667 -8455
rect 28861 10645 37610 10665
rect 28861 10611 28941 10645
rect 37530 10611 37610 10645
rect 28861 10591 37610 10611
rect 28861 10585 28935 10591
rect 28861 -8395 28881 10585
rect 28915 -8395 28935 10585
rect 28861 -8401 28935 -8395
rect 37536 10585 37610 10591
rect 37536 -8395 37556 10585
rect 37590 -8395 37610 10585
rect 37536 -8401 37610 -8395
rect 28861 -8421 37610 -8401
rect 28861 -8455 28941 -8421
rect 37530 -8455 37610 -8421
rect 28861 -8475 37610 -8455
<< psubdiffcont >>
rect 8686 -4505 8761 -4441
<< nsubdiffcont >>
rect -5371 10611 -2547 10645
rect -5431 -8395 -5397 10585
rect -2521 -8395 -2487 10585
rect -5371 -8455 -2547 -8421
rect -975 10611 27587 10645
rect -1035 -8395 -1001 10585
rect 27613 -8395 27647 10585
rect -975 -8455 27587 -8421
rect 28941 10611 37530 10645
rect 28881 -8395 28915 10585
rect 37556 -8395 37590 10585
rect 28941 -8455 37530 -8421
<< locali >>
rect -5431 10611 -5371 10645
rect -2547 10611 -2487 10645
rect -5431 10585 -5397 10611
rect -2521 10585 -2487 10611
rect -5431 -8421 -5397 -8395
rect -2521 -8421 -2487 -8395
rect -5431 -8455 -5371 -8421
rect -2547 -8455 -2487 -8421
rect -1035 10611 -975 10645
rect 27587 10611 27647 10645
rect -1035 10585 -1001 10611
rect 27613 10585 27647 10611
rect 8670 -4441 8776 -4425
rect 8670 -4505 8686 -4441
rect 8761 -4505 8776 -4441
rect 8670 -4521 8776 -4505
rect -1035 -8421 -1001 -8395
rect 27613 -8421 27647 -8395
rect -1035 -8455 -975 -8421
rect 27587 -8455 27647 -8421
rect 28881 10611 28941 10645
rect 37530 10611 37590 10645
rect 28881 10585 28915 10611
rect 28881 -8421 28915 -8395
rect 37556 10585 37590 10611
rect 37556 -8421 37590 -8395
rect 28881 -8455 28941 -8421
rect 37530 -8455 37590 -8421
<< viali >>
rect -4585 -798 -4551 -764
rect -4974 -1374 -4940 -1340
rect 8686 -4505 8761 -4441
<< metal1 >>
rect 16653 6636 16756 7080
rect 17848 6998 17858 7050
rect 17910 6998 17920 7050
rect 16653 6533 30380 6636
rect 17231 5947 17283 5953
rect 17283 5895 19463 5947
rect 19515 5895 19521 5947
rect 17231 5889 17283 5895
rect 17848 5716 17858 5768
rect 17910 5716 17920 5768
rect 19767 3249 19870 6533
rect 19020 3146 19870 3249
rect 19160 2845 19240 2851
rect 16812 2790 16822 2842
rect 18106 2790 18116 2842
rect 19240 2765 19450 2845
rect 19530 2765 19536 2845
rect 19160 2759 19240 2765
rect -5562 -1340 -4928 -1334
rect -5562 -1374 -4974 -1340
rect -4940 -1374 -4928 -1340
rect -4880 -1360 -4834 1230
rect -4253 327 -4243 379
rect -4059 327 -4049 379
rect -3413 -176 -3337 -170
rect -3413 -240 -3408 -176
rect -3344 -240 -3337 -176
rect -3413 -250 -3337 -240
rect -4604 -807 -4594 -755
rect -4542 -807 -4532 -755
rect -4734 -1048 -4724 -996
rect -4556 -1048 -4546 -996
rect -4547 -1266 -4537 -1090
rect -4485 -1266 -4475 -1090
rect -3433 -1267 -3423 -1090
rect -3371 -1267 -3361 -1090
rect -3074 -1325 -3028 1265
rect 18877 -851 18883 -727
rect 19007 -739 29120 -727
rect 19007 -839 28882 -739
rect 29120 -839 29130 -739
rect 19007 -851 29120 -839
rect 9397 -1238 19270 -1213
rect -2028 -1347 -2022 -1295
rect -1970 -1347 -250 -1295
rect 9397 -1310 9407 -1238
rect 9479 -1310 19270 -1238
rect 9397 -1337 19270 -1310
rect 19394 -1337 19404 -1213
rect -5562 -1380 -4928 -1374
rect -3423 -1396 -3371 -1390
rect -494 -1396 -442 -1390
rect -3371 -1448 -494 -1396
rect -3423 -1454 -3371 -1448
rect -494 -1454 -442 -1448
rect -1001 -1494 -949 -1488
rect -4543 -1546 -4537 -1494
rect -4485 -1546 -1001 -1494
rect -302 -1523 -250 -1347
rect -1001 -1552 -949 -1546
rect -308 -1575 -302 -1523
rect -250 -1575 -244 -1523
rect -2786 -1925 -138 -1918
rect -5598 -1974 -4883 -1928
rect -2786 -1977 -2780 -1925
rect -2728 -1977 -138 -1925
rect -86 -1977 -80 -1925
rect -2786 -1984 -138 -1977
rect 4494 -2367 4504 -2267
rect 4605 -2367 26531 -2267
rect 26631 -2367 26641 -2267
rect 8635 -2596 8645 -2496
rect 8744 -2596 26730 -2496
rect 26830 -2596 26840 -2496
rect 26778 -2602 26830 -2596
rect 9406 -2719 9416 -2663
rect 9472 -2719 9482 -2663
rect 13219 -2727 28694 -2714
rect -2732 -2817 -247 -2810
rect -5598 -2866 -4883 -2820
rect -2790 -2869 -2784 -2817
rect -2732 -2869 -305 -2817
rect -253 -2869 -247 -2817
rect -2732 -2876 -247 -2869
rect 13219 -2827 28579 -2727
rect 28679 -2827 28694 -2727
rect 13219 -2838 28694 -2827
rect 13219 -3026 13269 -2838
rect -138 -3084 -86 -3078
rect -86 -3135 272 -3085
rect -138 -3142 -86 -3136
rect -688 -3392 -682 -3326
rect -616 -3392 352 -3326
rect -2736 -3709 7 -3701
rect -5598 -3758 -4883 -3712
rect -2794 -3761 -2788 -3709
rect -2736 -3761 -50 -3709
rect 2 -3761 7 -3709
rect -2736 -3767 7 -3761
rect -305 -3988 -253 -3982
rect -253 -4039 189 -3989
rect -305 -4046 -253 -4040
rect 8674 -4441 8773 -4435
rect 8674 -4505 8686 -4441
rect 8761 -4505 8773 -4441
rect 8674 -4511 8773 -4505
rect -5598 -4650 -4883 -4604
rect -2776 -4662 -2770 -4596
rect -2704 -4662 -136 -4596
rect -70 -4662 -64 -4596
rect -501 -4730 8522 -4723
rect -501 -4782 -494 -4730
rect -442 -4782 8463 -4730
rect 8515 -4782 8522 -4730
rect -501 -4789 8522 -4782
rect -3855 -4910 -3845 -4858
rect -3069 -4910 -3059 -4858
rect -2774 -4916 -2768 -4850
rect -2702 -4916 -682 -4850
rect -616 -4916 -610 -4850
rect -1008 -5082 4184 -5075
rect -1008 -5134 -1001 -5082
rect -949 -5134 4126 -5082
rect 4178 -5134 4184 -5082
rect -1008 -5141 4184 -5134
rect 4097 -5142 4184 -5141
rect 8686 -5297 8761 -4511
rect 8965 -4566 19393 -4539
rect 8965 -4638 8991 -4566
rect 9063 -4638 19296 -4566
rect 19368 -4638 19393 -4566
rect 8965 -4663 19393 -4638
rect 18883 -4938 26437 -4919
rect 18883 -4940 26339 -4938
rect 18883 -5012 18902 -4940
rect 18974 -5010 26339 -4940
rect 26411 -5010 26437 -4938
rect 18974 -5012 26437 -5010
rect 18883 -5043 26437 -5012
rect 30277 -5401 30380 6533
rect 25619 -5504 30380 -5401
rect 25626 -5811 25636 -5759
rect 26033 -5811 26043 -5759
rect 4125 -6309 4135 -6257
rect 4187 -6309 4197 -6257
rect 8819 -6309 8829 -6257
rect 9226 -6309 9236 -6257
rect 8282 -6475 8292 -6423
rect 8689 -6475 8699 -6423
rect 25626 -6641 25636 -6589
rect 26033 -6641 26043 -6589
rect 25626 -6807 25636 -6755
rect 26033 -6807 26043 -6755
<< via1 >>
rect 17858 6998 17910 7050
rect 17231 5895 17283 5947
rect 19463 5895 19515 5947
rect 17858 5716 17910 5768
rect 16822 2790 18106 2842
rect 19160 2765 19240 2845
rect 19450 2765 19530 2845
rect -4243 327 -4059 379
rect -3408 -240 -3344 -176
rect -4594 -764 -4542 -755
rect -4594 -798 -4585 -764
rect -4585 -798 -4551 -764
rect -4551 -798 -4542 -764
rect -4594 -807 -4542 -798
rect -4724 -1048 -4556 -996
rect -4537 -1266 -4485 -1090
rect -3423 -1267 -3371 -1090
rect 18883 -851 19007 -727
rect 28882 -839 29120 -739
rect -2022 -1347 -1970 -1295
rect 9407 -1310 9479 -1238
rect 19270 -1337 19394 -1213
rect -3423 -1448 -3371 -1396
rect -494 -1448 -442 -1396
rect -4537 -1546 -4485 -1494
rect -1001 -1546 -949 -1494
rect -302 -1575 -250 -1523
rect -2780 -1977 -2728 -1925
rect -138 -1977 -86 -1925
rect 4504 -2367 4605 -2267
rect 26531 -2367 26631 -2267
rect 8645 -2596 8744 -2496
rect 26730 -2596 26830 -2496
rect 9416 -2719 9472 -2663
rect -2784 -2869 -2732 -2817
rect -305 -2869 -253 -2817
rect 28579 -2827 28679 -2727
rect -138 -3136 -86 -3084
rect -682 -3392 -616 -3326
rect -2788 -3761 -2736 -3709
rect -50 -3761 2 -3709
rect -305 -4040 -253 -3988
rect -2770 -4662 -2704 -4596
rect -136 -4662 -70 -4596
rect -494 -4782 -442 -4730
rect 8463 -4782 8515 -4730
rect -3845 -4910 -3069 -4858
rect -2768 -4916 -2702 -4850
rect -682 -4916 -616 -4850
rect -1001 -5134 -949 -5082
rect 4126 -5134 4178 -5082
rect 8991 -4638 9063 -4566
rect 19296 -4638 19368 -4566
rect 18902 -5012 18974 -4940
rect 26339 -5010 26411 -4938
rect 25636 -5811 26033 -5759
rect 4135 -6309 4187 -6257
rect 8829 -6309 9226 -6257
rect 8292 -6475 8689 -6423
rect 25636 -6641 26033 -6589
rect 25636 -6807 26033 -6755
<< metal2 >>
rect 17231 5947 17283 7177
rect 17858 7050 17910 7060
rect 17225 5895 17231 5947
rect 17283 5895 17289 5947
rect 17858 5768 17910 6998
rect 17858 5706 17910 5716
rect 19463 5947 19515 5953
rect 11086 3694 11138 3941
rect 11079 3684 11145 3694
rect 11079 3608 11145 3618
rect 18084 2928 19374 2986
rect 16822 2845 18106 2852
rect 16822 2842 19160 2845
rect 18106 2790 19160 2842
rect 16822 2787 19160 2790
rect 16822 2780 18106 2787
rect 18897 2765 19160 2787
rect 19240 2765 19246 2845
rect 9034 1546 9095 1549
rect 9027 1490 9036 1546
rect 9092 1490 9101 1546
rect -5534 379 -4059 389
rect -5534 327 -4243 379
rect -5534 317 -4059 327
rect -3948 -178 -3896 1257
rect -3408 -176 -3344 -166
rect -3408 -250 -3344 -240
rect -4594 -755 -4542 -745
rect -5559 -807 -4594 -755
rect -4594 -817 -4542 -807
rect -4724 -996 -4556 -986
rect -5561 -1048 -4724 -996
rect -4724 -1058 -4556 -1048
rect -4537 -1090 -4485 -1079
rect -4537 -1494 -4485 -1266
rect -3423 -1090 -3371 -1078
rect -3423 -1396 -3371 -1267
rect -2022 -1295 -1970 1244
rect 2464 -174 2530 -164
rect 2464 -250 2530 -240
rect 6580 -175 6646 -165
rect 2471 -1130 2523 -250
rect 6580 -251 6646 -241
rect 6587 -811 6639 -251
rect 9034 -1267 9095 1490
rect 18897 -721 18981 2765
rect 18883 -727 19007 -721
rect -2022 -1353 -1970 -1347
rect -3429 -1448 -3423 -1396
rect -3371 -1448 -3365 -1396
rect -501 -1448 -494 -1396
rect -442 -1448 -435 -1396
rect -1007 -1546 -1001 -1494
rect -949 -1546 -943 -1494
rect -4537 -1552 -4485 -1546
rect -3845 -1925 -2728 -1918
rect -3845 -1977 -2780 -1925
rect -3845 -1984 -2728 -1977
rect -3847 -2817 -2732 -2810
rect -3847 -2869 -2784 -2817
rect -3847 -2876 -2732 -2869
rect -3845 -3709 -2729 -3702
rect -3845 -3761 -2788 -3709
rect -2736 -3761 -2729 -3709
rect -3845 -3768 -2729 -3761
rect -2770 -4596 -2704 -4590
rect -3845 -4662 -2770 -4596
rect -2770 -4668 -2704 -4662
rect -3845 -4850 -3069 -4848
rect -2768 -4850 -2702 -4844
rect -3845 -4858 -2768 -4850
rect -3069 -4910 -2768 -4858
rect -3845 -4916 -2768 -4910
rect -3845 -4920 -3069 -4916
rect -2768 -4922 -2702 -4916
rect -1008 -5082 -942 -1546
rect -682 -3326 -616 -3320
rect -682 -4850 -616 -3392
rect -501 -4730 -435 -1448
rect -302 -1523 -250 -1517
rect 413 -1523 465 -1422
rect -250 -1575 465 -1523
rect -302 -1581 -250 -1575
rect -138 -1925 -86 -1919
rect -313 -2817 -247 -2810
rect -313 -2869 -305 -2817
rect -253 -2869 -247 -2817
rect -313 -3988 -247 -2869
rect -145 -3084 -79 -1977
rect 4505 -2257 4605 -1295
rect 8754 -1328 9095 -1267
rect 9380 -1238 9504 -1213
rect 9380 -1310 9407 -1238
rect 9479 -1310 9504 -1238
rect 8645 -1467 8697 -1413
rect 4504 -2267 4605 -2257
rect 4504 -2377 4605 -2367
rect 8644 -2496 8744 -1467
rect 8644 -2544 8645 -2496
rect 8645 -2606 8744 -2596
rect 9380 -2663 9504 -1310
rect 9415 -2719 9416 -2663
rect 9472 -2719 9473 -2663
rect 9415 -2720 9473 -2719
rect 9416 -2729 9472 -2720
rect -145 -3136 -138 -3084
rect -86 -3136 -79 -3084
rect -71 -3709 190 -3701
rect -71 -3761 -50 -3709
rect 2 -3761 190 -3709
rect -71 -3767 190 -3761
rect -313 -4040 -305 -3988
rect -253 -4040 -247 -3988
rect -313 -4046 -247 -4040
rect -131 -4239 -75 -4235
rect -136 -4244 -70 -4239
rect -136 -4300 -131 -4244
rect -75 -4300 -70 -4244
rect -136 -4596 -70 -4300
rect -136 -4668 -70 -4662
rect 8965 -4566 9089 -4539
rect 8965 -4638 8991 -4566
rect 9063 -4638 9089 -4566
rect -501 -4782 -494 -4730
rect -442 -4782 -435 -4730
rect -501 -4789 -435 -4782
rect 8456 -4730 8522 -4723
rect 8456 -4782 8463 -4730
rect 8515 -4782 8522 -4730
rect -682 -4922 -616 -4916
rect -1008 -5134 -1001 -5082
rect -949 -5134 -942 -5082
rect -1008 -5141 -942 -5134
rect 4126 -5082 4178 -5076
rect 4126 -6247 4178 -5134
rect 4126 -6255 4187 -6247
rect 4126 -6257 4200 -6255
rect 4126 -6307 4135 -6257
rect 4187 -6307 4200 -6257
rect 4135 -6319 4187 -6309
rect 8456 -6413 8522 -4782
rect 8965 -6247 9089 -4638
rect 18883 -4940 19007 -851
rect 19290 -1203 19374 2928
rect 19463 2851 19515 5895
rect 19450 2845 19530 2851
rect 19450 2759 19530 2765
rect 28882 -739 29120 -729
rect 29120 -839 29336 -739
rect 28882 -849 29120 -839
rect 19270 -1213 19394 -1203
rect 19270 -4566 19394 -1337
rect 28579 -2062 32605 -1962
rect 19270 -4638 19296 -4566
rect 19368 -4638 19394 -4566
rect 19270 -4662 19394 -4638
rect 26531 -2267 26631 -2257
rect 18883 -5012 18902 -4940
rect 18974 -5012 19007 -4940
rect 18883 -5022 19007 -5012
rect 26313 -4938 26437 -4919
rect 26313 -5010 26339 -4938
rect 26411 -5010 26437 -4938
rect 26313 -5749 26437 -5010
rect 25636 -5759 26437 -5749
rect 26033 -5811 26437 -5759
rect 25636 -5821 26437 -5811
rect 8829 -6257 9226 -6247
rect 8829 -6319 9226 -6309
rect 8292 -6423 8689 -6413
rect 8292 -6485 8689 -6475
rect 26531 -6579 26631 -2367
rect 25636 -6589 26631 -6579
rect 26033 -6641 26631 -6589
rect 25636 -6651 26631 -6641
rect 26730 -2495 26830 -2486
rect 26730 -2496 26836 -2495
rect 26830 -2596 26836 -2496
rect 26730 -2597 26836 -2596
rect 26730 -6745 26830 -2597
rect 28579 -2727 28679 -2062
rect 28573 -2827 28579 -2727
rect 28679 -2827 28685 -2727
rect 25636 -6755 26830 -6745
rect 25634 -6807 25636 -6755
rect 26033 -6807 26830 -6755
rect 25636 -6817 26830 -6807
<< via2 >>
rect 11079 3618 11145 3684
rect 9036 1490 9092 1546
rect -3408 -240 -3344 -176
rect 2464 -240 2530 -174
rect 6580 -241 6646 -175
rect 9416 -2719 9472 -2663
rect -131 -4300 -75 -4244
<< metal3 >>
rect 11062 3684 11162 3699
rect 11062 3618 11079 3684
rect 11145 3618 11162 3684
rect 11062 3599 11162 3618
rect 9031 1546 9097 1551
rect 9031 1490 9036 1546
rect 9092 1490 9097 1546
rect 9031 1485 9097 1490
rect -3428 -176 -3328 -157
rect -3428 -240 -3408 -176
rect -3344 -240 -3328 -176
rect -3428 -257 -3328 -240
rect 2449 -174 2549 -157
rect 2449 -240 2464 -174
rect 2530 -240 2549 -174
rect 2449 -257 2549 -240
rect 6563 -175 6663 -158
rect 6563 -241 6580 -175
rect 6646 -241 6663 -175
rect 6563 -258 6663 -241
rect 9396 -2659 9496 -2641
rect 9396 -2723 9412 -2659
rect 9476 -2723 9496 -2659
rect 9396 -2741 9496 -2723
rect -136 -4244 2600 -4239
rect -136 -4300 -131 -4244
rect -75 -4300 2600 -4244
rect -136 -4305 2600 -4300
<< via3 >>
rect 11079 3618 11145 3684
rect -3408 -240 -3344 -176
rect 2464 -240 2530 -174
rect 6580 -241 6646 -175
rect 9412 -2663 9476 -2659
rect 9412 -2719 9416 -2663
rect 9416 -2719 9472 -2663
rect 9472 -2719 9476 -2663
rect 9412 -2723 9476 -2719
<< metal4 >>
rect 11078 3684 11146 3685
rect 11078 3682 11079 3684
rect 8653 3618 11079 3682
rect 11145 3682 11146 3684
rect 15890 3682 15954 4789
rect 11145 3618 15954 3682
rect 2463 -174 2531 -173
rect -3409 -176 -3343 -175
rect 2463 -176 2464 -174
rect -3409 -240 -3408 -176
rect -3344 -240 2464 -176
rect 2530 -176 2531 -174
rect 6579 -175 6647 -174
rect 6579 -176 6580 -175
rect 2530 -240 6580 -176
rect -3409 -241 -3343 -240
rect 2463 -241 2531 -240
rect 6579 -241 6580 -240
rect 6646 -176 6647 -175
rect 8653 -176 8717 3618
rect 11078 3617 11146 3618
rect 6646 -240 8717 -176
rect 6646 -241 6647 -240
rect 6579 -242 6647 -241
rect 9411 -2659 9477 -2658
rect 9411 -2723 9412 -2659
rect 9476 -2723 9477 -2659
rect 9411 -2973 9477 -2723
use bjt  bjt_0
timestamp 1764413320
transform -1 0 36957 0 -1 2857
box 0 0 7749 7292
use digital  digital_0
timestamp 1764411030
transform 1 0 -4922 0 1 -4244
box -108 -870 2044 4722
use op5  op5_0
timestamp 1762874782
transform 1 0 9786 0 1 -6121
box -9786 6121 9272 13721
use pmos_current_bgr  pmos_current_bgr_0
timestamp 1762875002
transform 1 0 425 0 1 -1186
box -227 -676 8487 506
use res_trim  res_trim_0
timestamp 1762873293
transform 0 1 101 -1 0 -2857
box -31 -51 1533 15873
use resist_const  resist_const_0
timestamp 1762877483
transform -1 0 28465 0 -1 -9225
box 2257 -4057 28483 -2103
use startupcir  startupcir_0
timestamp 1762846550
transform -1 0 21906 0 -1 7909
box -20 -1581 21888 938
<< labels >>
flabel metal2 -3923 1228 -3923 1228 0 FreeSans 1600 0 0 0 avdd
port 0 nsew
flabel metal1 -5553 -1950 -5553 -1950 0 FreeSans 1600 0 0 0 trim0
port 5 nsew
flabel metal1 -5553 -2846 -5553 -2846 0 FreeSans 1600 0 0 0 trim1
port 6 nsew
flabel metal1 -5551 -3734 -5551 -3734 0 FreeSans 1600 0 0 0 trim2
port 7 nsew
flabel metal1 -5553 -4629 -5553 -4629 0 FreeSans 1600 0 0 0 trim3
port 8 nsew
flabel metal1 -3054 1242 -3054 1242 0 FreeSans 1600 0 0 0 vbgsc
port 9 nsew
flabel metal1 -4856 1187 -4856 1187 0 FreeSans 1600 0 0 0 vbgtc
port 10 nsew
flabel metal2 -5533 -782 -5533 -782 0 FreeSans 1600 0 0 0 dvdd
port 2 nsew
flabel metal1 -5531 -1358 -5531 -1358 0 FreeSans 1600 0 0 0 dvss
port 3 nsew
flabel metal2 -1992 1209 -1992 1209 0 FreeSans 1600 0 0 0 vref
port 12 nsew
flabel metal2 -5533 -1027 -5533 -1027 0 FreeSans 1600 0 0 0 vena
port 11 nsew
flabel metal2 -5501 350 -5501 350 0 FreeSans 1600 0 0 0 ena
port 4 nsew
flabel metal1 30340 5347 30340 5347 0 FreeSans 1600 0 0 0 avss
port 1 nsew
<< end >>
