magic
tech sky130A
magscale 1 2
timestamp 1717985588
<< nwell >>
rect -227 -1493 8585 556
<< nsubdiff >>
rect -191 486 -131 520
rect 8489 486 8549 520
rect -191 460 -157 486
rect 8515 460 8549 486
rect -191 -1423 -157 -1397
rect 8515 -1423 8549 -1397
rect -191 -1457 -131 -1423
rect 8489 -1457 8549 -1423
<< nsubdiffcont >>
rect -131 486 8489 520
rect -191 -1397 -157 460
rect 8515 -1397 8549 460
rect -131 -1457 8489 -1423
<< poly >>
rect -58 426 34 442
rect -58 392 -42 426
rect -8 392 34 426
rect -58 376 34 392
rect 4 368 34 376
rect 8324 426 8416 442
rect 8324 392 8366 426
rect 8400 392 8416 426
rect 8324 376 8416 392
rect 8324 345 8354 376
rect 4 -436 34 -348
rect -58 -452 34 -436
rect -58 -486 -42 -452
rect -8 -486 34 -452
rect -58 -502 34 -486
rect 4 -592 34 -502
rect 92 -540 8266 -398
rect 8324 -436 8354 -346
rect 8324 -452 8416 -436
rect 8324 -486 8366 -452
rect 8400 -486 8416 -452
rect 8324 -502 8416 -486
rect 8324 -578 8354 -502
rect 4 -1314 34 -1298
rect -58 -1330 34 -1314
rect -58 -1364 -42 -1330
rect -8 -1364 34 -1330
rect -58 -1380 34 -1364
rect 8324 -1314 8354 -1283
rect 8324 -1330 8416 -1314
rect 8324 -1364 8366 -1330
rect 8400 -1364 8416 -1330
rect 8324 -1380 8416 -1364
<< polycont >>
rect -42 392 -8 426
rect 8366 392 8400 426
rect -42 -486 -8 -452
rect 8366 -486 8400 -452
rect -42 -1364 -8 -1330
rect 8366 -1364 8400 -1330
<< locali >>
rect -191 486 -131 520
rect 8489 486 8549 520
rect -191 460 -157 486
rect 8515 460 8549 486
rect -42 426 -8 442
rect -42 343 -8 392
rect 8366 426 8400 442
rect 8366 345 8400 392
rect -42 -452 -8 -436
rect -42 -502 -8 -486
rect 8366 -452 8400 -436
rect 8366 -502 8400 -486
rect -42 -1330 -8 -1286
rect -42 -1380 -8 -1364
rect 8366 -1330 8400 -1283
rect 8366 -1380 8400 -1364
rect -191 -1423 -157 -1397
rect 8515 -1423 8549 -1397
rect -191 -1457 -131 -1423
rect 8489 -1457 8549 -1423
<< viali >>
rect -42 486 -8 520
rect 2104 486 2138 520
rect 4162 486 4196 520
rect 6220 486 6254 520
rect 8366 486 8400 520
rect -42 392 -8 426
rect 8366 392 8400 426
rect -191 -486 -157 -452
rect -42 -486 -8 -452
rect 8366 -486 8400 -452
rect 8515 -486 8549 -452
rect -42 -1364 -8 -1330
rect 8366 -1364 8400 -1330
rect -42 -1457 -8 -1423
rect 2104 -1457 2138 -1423
rect 4162 -1457 4196 -1423
rect 6220 -1457 6254 -1423
rect 8366 -1457 8400 -1423
<< metal1 >>
rect -48 520 -2 532
rect -48 486 -42 520
rect -8 486 -2 520
rect -48 426 -2 486
rect -48 392 -42 426
rect -8 392 -2 426
rect -48 342 -2 392
rect 2098 520 2144 532
rect 2098 486 2104 520
rect 2138 486 2144 520
rect 2098 333 2144 486
rect 4156 520 4202 532
rect 4156 486 4162 520
rect 4196 486 4202 520
rect 27 157 37 333
rect 89 157 99 333
rect 2085 157 2095 333
rect 2147 157 2157 333
rect 4156 327 4202 486
rect 6214 520 6260 532
rect 6214 486 6220 520
rect 6254 486 6260 520
rect 6214 333 6260 486
rect 8360 520 8406 532
rect 8360 486 8366 520
rect 8400 486 8406 520
rect 8360 426 8406 486
rect 8360 392 8366 426
rect 8400 392 8406 426
rect 8360 345 8406 392
rect 6201 157 6211 333
rect 6263 157 6273 333
rect 8259 157 8269 333
rect 8321 157 8331 333
rect 4156 104 4202 152
rect -152 -19 -142 33
rect -90 30 -80 33
rect 588 30 1596 67
rect 3633 58 4730 104
rect 6762 30 7770 62
rect 8438 30 8448 33
rect -90 -16 8448 30
rect -90 -19 -80 -16
rect 8438 -19 8448 -16
rect 8500 -19 8510 33
rect 590 -96 600 -44
rect 1584 -47 1594 -44
rect 6764 -47 6774 -44
rect 1584 -93 6774 -47
rect 1584 -96 1594 -93
rect 6764 -96 6774 -93
rect 7758 -96 7768 -44
rect -48 -440 -2 -313
rect -197 -452 -2 -440
rect 40 -443 86 -320
rect 2085 -322 2095 -146
rect 2147 -322 2157 -146
rect 4143 -322 4153 -146
rect 4205 -322 4215 -146
rect 6201 -322 6211 -146
rect 6263 -322 6273 -146
rect -197 -486 -191 -452
rect -157 -486 -42 -452
rect -8 -486 -2 -452
rect -197 -498 -2 -486
rect 27 -495 37 -443
rect 89 -495 99 -443
rect 588 -452 1596 -414
rect 6762 -452 7770 -419
rect 8272 -443 8318 -316
rect 8360 -440 8406 -309
rect 588 -486 7770 -452
rect -48 -614 -2 -498
rect 40 -618 86 -495
rect 588 -523 1596 -486
rect 6762 -528 7770 -486
rect 8259 -495 8269 -443
rect 8321 -495 8331 -443
rect 8360 -452 8555 -440
rect 8360 -486 8366 -452
rect 8400 -486 8515 -452
rect 8549 -486 8555 -452
rect 8272 -614 8318 -495
rect 8360 -498 8555 -486
rect 8360 -610 8406 -498
rect 2085 -792 2095 -616
rect 2147 -792 2157 -616
rect 4143 -792 4153 -616
rect 4205 -792 4215 -616
rect 6201 -792 6211 -616
rect 6263 -792 6273 -616
rect 590 -894 600 -842
rect 1584 -845 1594 -842
rect 1584 -891 6762 -845
rect 1584 -894 1594 -891
rect 6764 -894 6774 -842
rect 7758 -894 7768 -842
rect -152 -971 -142 -919
rect -90 -922 -80 -919
rect 8438 -922 8448 -919
rect -90 -968 8448 -922
rect -90 -971 -80 -968
rect 588 -1009 1596 -968
rect 3639 -1042 4736 -996
rect 6762 -1001 7770 -968
rect 8438 -971 8448 -968
rect 8500 -971 8510 -919
rect -48 -1330 -2 -1250
rect 27 -1271 37 -1095
rect 89 -1271 99 -1095
rect 2085 -1271 2095 -1095
rect 2147 -1271 2157 -1095
rect 4156 -1097 4202 -1042
rect -48 -1364 -42 -1330
rect -8 -1364 -2 -1330
rect -48 -1423 -2 -1364
rect -48 -1457 -42 -1423
rect -8 -1457 -2 -1423
rect -48 -1469 -2 -1457
rect 2098 -1423 2144 -1271
rect 2098 -1457 2104 -1423
rect 2138 -1457 2144 -1423
rect 2098 -1469 2144 -1457
rect 4156 -1423 4202 -1251
rect 6201 -1271 6211 -1095
rect 6263 -1271 6273 -1095
rect 8259 -1271 8269 -1095
rect 8321 -1271 8331 -1095
rect 4156 -1457 4162 -1423
rect 4196 -1457 4202 -1423
rect 4156 -1469 4202 -1457
rect 6214 -1423 6260 -1271
rect 6214 -1457 6220 -1423
rect 6254 -1457 6260 -1423
rect 6214 -1469 6260 -1457
rect 8360 -1330 8406 -1283
rect 8360 -1364 8366 -1330
rect 8400 -1364 8406 -1330
rect 8360 -1423 8406 -1364
rect 8360 -1457 8366 -1423
rect 8400 -1457 8406 -1423
rect 8360 -1469 8406 -1457
<< via1 >>
rect 37 157 89 333
rect 2095 157 2147 333
rect 6211 157 6263 333
rect 8269 157 8321 333
rect -142 -19 -90 33
rect 8448 -19 8500 33
rect 600 -96 1584 -44
rect 6774 -96 7758 -44
rect 2095 -322 2147 -146
rect 4153 -322 4205 -146
rect 6211 -322 6263 -146
rect 37 -495 89 -443
rect 8269 -495 8321 -443
rect 2095 -792 2147 -616
rect 4153 -792 4205 -616
rect 6211 -792 6263 -616
rect 600 -894 1584 -842
rect 6774 -894 7758 -842
rect -142 -971 -90 -919
rect 8448 -971 8500 -919
rect 37 -1271 89 -1095
rect 2095 -1271 2147 -1095
rect 6211 -1271 6263 -1095
rect 8269 -1271 8321 -1095
<< metal2 >>
rect 37 383 8321 435
rect 37 343 89 383
rect 8269 343 8321 383
rect 35 333 91 343
rect 35 147 91 157
rect 2095 333 2147 343
rect -142 33 -90 43
rect -142 -919 -90 -19
rect 600 -42 1584 -32
rect 600 -108 1584 -98
rect 2095 -146 2147 157
rect 6211 333 6263 343
rect 35 -441 91 -431
rect 35 -507 91 -497
rect 2095 -616 2147 -322
rect 600 -840 1584 -830
rect 600 -906 1584 -896
rect -142 -981 -90 -971
rect 35 -1095 91 -1085
rect 35 -1281 91 -1271
rect 2095 -1095 2147 -792
rect 4153 -146 4205 -136
rect 4153 -616 4205 -322
rect 4153 -802 4205 -792
rect 6211 -146 6263 157
rect 8267 333 8323 343
rect 8267 147 8323 157
rect 8448 33 8500 43
rect 6774 -42 7758 -32
rect 6774 -108 7758 -98
rect 6211 -616 6263 -322
rect 8267 -441 8323 -431
rect 8267 -507 8323 -497
rect 2095 -1281 2147 -1271
rect 6211 -1095 6263 -792
rect 6774 -840 7758 -830
rect 6774 -906 7758 -896
rect 8448 -919 8500 -19
rect 8448 -981 8500 -971
rect 6211 -1281 6263 -1271
rect 8267 -1095 8323 -1085
rect 8267 -1281 8323 -1271
rect 37 -1321 89 -1281
rect 8269 -1321 8321 -1281
rect 37 -1373 8321 -1321
<< via2 >>
rect 35 157 37 333
rect 37 157 89 333
rect 89 157 91 333
rect 600 -44 1584 -42
rect 600 -96 1584 -44
rect 600 -98 1584 -96
rect 35 -443 91 -441
rect 35 -495 37 -443
rect 37 -495 89 -443
rect 89 -495 91 -443
rect 35 -497 91 -495
rect 600 -842 1584 -840
rect 600 -894 1584 -842
rect 600 -896 1584 -894
rect 35 -1271 37 -1095
rect 37 -1271 89 -1095
rect 89 -1271 91 -1095
rect 8267 157 8269 333
rect 8269 157 8321 333
rect 8321 157 8323 333
rect 6774 -44 7758 -42
rect 6774 -96 7758 -44
rect 6774 -98 7758 -96
rect 8267 -443 8323 -441
rect 8267 -495 8269 -443
rect 8269 -495 8321 -443
rect 8321 -495 8323 -443
rect 8267 -497 8323 -495
rect 6774 -842 7758 -840
rect 6774 -894 7758 -842
rect 6774 -896 7758 -894
rect 8267 -1271 8269 -1095
rect 8269 -1271 8321 -1095
rect 8321 -1271 8323 -1095
<< metal3 >>
rect 25 333 101 338
rect 25 157 35 333
rect 91 157 101 333
rect 25 152 101 157
rect 8257 333 8333 338
rect 8257 157 8267 333
rect 8323 157 8333 333
rect 8257 152 8333 157
rect 33 43 93 152
rect 8265 43 8325 152
rect -142 -17 650 43
rect -142 -921 -82 -17
rect 590 -37 650 -17
rect 7708 -17 8500 43
rect 7708 -37 7768 -17
rect 590 -42 1594 -37
rect 590 -98 600 -42
rect 1584 -98 1594 -42
rect 590 -103 1594 -98
rect 6764 -42 7768 -37
rect 6764 -98 6774 -42
rect 7758 -98 7768 -42
rect 6764 -103 7768 -98
rect 25 -439 101 -436
rect 8257 -439 8333 -436
rect 25 -441 8333 -439
rect 25 -497 35 -441
rect 91 -497 8267 -441
rect 8323 -497 8333 -441
rect 25 -499 8333 -497
rect 25 -502 101 -499
rect 8257 -502 8333 -499
rect 590 -840 1594 -835
rect 590 -896 600 -840
rect 1584 -896 1594 -840
rect 590 -901 1594 -896
rect 6764 -840 7768 -835
rect 6764 -896 6774 -840
rect 7758 -896 7768 -840
rect 6764 -901 7768 -896
rect 590 -921 650 -901
rect -142 -981 650 -921
rect 7708 -921 7768 -901
rect 8440 -921 8500 -17
rect 7708 -981 8500 -921
rect 33 -1090 93 -981
rect 8265 -1090 8325 -981
rect 25 -1095 101 -1090
rect 25 -1271 35 -1095
rect 91 -1271 101 -1095
rect 25 -1276 101 -1271
rect 8257 -1095 8333 -1090
rect 8257 -1271 8267 -1095
rect 8323 -1271 8333 -1095
rect 8257 -1276 8333 -1271
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_0
timestamp 1717765832
transform 1 0 19 0 1 -704
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_1
timestamp 1717765832
transform 1 0 8339 0 1 -1183
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_2
timestamp 1717765832
transform 1 0 8339 0 1 -704
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_3
timestamp 1717765832
transform 1 0 8339 0 1 -234
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_4
timestamp 1717765832
transform 1 0 8339 0 1 245
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_5
timestamp 1717765832
transform 1 0 19 0 1 245
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_6
timestamp 1717765832
transform 1 0 19 0 1 -234
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_8
timestamp 1717765832
transform 1 0 19 0 1 -1183
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_8WJJP2  sky130_fd_pr__pfet_01v8_8WJJP2_1
timestamp 1717408091
transform 1 0 4179 0 1 -1147
box -4181 -198 4181 164
use sky130_fd_pr__pfet_01v8_C2SJBD  sky130_fd_pr__pfet_01v8_C2SJBD_0
timestamp 1717408091
transform 1 0 4179 0 1 209
box -4181 -164 4181 198
use sky130_fd_pr__pfet_01v8_HVJJBB  sky130_fd_pr__pfet_01v8_HVJJBB_0
timestamp 1717985045
transform 1 0 4179 0 1 -234
box -4181 -200 4181 200
use sky130_fd_pr__pfet_01v8_HVJJBB  sky130_fd_pr__pfet_01v8_HVJJBB_1
timestamp 1717985045
transform 1 0 4179 0 1 -704
box -4181 -200 4181 200
<< labels >>
flabel metal3 8286 74 8286 74 0 FreeSans 800 0 0 0 D10
port 0 nsew
flabel metal1 8289 -389 8289 -389 0 FreeSans 800 0 0 0 D2
port 1 nsew
flabel metal2 4178 -374 4178 -374 0 FreeSans 800 0 0 0 D1
port 2 nsew
flabel metal1 6234 -1407 6234 -1407 0 FreeSans 800 0 0 0 vdde
port 3 nsew
flabel metal1 7457 29 7457 29 0 FreeSans 800 0 0 0 G10
port 4 nsew
<< end >>
