magic
tech sky130A
magscale 1 2
timestamp 1716351939
<< nwell >>
rect -511 -2235 511 2235
<< nsubdiff >>
rect -475 2165 -379 2199
rect 379 2165 475 2199
rect -475 2103 -441 2165
rect 441 2103 475 2165
rect -475 -2165 -441 -2103
rect 441 -2165 475 -2103
rect -475 -2199 -379 -2165
rect 379 -2199 475 -2165
<< nsubdiffcont >>
rect -379 2165 379 2199
rect -475 -2103 -441 2103
rect 441 -2103 475 2103
rect -379 -2199 379 -2165
<< xpolycontact >>
rect -284 1628 -214 2060
rect -284 1108 -214 1540
rect -118 1628 -48 2060
rect -118 1108 -48 1540
rect 48 1628 118 2060
rect 48 1108 118 1540
rect 214 1628 284 2060
rect 214 1108 284 1540
rect -284 572 -214 1004
rect -284 52 -214 484
rect -118 572 -48 1004
rect -118 52 -48 484
rect 48 572 118 1004
rect 48 52 118 484
rect 214 572 284 1004
rect 214 52 284 484
rect -284 -484 -214 -52
rect -284 -1004 -214 -572
rect -118 -484 -48 -52
rect -118 -1004 -48 -572
rect 48 -484 118 -52
rect 48 -1004 118 -572
rect 214 -484 284 -52
rect 214 -1004 284 -572
rect -284 -1540 -214 -1108
rect -284 -2060 -214 -1628
rect -118 -1540 -48 -1108
rect -118 -2060 -48 -1628
rect 48 -1540 118 -1108
rect 48 -2060 118 -1628
rect 214 -1540 284 -1108
rect 214 -2060 284 -1628
<< ppolyres >>
rect -284 1540 -214 1628
rect -118 1540 -48 1628
rect 48 1540 118 1628
rect 214 1540 284 1628
rect -284 484 -214 572
rect -118 484 -48 572
rect 48 484 118 572
rect 214 484 284 572
rect -284 -572 -214 -484
rect -118 -572 -48 -484
rect 48 -572 118 -484
rect 214 -572 284 -484
rect -284 -1628 -214 -1540
rect -118 -1628 -48 -1540
rect 48 -1628 118 -1540
rect 214 -1628 284 -1540
<< locali >>
rect -475 2165 -379 2199
rect 379 2165 475 2199
rect -475 2103 -441 2165
rect 441 2103 475 2165
rect -475 -2165 -441 -2103
rect 441 -2165 475 -2103
rect -475 -2199 -379 -2165
rect 379 -2199 475 -2165
<< viali >>
rect -268 1645 -230 2042
rect -102 1645 -64 2042
rect 64 1645 102 2042
rect 230 1645 268 2042
rect -268 1126 -230 1523
rect -102 1126 -64 1523
rect 64 1126 102 1523
rect 230 1126 268 1523
rect -268 589 -230 986
rect -102 589 -64 986
rect 64 589 102 986
rect 230 589 268 986
rect -268 70 -230 467
rect -102 70 -64 467
rect 64 70 102 467
rect 230 70 268 467
rect -268 -467 -230 -70
rect -102 -467 -64 -70
rect 64 -467 102 -70
rect 230 -467 268 -70
rect -268 -986 -230 -589
rect -102 -986 -64 -589
rect 64 -986 102 -589
rect 230 -986 268 -589
rect -268 -1523 -230 -1126
rect -102 -1523 -64 -1126
rect 64 -1523 102 -1126
rect 230 -1523 268 -1126
rect -268 -2042 -230 -1645
rect -102 -2042 -64 -1645
rect 64 -2042 102 -1645
rect 230 -2042 268 -1645
<< metal1 >>
rect -274 2042 -224 2054
rect -274 1645 -268 2042
rect -230 1645 -224 2042
rect -274 1633 -224 1645
rect -108 2042 -58 2054
rect -108 1645 -102 2042
rect -64 1645 -58 2042
rect -108 1633 -58 1645
rect 58 2042 108 2054
rect 58 1645 64 2042
rect 102 1645 108 2042
rect 58 1633 108 1645
rect 224 2042 274 2054
rect 224 1645 230 2042
rect 268 1645 274 2042
rect 224 1633 274 1645
rect -274 1523 -224 1535
rect -274 1126 -268 1523
rect -230 1126 -224 1523
rect -274 1114 -224 1126
rect -108 1523 -58 1535
rect -108 1126 -102 1523
rect -64 1126 -58 1523
rect -108 1114 -58 1126
rect 58 1523 108 1535
rect 58 1126 64 1523
rect 102 1126 108 1523
rect 58 1114 108 1126
rect 224 1523 274 1535
rect 224 1126 230 1523
rect 268 1126 274 1523
rect 224 1114 274 1126
rect -274 986 -224 998
rect -274 589 -268 986
rect -230 589 -224 986
rect -274 577 -224 589
rect -108 986 -58 998
rect -108 589 -102 986
rect -64 589 -58 986
rect -108 577 -58 589
rect 58 986 108 998
rect 58 589 64 986
rect 102 589 108 986
rect 58 577 108 589
rect 224 986 274 998
rect 224 589 230 986
rect 268 589 274 986
rect 224 577 274 589
rect -274 467 -224 479
rect -274 70 -268 467
rect -230 70 -224 467
rect -274 58 -224 70
rect -108 467 -58 479
rect -108 70 -102 467
rect -64 70 -58 467
rect -108 58 -58 70
rect 58 467 108 479
rect 58 70 64 467
rect 102 70 108 467
rect 58 58 108 70
rect 224 467 274 479
rect 224 70 230 467
rect 268 70 274 467
rect 224 58 274 70
rect -274 -70 -224 -58
rect -274 -467 -268 -70
rect -230 -467 -224 -70
rect -274 -479 -224 -467
rect -108 -70 -58 -58
rect -108 -467 -102 -70
rect -64 -467 -58 -70
rect -108 -479 -58 -467
rect 58 -70 108 -58
rect 58 -467 64 -70
rect 102 -467 108 -70
rect 58 -479 108 -467
rect 224 -70 274 -58
rect 224 -467 230 -70
rect 268 -467 274 -70
rect 224 -479 274 -467
rect -274 -589 -224 -577
rect -274 -986 -268 -589
rect -230 -986 -224 -589
rect -274 -998 -224 -986
rect -108 -589 -58 -577
rect -108 -986 -102 -589
rect -64 -986 -58 -589
rect -108 -998 -58 -986
rect 58 -589 108 -577
rect 58 -986 64 -589
rect 102 -986 108 -589
rect 58 -998 108 -986
rect 224 -589 274 -577
rect 224 -986 230 -589
rect 268 -986 274 -589
rect 224 -998 274 -986
rect -274 -1126 -224 -1114
rect -274 -1523 -268 -1126
rect -230 -1523 -224 -1126
rect -274 -1535 -224 -1523
rect -108 -1126 -58 -1114
rect -108 -1523 -102 -1126
rect -64 -1523 -58 -1126
rect -108 -1535 -58 -1523
rect 58 -1126 108 -1114
rect 58 -1523 64 -1126
rect 102 -1523 108 -1126
rect 58 -1535 108 -1523
rect 224 -1126 274 -1114
rect 224 -1523 230 -1126
rect 268 -1523 274 -1126
rect 224 -1535 274 -1523
rect -274 -1645 -224 -1633
rect -274 -2042 -268 -1645
rect -230 -2042 -224 -1645
rect -274 -2054 -224 -2042
rect -108 -1645 -58 -1633
rect -108 -2042 -102 -1645
rect -64 -2042 -58 -1645
rect -108 -2054 -58 -2042
rect 58 -1645 108 -1633
rect 58 -2042 64 -1645
rect 102 -2042 108 -1645
rect 58 -2054 108 -2042
rect 224 -1645 274 -1633
rect 224 -2042 230 -1645
rect 268 -2042 274 -1645
rect 224 -2054 274 -2042
<< properties >>
string FIXED_BBOX -458 -2182 458 2182
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.350 l 0.6 m 4 nx 4 wmin 0.350 lmin 0.50 rho 319.8 val 1.661k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.350 vias 1 n_guard 1 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
