magic
tech sky130A
magscale 1 2
timestamp 1717227529
<< nwell >>
rect -812 -537 812 537
<< pmos >>
rect -616 118 -416 318
rect -358 118 -158 318
rect -100 118 100 318
rect 158 118 358 318
rect 416 118 616 318
rect -616 -318 -416 -118
rect -358 -318 -158 -118
rect -100 -318 100 -118
rect 158 -318 358 -118
rect 416 -318 616 -118
<< pdiff >>
rect -674 306 -616 318
rect -674 130 -662 306
rect -628 130 -616 306
rect -674 118 -616 130
rect -416 306 -358 318
rect -416 130 -404 306
rect -370 130 -358 306
rect -416 118 -358 130
rect -158 306 -100 318
rect -158 130 -146 306
rect -112 130 -100 306
rect -158 118 -100 130
rect 100 306 158 318
rect 100 130 112 306
rect 146 130 158 306
rect 100 118 158 130
rect 358 306 416 318
rect 358 130 370 306
rect 404 130 416 306
rect 358 118 416 130
rect 616 306 674 318
rect 616 130 628 306
rect 662 130 674 306
rect 616 118 674 130
rect -674 -130 -616 -118
rect -674 -306 -662 -130
rect -628 -306 -616 -130
rect -674 -318 -616 -306
rect -416 -130 -358 -118
rect -416 -306 -404 -130
rect -370 -306 -358 -130
rect -416 -318 -358 -306
rect -158 -130 -100 -118
rect -158 -306 -146 -130
rect -112 -306 -100 -130
rect -158 -318 -100 -306
rect 100 -130 158 -118
rect 100 -306 112 -130
rect 146 -306 158 -130
rect 100 -318 158 -306
rect 358 -130 416 -118
rect 358 -306 370 -130
rect 404 -306 416 -130
rect 358 -318 416 -306
rect 616 -130 674 -118
rect 616 -306 628 -130
rect 662 -306 674 -130
rect 616 -318 674 -306
<< pdiffc >>
rect -662 130 -628 306
rect -404 130 -370 306
rect -146 130 -112 306
rect 112 130 146 306
rect 370 130 404 306
rect 628 130 662 306
rect -662 -306 -628 -130
rect -404 -306 -370 -130
rect -146 -306 -112 -130
rect 112 -306 146 -130
rect 370 -306 404 -130
rect 628 -306 662 -130
<< nsubdiff >>
rect -776 467 -680 501
rect 680 467 776 501
rect -776 405 -742 467
rect 742 405 776 467
rect -776 -467 -742 -405
rect 742 -467 776 -405
rect -776 -501 -680 -467
rect 680 -501 776 -467
<< nsubdiffcont >>
rect -680 467 680 501
rect -776 -405 -742 405
rect 742 -405 776 405
rect -680 -501 680 -467
<< poly >>
rect -616 399 -416 415
rect -616 365 -600 399
rect -432 365 -416 399
rect -616 318 -416 365
rect -358 399 -158 415
rect -358 365 -342 399
rect -174 365 -158 399
rect -358 318 -158 365
rect -100 399 100 415
rect -100 365 -84 399
rect 84 365 100 399
rect -100 318 100 365
rect 158 399 358 415
rect 158 365 174 399
rect 342 365 358 399
rect 158 318 358 365
rect 416 399 616 415
rect 416 365 432 399
rect 600 365 616 399
rect 416 318 616 365
rect -616 71 -416 118
rect -616 37 -600 71
rect -432 37 -416 71
rect -616 21 -416 37
rect -358 71 -158 118
rect -358 37 -342 71
rect -174 37 -158 71
rect -358 21 -158 37
rect -100 71 100 118
rect -100 37 -84 71
rect 84 37 100 71
rect -100 21 100 37
rect 158 71 358 118
rect 158 37 174 71
rect 342 37 358 71
rect 158 21 358 37
rect 416 71 616 118
rect 416 37 432 71
rect 600 37 616 71
rect 416 21 616 37
rect -616 -37 -416 -21
rect -616 -71 -600 -37
rect -432 -71 -416 -37
rect -616 -118 -416 -71
rect -358 -37 -158 -21
rect -358 -71 -342 -37
rect -174 -71 -158 -37
rect -358 -118 -158 -71
rect -100 -37 100 -21
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -100 -118 100 -71
rect 158 -37 358 -21
rect 158 -71 174 -37
rect 342 -71 358 -37
rect 158 -118 358 -71
rect 416 -37 616 -21
rect 416 -71 432 -37
rect 600 -71 616 -37
rect 416 -118 616 -71
rect -616 -365 -416 -318
rect -616 -399 -600 -365
rect -432 -399 -416 -365
rect -616 -415 -416 -399
rect -358 -365 -158 -318
rect -358 -399 -342 -365
rect -174 -399 -158 -365
rect -358 -415 -158 -399
rect -100 -365 100 -318
rect -100 -399 -84 -365
rect 84 -399 100 -365
rect -100 -415 100 -399
rect 158 -365 358 -318
rect 158 -399 174 -365
rect 342 -399 358 -365
rect 158 -415 358 -399
rect 416 -365 616 -318
rect 416 -399 432 -365
rect 600 -399 616 -365
rect 416 -415 616 -399
<< polycont >>
rect -600 365 -432 399
rect -342 365 -174 399
rect -84 365 84 399
rect 174 365 342 399
rect 432 365 600 399
rect -600 37 -432 71
rect -342 37 -174 71
rect -84 37 84 71
rect 174 37 342 71
rect 432 37 600 71
rect -600 -71 -432 -37
rect -342 -71 -174 -37
rect -84 -71 84 -37
rect 174 -71 342 -37
rect 432 -71 600 -37
rect -600 -399 -432 -365
rect -342 -399 -174 -365
rect -84 -399 84 -365
rect 174 -399 342 -365
rect 432 -399 600 -365
<< locali >>
rect -776 467 -680 501
rect 680 467 776 501
rect -776 405 -742 467
rect 742 405 776 467
rect -616 365 -600 399
rect -432 365 -416 399
rect -358 365 -342 399
rect -174 365 -158 399
rect -100 365 -84 399
rect 84 365 100 399
rect 158 365 174 399
rect 342 365 358 399
rect 416 365 432 399
rect 600 365 616 399
rect -662 306 -628 322
rect -662 114 -628 130
rect -404 306 -370 322
rect -404 114 -370 130
rect -146 306 -112 322
rect -146 114 -112 130
rect 112 306 146 322
rect 112 114 146 130
rect 370 306 404 322
rect 370 114 404 130
rect 628 306 662 322
rect 628 114 662 130
rect -616 37 -600 71
rect -432 37 -416 71
rect -358 37 -342 71
rect -174 37 -158 71
rect -100 37 -84 71
rect 84 37 100 71
rect 158 37 174 71
rect 342 37 358 71
rect 416 37 432 71
rect 600 37 616 71
rect -616 -71 -600 -37
rect -432 -71 -416 -37
rect -358 -71 -342 -37
rect -174 -71 -158 -37
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect 158 -71 174 -37
rect 342 -71 358 -37
rect 416 -71 432 -37
rect 600 -71 616 -37
rect -662 -130 -628 -114
rect -662 -322 -628 -306
rect -404 -130 -370 -114
rect -404 -322 -370 -306
rect -146 -130 -112 -114
rect -146 -322 -112 -306
rect 112 -130 146 -114
rect 112 -322 146 -306
rect 370 -130 404 -114
rect 370 -322 404 -306
rect 628 -130 662 -114
rect 628 -322 662 -306
rect -616 -399 -600 -365
rect -432 -399 -416 -365
rect -358 -399 -342 -365
rect -174 -399 -158 -365
rect -100 -399 -84 -365
rect 84 -399 100 -365
rect 158 -399 174 -365
rect 342 -399 358 -365
rect 416 -399 432 -365
rect 600 -399 616 -365
rect -776 -467 -742 -405
rect 742 -467 776 -405
rect -776 -501 -680 -467
rect 680 -501 776 -467
<< viali >>
rect -600 365 -432 399
rect -342 365 -174 399
rect -84 365 84 399
rect 174 365 342 399
rect 432 365 600 399
rect -662 130 -628 306
rect -404 130 -370 306
rect -146 130 -112 306
rect 112 130 146 306
rect 370 130 404 306
rect 628 130 662 306
rect -600 37 -432 71
rect -342 37 -174 71
rect -84 37 84 71
rect 174 37 342 71
rect 432 37 600 71
rect -600 -71 -432 -37
rect -342 -71 -174 -37
rect -84 -71 84 -37
rect 174 -71 342 -37
rect 432 -71 600 -37
rect -662 -306 -628 -130
rect -404 -306 -370 -130
rect -146 -306 -112 -130
rect 112 -306 146 -130
rect 370 -306 404 -130
rect 628 -306 662 -130
rect -600 -399 -432 -365
rect -342 -399 -174 -365
rect -84 -399 84 -365
rect 174 -399 342 -365
rect 432 -399 600 -365
<< metal1 >>
rect -612 399 -420 405
rect -612 365 -600 399
rect -432 365 -420 399
rect -612 359 -420 365
rect -354 399 -162 405
rect -354 365 -342 399
rect -174 365 -162 399
rect -354 359 -162 365
rect -96 399 96 405
rect -96 365 -84 399
rect 84 365 96 399
rect -96 359 96 365
rect 162 399 354 405
rect 162 365 174 399
rect 342 365 354 399
rect 162 359 354 365
rect 420 399 612 405
rect 420 365 432 399
rect 600 365 612 399
rect 420 359 612 365
rect -668 306 -622 318
rect -668 130 -662 306
rect -628 130 -622 306
rect -668 118 -622 130
rect -410 306 -364 318
rect -410 130 -404 306
rect -370 130 -364 306
rect -410 118 -364 130
rect -152 306 -106 318
rect -152 130 -146 306
rect -112 130 -106 306
rect -152 118 -106 130
rect 106 306 152 318
rect 106 130 112 306
rect 146 130 152 306
rect 106 118 152 130
rect 364 306 410 318
rect 364 130 370 306
rect 404 130 410 306
rect 364 118 410 130
rect 622 306 668 318
rect 622 130 628 306
rect 662 130 668 306
rect 622 118 668 130
rect -612 71 -420 77
rect -612 37 -600 71
rect -432 37 -420 71
rect -612 31 -420 37
rect -354 71 -162 77
rect -354 37 -342 71
rect -174 37 -162 71
rect -354 31 -162 37
rect -96 71 96 77
rect -96 37 -84 71
rect 84 37 96 71
rect -96 31 96 37
rect 162 71 354 77
rect 162 37 174 71
rect 342 37 354 71
rect 162 31 354 37
rect 420 71 612 77
rect 420 37 432 71
rect 600 37 612 71
rect 420 31 612 37
rect -612 -37 -420 -31
rect -612 -71 -600 -37
rect -432 -71 -420 -37
rect -612 -77 -420 -71
rect -354 -37 -162 -31
rect -354 -71 -342 -37
rect -174 -71 -162 -37
rect -354 -77 -162 -71
rect -96 -37 96 -31
rect -96 -71 -84 -37
rect 84 -71 96 -37
rect -96 -77 96 -71
rect 162 -37 354 -31
rect 162 -71 174 -37
rect 342 -71 354 -37
rect 162 -77 354 -71
rect 420 -37 612 -31
rect 420 -71 432 -37
rect 600 -71 612 -37
rect 420 -77 612 -71
rect -668 -130 -622 -118
rect -668 -306 -662 -130
rect -628 -306 -622 -130
rect -668 -318 -622 -306
rect -410 -130 -364 -118
rect -410 -306 -404 -130
rect -370 -306 -364 -130
rect -410 -318 -364 -306
rect -152 -130 -106 -118
rect -152 -306 -146 -130
rect -112 -306 -106 -130
rect -152 -318 -106 -306
rect 106 -130 152 -118
rect 106 -306 112 -130
rect 146 -306 152 -130
rect 106 -318 152 -306
rect 364 -130 410 -118
rect 364 -306 370 -130
rect 404 -306 410 -130
rect 364 -318 410 -306
rect 622 -130 668 -118
rect 622 -306 628 -130
rect 662 -306 668 -130
rect 622 -318 668 -306
rect -612 -365 -420 -359
rect -612 -399 -600 -365
rect -432 -399 -420 -365
rect -612 -405 -420 -399
rect -354 -365 -162 -359
rect -354 -399 -342 -365
rect -174 -399 -162 -365
rect -354 -405 -162 -399
rect -96 -365 96 -359
rect -96 -399 -84 -365
rect 84 -399 96 -365
rect -96 -405 96 -399
rect 162 -365 354 -359
rect 162 -399 174 -365
rect 342 -399 354 -365
rect 162 -405 354 -399
rect 420 -365 612 -359
rect 420 -399 432 -365
rect 600 -399 612 -365
rect 420 -405 612 -399
<< properties >>
string FIXED_BBOX -759 -484 759 484
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 1 m 2 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
