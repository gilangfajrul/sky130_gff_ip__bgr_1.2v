magic
tech sky130A
magscale 1 2
timestamp 1720284156
<< xpolycontact >>
rect -450 1352 -380 1784
rect -450 52 -380 484
rect -284 1352 -214 1784
rect -284 52 -214 484
rect -118 1352 -48 1784
rect -118 52 -48 484
rect 48 1352 118 1784
rect 48 52 118 484
rect 214 1352 284 1784
rect 214 52 284 484
rect 380 1352 450 1784
rect 380 52 450 484
rect -450 -484 -380 -52
rect -450 -1784 -380 -1352
rect -284 -484 -214 -52
rect -284 -1784 -214 -1352
rect -118 -484 -48 -52
rect -118 -1784 -48 -1352
rect 48 -484 118 -52
rect 48 -1784 118 -1352
rect 214 -484 284 -52
rect 214 -1784 284 -1352
rect 380 -484 450 -52
rect 380 -1784 450 -1352
<< ppolyres >>
rect -450 484 -380 1352
rect -284 484 -214 1352
rect -118 484 -48 1352
rect 48 484 118 1352
rect 214 484 284 1352
rect 380 484 450 1352
rect -450 -1352 -380 -484
rect -284 -1352 -214 -484
rect -118 -1352 -48 -484
rect 48 -1352 118 -484
rect 214 -1352 284 -484
rect 380 -1352 450 -484
<< viali >>
rect -434 1369 -396 1766
rect -268 1369 -230 1766
rect -102 1369 -64 1766
rect 64 1369 102 1766
rect 230 1369 268 1766
rect 396 1369 434 1766
rect -434 70 -396 467
rect -268 70 -230 467
rect -102 70 -64 467
rect 64 70 102 467
rect 230 70 268 467
rect 396 70 434 467
rect -434 -467 -396 -70
rect -268 -467 -230 -70
rect -102 -467 -64 -70
rect 64 -467 102 -70
rect 230 -467 268 -70
rect 396 -467 434 -70
rect -434 -1766 -396 -1369
rect -268 -1766 -230 -1369
rect -102 -1766 -64 -1369
rect 64 -1766 102 -1369
rect 230 -1766 268 -1369
rect 396 -1766 434 -1369
<< metal1 >>
rect -440 1766 -390 1778
rect -440 1369 -434 1766
rect -396 1369 -390 1766
rect -440 1357 -390 1369
rect -274 1766 -224 1778
rect -274 1369 -268 1766
rect -230 1369 -224 1766
rect -274 1357 -224 1369
rect -108 1766 -58 1778
rect -108 1369 -102 1766
rect -64 1369 -58 1766
rect -108 1357 -58 1369
rect 58 1766 108 1778
rect 58 1369 64 1766
rect 102 1369 108 1766
rect 58 1357 108 1369
rect 224 1766 274 1778
rect 224 1369 230 1766
rect 268 1369 274 1766
rect 224 1357 274 1369
rect 390 1766 440 1778
rect 390 1369 396 1766
rect 434 1369 440 1766
rect 390 1357 440 1369
rect -440 467 -390 479
rect -440 70 -434 467
rect -396 70 -390 467
rect -440 58 -390 70
rect -274 467 -224 479
rect -274 70 -268 467
rect -230 70 -224 467
rect -274 58 -224 70
rect -108 467 -58 479
rect -108 70 -102 467
rect -64 70 -58 467
rect -108 58 -58 70
rect 58 467 108 479
rect 58 70 64 467
rect 102 70 108 467
rect 58 58 108 70
rect 224 467 274 479
rect 224 70 230 467
rect 268 70 274 467
rect 224 58 274 70
rect 390 467 440 479
rect 390 70 396 467
rect 434 70 440 467
rect 390 58 440 70
rect -440 -70 -390 -58
rect -440 -467 -434 -70
rect -396 -467 -390 -70
rect -440 -479 -390 -467
rect -274 -70 -224 -58
rect -274 -467 -268 -70
rect -230 -467 -224 -70
rect -274 -479 -224 -467
rect -108 -70 -58 -58
rect -108 -467 -102 -70
rect -64 -467 -58 -70
rect -108 -479 -58 -467
rect 58 -70 108 -58
rect 58 -467 64 -70
rect 102 -467 108 -70
rect 58 -479 108 -467
rect 224 -70 274 -58
rect 224 -467 230 -70
rect 268 -467 274 -70
rect 224 -479 274 -467
rect 390 -70 440 -58
rect 390 -467 396 -70
rect 434 -467 440 -70
rect 390 -479 440 -467
rect -440 -1369 -390 -1357
rect -440 -1766 -434 -1369
rect -396 -1766 -390 -1369
rect -440 -1778 -390 -1766
rect -274 -1369 -224 -1357
rect -274 -1766 -268 -1369
rect -230 -1766 -224 -1369
rect -274 -1778 -224 -1766
rect -108 -1369 -58 -1357
rect -108 -1766 -102 -1369
rect -64 -1766 -58 -1369
rect -108 -1778 -58 -1766
rect 58 -1369 108 -1357
rect 58 -1766 64 -1369
rect 102 -1766 108 -1369
rect 58 -1778 108 -1766
rect 224 -1369 274 -1357
rect 224 -1766 230 -1369
rect 268 -1766 274 -1369
rect 224 -1778 274 -1766
rect 390 -1369 440 -1357
rect 390 -1766 396 -1369
rect 434 -1766 440 -1369
rect 390 -1778 440 -1766
<< properties >>
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.350 l 4.5 m 2 nx 6 wmin 0.350 lmin 0.50 rho 319.8 val 5.224k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
