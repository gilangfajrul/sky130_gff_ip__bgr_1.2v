magic
tech sky130A
magscale 1 2
timestamp 1764413320
<< viali >>
rect 41 7178 1299 7250
rect 41 6064 113 7178
rect 189 7031 1151 7103
rect 189 6213 261 7031
rect 1079 6213 1151 7031
rect 189 6141 1151 6213
rect 1227 6064 1299 7178
rect 41 5992 1299 6064
rect 1529 7178 2787 7250
rect 1529 6064 1601 7178
rect 1677 7031 2639 7103
rect 1677 6213 1749 7031
rect 2567 6213 2639 7031
rect 1677 6141 2639 6213
rect 2715 6064 2787 7178
rect 1529 5992 2787 6064
rect 3017 7178 4275 7250
rect 3017 6064 3089 7178
rect 3165 7031 4127 7103
rect 3165 6213 3237 7031
rect 4055 6213 4127 7031
rect 3165 6141 4127 6213
rect 4203 6064 4275 7178
rect 3017 5992 4275 6064
rect 4505 7178 5763 7250
rect 4505 6064 4577 7178
rect 4653 7031 5615 7103
rect 4653 6213 4725 7031
rect 5543 6213 5615 7031
rect 4653 6141 5615 6213
rect 5691 6064 5763 7178
rect 4505 5992 5763 6064
rect 5993 7178 7251 7250
rect 5993 6064 6065 7178
rect 6141 7031 7103 7103
rect 6141 6213 6213 7031
rect 7031 6213 7103 7031
rect 6141 6141 7103 6213
rect 7179 6064 7251 7178
rect 5993 5992 7251 6064
rect 41 5690 1299 5762
rect 41 4576 113 5690
rect 189 5543 1151 5615
rect 189 4725 261 5543
rect 1079 4725 1151 5543
rect 189 4653 1151 4725
rect 1227 4576 1299 5690
rect 41 4504 1299 4576
rect 1529 5690 2787 5762
rect 1529 4576 1601 5690
rect 1677 5543 2639 5615
rect 1677 4725 1749 5543
rect 2567 4725 2639 5543
rect 1677 4653 2639 4725
rect 2715 4576 2787 5690
rect 1529 4504 2787 4576
rect 3017 5690 4275 5762
rect 3017 4576 3089 5690
rect 3165 5543 4127 5615
rect 3165 4725 3237 5543
rect 4055 4725 4127 5543
rect 3165 4653 4127 4725
rect 4203 4576 4275 5690
rect 3017 4504 4275 4576
rect 4505 5690 5763 5762
rect 4505 4576 4577 5690
rect 4653 5543 5615 5615
rect 4653 4725 4725 5543
rect 5543 4725 5615 5543
rect 4653 4653 5615 4725
rect 5691 4576 5763 5690
rect 4505 4504 5763 4576
rect 5993 5690 7251 5762
rect 5993 4576 6065 5690
rect 6141 5543 7103 5615
rect 6141 4725 6213 5543
rect 7031 4725 7103 5543
rect 6141 4653 7103 4725
rect 7179 4576 7251 5690
rect 5993 4504 7251 4576
rect 41 4202 1299 4274
rect 41 3088 113 4202
rect 189 4055 1151 4127
rect 189 3237 261 4055
rect 1079 3237 1151 4055
rect 189 3165 1151 3237
rect 1227 3088 1299 4202
rect 41 3016 1299 3088
rect 1529 4202 2787 4274
rect 1529 3088 1601 4202
rect 1677 4055 2639 4127
rect 1677 3237 1749 4055
rect 2567 3237 2639 4055
rect 1677 3165 2639 3237
rect 2715 3088 2787 4202
rect 1529 3016 2787 3088
rect 3017 4202 4275 4274
rect 3017 3088 3089 4202
rect 3165 4055 4127 4127
rect 3165 3237 3237 4055
rect 4055 3237 4127 4055
rect 3165 3165 4127 3237
rect 4203 3088 4275 4202
rect 3017 3016 4275 3088
rect 4505 4202 5763 4274
rect 4505 3088 4577 4202
rect 4653 4055 5615 4127
rect 4653 3237 4725 4055
rect 5543 3237 5615 4055
rect 4653 3165 5615 3237
rect 5691 3088 5763 4202
rect 4505 3016 5763 3088
rect 5993 4202 7251 4274
rect 5993 3088 6065 4202
rect 6141 4055 7103 4127
rect 6141 3237 6213 4055
rect 7031 3237 7103 4055
rect 6141 3165 7103 3237
rect 7179 3088 7251 4202
rect 5993 3016 7251 3088
rect 41 2714 1299 2786
rect 41 1600 113 2714
rect 189 2567 1151 2639
rect 189 1749 261 2567
rect 1079 1749 1151 2567
rect 189 1677 1151 1749
rect 1227 1600 1299 2714
rect 41 1528 1299 1600
rect 1529 2714 2787 2786
rect 1529 1600 1601 2714
rect 1677 2567 2639 2639
rect 1677 1749 1749 2567
rect 2567 1749 2639 2567
rect 1677 1677 2639 1749
rect 2715 1600 2787 2714
rect 1529 1528 2787 1600
rect 3017 2714 4275 2786
rect 3017 1600 3089 2714
rect 3165 2567 4127 2639
rect 3165 1749 3237 2567
rect 4055 1749 4127 2567
rect 3165 1677 4127 1749
rect 4203 1600 4275 2714
rect 3017 1528 4275 1600
rect 4505 2714 5763 2786
rect 4505 1600 4577 2714
rect 4653 2567 5615 2639
rect 4653 1749 4725 2567
rect 5543 1749 5615 2567
rect 4653 1677 5615 1749
rect 5691 1600 5763 2714
rect 4505 1528 5763 1600
rect 5993 2714 7251 2786
rect 5993 1600 6065 2714
rect 6141 2567 7103 2639
rect 6141 1749 6213 2567
rect 7031 1749 7103 2567
rect 6141 1677 7103 1749
rect 7179 1600 7251 2714
rect 5993 1528 7251 1600
rect 41 1226 1299 1298
rect 41 112 113 1226
rect 189 1079 1151 1151
rect 189 261 261 1079
rect 1079 261 1151 1079
rect 189 189 1151 261
rect 1227 112 1299 1226
rect 41 40 1299 112
rect 1529 1226 2787 1298
rect 1529 112 1601 1226
rect 1677 1079 2639 1151
rect 1677 261 1749 1079
rect 2567 261 2639 1079
rect 1677 189 2639 261
rect 2715 112 2787 1226
rect 1529 40 2787 112
rect 3017 1226 4275 1298
rect 3017 112 3089 1226
rect 3165 1079 4127 1151
rect 3165 261 3237 1079
rect 4055 261 4127 1079
rect 3165 189 4127 261
rect 4203 112 4275 1226
rect 3017 40 4275 112
rect 4505 1226 5763 1298
rect 4505 112 4577 1226
rect 4653 1079 5615 1151
rect 4653 261 4725 1079
rect 5543 261 5615 1079
rect 4653 189 5615 261
rect 5691 112 5763 1226
rect 4505 40 5763 112
rect 5993 1226 7251 1298
rect 5993 112 6065 1226
rect 6141 1079 7103 1151
rect 6141 261 6213 1079
rect 7031 261 7103 1079
rect 6141 189 7103 261
rect 7179 112 7251 1226
rect 5993 40 7251 112
<< metal1 >>
rect 35 7256 119 7262
rect 1221 7256 1305 7262
rect 1523 7256 1607 7262
rect 2709 7256 2793 7262
rect 3011 7256 3095 7262
rect 4197 7256 4281 7262
rect 4499 7256 4583 7262
rect 5685 7256 5769 7262
rect 5987 7256 6071 7262
rect 7173 7256 7257 7262
rect 29 7250 1311 7256
rect 29 7172 41 7250
rect 35 6070 41 7172
rect 29 5992 41 6070
rect 113 7172 1227 7178
rect 113 6070 119 7172
rect 183 7109 267 7115
rect 1073 7109 1157 7115
rect 177 7103 1163 7109
rect 177 7025 189 7103
rect 183 6219 189 7025
rect 177 6141 189 6219
rect 261 7025 1079 7031
rect 261 6219 267 7025
rect 1073 6673 1079 7025
rect 364 6573 1079 6673
rect 620 6219 720 6573
rect 1073 6219 1079 6573
rect 261 6213 1079 6219
rect 1151 7025 1163 7103
rect 1151 6673 1157 7025
rect 1221 6673 1227 7172
rect 1151 6573 1227 6673
rect 1151 6219 1157 6573
rect 1151 6141 1163 6219
rect 177 6135 1163 6141
rect 183 6129 267 6135
rect 620 6070 720 6135
rect 1073 6129 1157 6135
rect 1221 6070 1227 6573
rect 113 6064 1227 6070
rect 1299 7172 1311 7250
rect 1517 7250 2799 7256
rect 1517 7172 1529 7250
rect 1299 6673 1305 7172
rect 1523 6673 1529 7172
rect 1299 6573 1529 6673
rect 1299 6070 1305 6573
rect 1523 6070 1529 6573
rect 1299 5992 1311 6070
rect 29 5986 1311 5992
rect 1517 5992 1529 6070
rect 1601 7172 2715 7178
rect 1601 6673 1607 7172
rect 1671 7109 1755 7115
rect 2561 7109 2645 7115
rect 1665 7103 2651 7109
rect 1665 7025 1677 7103
rect 1671 6673 1677 7025
rect 1601 6573 1677 6673
rect 1601 6070 1607 6573
rect 1671 6219 1677 6573
rect 1665 6141 1677 6219
rect 1749 7025 2567 7031
rect 1749 6673 1755 7025
rect 2561 6673 2567 7025
rect 1749 6573 2567 6673
rect 1749 6219 1755 6573
rect 2561 6219 2567 6573
rect 1749 6213 2567 6219
rect 2639 7025 2651 7103
rect 2639 6673 2645 7025
rect 2709 6673 2715 7172
rect 2639 6573 2715 6673
rect 2639 6219 2645 6573
rect 2639 6141 2651 6219
rect 1665 6135 2651 6141
rect 1671 6129 1755 6135
rect 2561 6129 2645 6135
rect 2709 6070 2715 6573
rect 1601 6064 2715 6070
rect 2787 7172 2799 7250
rect 3005 7250 4287 7256
rect 3005 7172 3017 7250
rect 2787 6673 2793 7172
rect 3011 6673 3017 7172
rect 2787 6573 3017 6673
rect 2787 6070 2793 6573
rect 3011 6070 3017 6573
rect 2787 5992 2799 6070
rect 1517 5986 2799 5992
rect 3005 5992 3017 6070
rect 3089 7172 4203 7178
rect 3089 6673 3095 7172
rect 3159 7109 3243 7115
rect 4049 7109 4133 7115
rect 3153 7103 4139 7109
rect 3153 7025 3165 7103
rect 3159 6673 3165 7025
rect 3089 6573 3165 6673
rect 3089 6070 3095 6573
rect 3159 6219 3165 6573
rect 3153 6141 3165 6219
rect 3237 7025 4055 7031
rect 3237 6673 3243 7025
rect 4049 6673 4055 7025
rect 3237 6573 4055 6673
rect 3237 6219 3243 6573
rect 4049 6219 4055 6573
rect 3237 6213 4055 6219
rect 4127 7025 4139 7103
rect 4127 6673 4133 7025
rect 4197 6673 4203 7172
rect 4127 6573 4203 6673
rect 4127 6219 4133 6573
rect 4127 6141 4139 6219
rect 3153 6135 4139 6141
rect 3159 6129 3243 6135
rect 4049 6129 4133 6135
rect 4197 6070 4203 6573
rect 3089 6064 4203 6070
rect 4275 7172 4287 7250
rect 4493 7250 5775 7256
rect 4493 7172 4505 7250
rect 4275 6673 4281 7172
rect 4499 6673 4505 7172
rect 4275 6573 4505 6673
rect 4275 6070 4281 6573
rect 4499 6070 4505 6573
rect 4275 5992 4287 6070
rect 3005 5986 4287 5992
rect 4493 5992 4505 6070
rect 4577 7172 5691 7178
rect 4577 6673 4583 7172
rect 4647 7109 4731 7115
rect 5537 7109 5621 7115
rect 4641 7103 5627 7109
rect 4641 7025 4653 7103
rect 4647 6673 4653 7025
rect 4577 6573 4653 6673
rect 4577 6070 4583 6573
rect 4647 6219 4653 6573
rect 4641 6141 4653 6219
rect 4725 7025 5543 7031
rect 4725 6673 4731 7025
rect 5537 6673 5543 7025
rect 4725 6573 5543 6673
rect 4725 6219 4731 6573
rect 5537 6219 5543 6573
rect 4725 6213 5543 6219
rect 5615 7025 5627 7103
rect 5615 6673 5621 7025
rect 5685 6673 5691 7172
rect 5615 6573 5691 6673
rect 5615 6219 5621 6573
rect 5615 6141 5627 6219
rect 4641 6135 5627 6141
rect 4647 6129 4731 6135
rect 5537 6129 5621 6135
rect 5685 6070 5691 6573
rect 4577 6064 5691 6070
rect 5763 7172 5775 7250
rect 5981 7250 7263 7256
rect 5981 7172 5993 7250
rect 5763 6673 5769 7172
rect 5987 6673 5993 7172
rect 5763 6573 5993 6673
rect 5763 6070 5769 6573
rect 5987 6070 5993 6573
rect 5763 5992 5775 6070
rect 4493 5986 5775 5992
rect 5981 5992 5993 6070
rect 6065 7172 7179 7178
rect 6065 6673 6071 7172
rect 6135 7109 6219 7115
rect 7025 7109 7109 7115
rect 6129 7103 7115 7109
rect 6129 7025 6141 7103
rect 6135 6673 6141 7025
rect 6065 6573 6141 6673
rect 6065 6070 6071 6573
rect 6135 6219 6141 6573
rect 6129 6141 6141 6219
rect 6213 7025 7031 7031
rect 6213 6673 6219 7025
rect 6213 6573 6672 6673
rect 6213 6219 6219 6573
rect 6572 6219 6672 6573
rect 7025 6219 7031 7025
rect 6213 6213 7031 6219
rect 7103 7025 7115 7103
rect 7103 6219 7109 7025
rect 7103 6141 7115 6219
rect 6129 6135 7115 6141
rect 6135 6129 6219 6135
rect 6572 6070 6672 6135
rect 7025 6129 7109 6135
rect 7173 6070 7179 7172
rect 6065 6064 7179 6070
rect 7251 7172 7263 7250
rect 7251 6070 7257 7172
rect 7251 5992 7263 6070
rect 5981 5986 7263 5992
rect 35 5980 119 5986
rect 35 5768 119 5774
rect 620 5768 720 5986
rect 1221 5980 1305 5986
rect 1523 5980 1607 5986
rect 2709 5980 2793 5986
rect 3011 5980 3095 5986
rect 4197 5980 4281 5986
rect 4499 5980 4583 5986
rect 5685 5980 5769 5986
rect 5987 5980 6071 5986
rect 1221 5768 1305 5774
rect 1523 5768 1607 5774
rect 2709 5768 2793 5774
rect 3011 5768 3095 5774
rect 4197 5768 4281 5774
rect 4499 5768 4583 5774
rect 5685 5768 5769 5774
rect 5987 5768 6071 5774
rect 6572 5768 6672 5986
rect 7173 5980 7257 5986
rect 7173 5768 7257 5774
rect 29 5762 1311 5768
rect 29 5684 41 5762
rect 35 4582 41 5684
rect 29 4504 41 4582
rect 113 5684 1227 5690
rect 113 4582 119 5684
rect 183 5621 267 5627
rect 620 5621 720 5684
rect 1221 5627 1227 5684
rect 1073 5621 1227 5627
rect 177 5615 1227 5621
rect 177 5537 189 5615
rect 183 4731 189 5537
rect 177 4653 189 4731
rect 261 5537 1079 5543
rect 261 4731 267 5537
rect 620 4731 720 5537
rect 1073 4731 1079 5537
rect 261 4725 1079 4731
rect 1151 5527 1227 5615
rect 1151 4741 1157 5527
rect 1221 4741 1227 5527
rect 1151 4653 1227 4741
rect 177 4647 1227 4653
rect 183 4641 267 4647
rect 620 4582 720 4647
rect 1073 4641 1227 4647
rect 1221 4582 1227 4641
rect 113 4576 1227 4582
rect 1299 5684 1311 5762
rect 1517 5762 2799 5768
rect 1517 5684 1529 5762
rect 1299 5627 1305 5684
rect 1523 5627 1529 5684
rect 1299 5527 1529 5627
rect 1299 4741 1305 5527
rect 1523 4741 1529 5527
rect 1299 4641 1529 4741
rect 1299 4582 1305 4641
rect 1523 4582 1529 4641
rect 1299 4504 1311 4582
rect 29 4498 1311 4504
rect 1517 4504 1529 4582
rect 1601 5684 2715 5690
rect 1601 5627 1607 5684
rect 2709 5627 2715 5684
rect 1601 5615 2715 5627
rect 1601 5527 1677 5615
rect 1601 4741 1607 5527
rect 1671 4741 1677 5527
rect 1601 4653 1677 4741
rect 1749 5527 2567 5543
rect 1749 4741 1755 5527
rect 1843 4829 1853 5439
rect 2463 4829 2473 5439
rect 2561 4741 2567 5527
rect 1749 4725 2567 4741
rect 2639 5527 2715 5615
rect 2639 4741 2645 5527
rect 2709 4741 2715 5527
rect 2639 4653 2715 4741
rect 1601 4641 2715 4653
rect 1601 4582 1607 4641
rect 2709 4582 2715 4641
rect 1601 4576 2715 4582
rect 2787 5684 2799 5762
rect 3005 5762 4287 5768
rect 3005 5684 3017 5762
rect 2787 5627 2793 5684
rect 3011 5627 3017 5684
rect 2787 5527 3017 5627
rect 2787 4741 2793 5527
rect 3011 4741 3017 5527
rect 2787 4641 3017 4741
rect 2787 4582 2793 4641
rect 3011 4582 3017 4641
rect 2787 4504 2799 4582
rect 1517 4498 2799 4504
rect 3005 4504 3017 4582
rect 3089 5684 4203 5690
rect 3089 5627 3095 5684
rect 4197 5627 4203 5684
rect 3089 5615 4203 5627
rect 3089 5527 3165 5615
rect 3089 4741 3095 5527
rect 3159 4741 3165 5527
rect 3089 4653 3165 4741
rect 3237 5527 4055 5543
rect 3237 4741 3243 5527
rect 3331 4829 3341 5439
rect 3951 4829 3961 5439
rect 4049 4741 4055 5527
rect 3237 4725 4055 4741
rect 4127 5527 4203 5615
rect 4127 4741 4133 5527
rect 4197 4741 4203 5527
rect 4127 4653 4203 4741
rect 3089 4641 4203 4653
rect 3089 4582 3095 4641
rect 4197 4582 4203 4641
rect 3089 4576 4203 4582
rect 4275 5684 4287 5762
rect 4493 5762 5775 5768
rect 4493 5684 4505 5762
rect 4275 5627 4281 5684
rect 4499 5627 4505 5684
rect 4275 5527 4505 5627
rect 4275 4741 4281 5527
rect 4499 4741 4505 5527
rect 4275 4641 4505 4741
rect 4275 4582 4281 4641
rect 4499 4582 4505 4641
rect 4275 4504 4287 4582
rect 3005 4498 4287 4504
rect 4493 4504 4505 4582
rect 4577 5684 5691 5690
rect 4577 5627 4583 5684
rect 5685 5627 5691 5684
rect 4577 5615 5691 5627
rect 4577 5527 4653 5615
rect 4577 4741 4583 5527
rect 4647 4741 4653 5527
rect 4577 4653 4653 4741
rect 4725 5527 5543 5543
rect 4725 4741 4731 5527
rect 4819 4829 4829 5439
rect 5439 4829 5449 5439
rect 5537 4741 5543 5527
rect 4725 4725 5543 4741
rect 5615 5527 5691 5615
rect 5615 4741 5621 5527
rect 5685 4741 5691 5527
rect 5615 4653 5691 4741
rect 4577 4641 5691 4653
rect 4577 4582 4583 4641
rect 5685 4582 5691 4641
rect 4577 4576 5691 4582
rect 5763 5684 5775 5762
rect 5981 5762 7263 5768
rect 5981 5684 5993 5762
rect 5763 5627 5769 5684
rect 5987 5627 5993 5684
rect 5763 5527 5993 5627
rect 5763 4741 5769 5527
rect 5987 4741 5993 5527
rect 5763 4641 5993 4741
rect 5763 4582 5769 4641
rect 5987 4582 5993 4641
rect 5763 4504 5775 4582
rect 4493 4498 5775 4504
rect 5981 4504 5993 4582
rect 6065 5684 7179 5690
rect 6065 5627 6071 5684
rect 6065 5621 6219 5627
rect 6572 5621 6672 5684
rect 7025 5621 7109 5627
rect 6065 5615 7115 5621
rect 6065 5527 6141 5615
rect 6065 4741 6071 5527
rect 6135 4741 6141 5527
rect 6065 4653 6141 4741
rect 6213 5537 7031 5543
rect 6213 4731 6219 5537
rect 6572 4731 6672 5537
rect 7025 4731 7031 5537
rect 6213 4725 7031 4731
rect 7103 5537 7115 5615
rect 7103 4731 7109 5537
rect 7103 4653 7115 4731
rect 6065 4647 7115 4653
rect 6065 4641 6219 4647
rect 6065 4582 6071 4641
rect 6572 4582 6672 4647
rect 7025 4641 7109 4647
rect 7173 4582 7179 5684
rect 6065 4576 7179 4582
rect 7251 5684 7263 5762
rect 7251 4582 7257 5684
rect 7251 4504 7263 4582
rect 5981 4498 7263 4504
rect 35 4492 119 4498
rect 35 4280 119 4286
rect 620 4280 720 4498
rect 1221 4492 1305 4498
rect 1523 4492 1607 4498
rect 2709 4492 2793 4498
rect 3011 4492 3095 4498
rect 4197 4492 4281 4498
rect 4499 4492 4583 4498
rect 5685 4492 5769 4498
rect 5987 4492 6071 4498
rect 1221 4280 1305 4286
rect 1523 4280 1607 4286
rect 2709 4280 2793 4286
rect 3011 4280 3095 4286
rect 4197 4280 4281 4286
rect 4499 4280 4583 4286
rect 5685 4280 5769 4286
rect 5987 4280 6071 4286
rect 6572 4280 6672 4498
rect 7173 4492 7257 4498
rect 7173 4280 7257 4286
rect 29 4274 1311 4280
rect 29 4196 41 4274
rect 35 3094 41 4196
rect 29 3016 41 3094
rect 113 4196 1227 4202
rect 113 3094 119 4196
rect 183 4133 267 4139
rect 620 4133 720 4196
rect 1221 4139 1227 4196
rect 1073 4133 1227 4139
rect 177 4127 1227 4133
rect 177 4049 189 4127
rect 183 3243 189 4049
rect 177 3165 189 3243
rect 261 4049 1079 4055
rect 261 3243 267 4049
rect 620 3243 720 4049
rect 1073 3243 1079 4049
rect 261 3237 1079 3243
rect 1151 4039 1227 4127
rect 1151 3253 1157 4039
rect 1221 3253 1227 4039
rect 1151 3165 1227 3253
rect 177 3159 1227 3165
rect 183 3153 267 3159
rect 620 3094 720 3159
rect 1073 3153 1227 3159
rect 1221 3094 1227 3153
rect 113 3088 1227 3094
rect 1299 4196 1311 4274
rect 1517 4274 2799 4280
rect 1517 4196 1529 4274
rect 1299 4139 1305 4196
rect 1523 4139 1529 4196
rect 1299 4039 1529 4139
rect 1299 3253 1305 4039
rect 1523 3253 1529 4039
rect 1299 3153 1529 3253
rect 1299 3094 1305 3153
rect 1523 3094 1529 3153
rect 1299 3016 1311 3094
rect 29 3010 1311 3016
rect 1517 3016 1529 3094
rect 1601 4196 2715 4202
rect 1601 4139 1607 4196
rect 2709 4139 2715 4196
rect 1601 4127 2715 4139
rect 1601 4039 1677 4127
rect 1601 3253 1607 4039
rect 1671 3253 1677 4039
rect 1601 3165 1677 3253
rect 1749 4039 2567 4055
rect 1749 3253 1755 4039
rect 1843 3341 1853 3951
rect 2463 3341 2473 3951
rect 2561 3253 2567 4039
rect 1749 3237 2567 3253
rect 2639 4039 2715 4127
rect 2639 3253 2645 4039
rect 2709 3253 2715 4039
rect 2639 3165 2715 3253
rect 1601 3153 2715 3165
rect 1601 3094 1607 3153
rect 2709 3094 2715 3153
rect 1601 3088 2715 3094
rect 2787 4196 2799 4274
rect 3005 4274 4287 4280
rect 3005 4196 3017 4274
rect 2787 4139 2793 4196
rect 3011 4139 3017 4196
rect 2787 4039 3017 4139
rect 2787 3253 2793 4039
rect 3011 3253 3017 4039
rect 2787 3153 3017 3253
rect 2787 3094 2793 3153
rect 3011 3094 3017 3153
rect 2787 3016 2799 3094
rect 1517 3010 2799 3016
rect 3005 3016 3017 3094
rect 3089 4196 4203 4202
rect 3089 4139 3095 4196
rect 4197 4139 4203 4196
rect 3089 4127 4203 4139
rect 3089 4039 3165 4127
rect 3089 3253 3095 4039
rect 3159 3253 3165 4039
rect 3089 3165 3165 3253
rect 3237 4039 4055 4055
rect 3237 3253 3243 4039
rect 3331 3341 3341 3951
rect 3951 3341 3961 3951
rect 4049 3253 4055 4039
rect 3237 3237 4055 3253
rect 4127 4039 4203 4127
rect 4127 3253 4133 4039
rect 4197 3253 4203 4039
rect 4127 3165 4203 3253
rect 3089 3153 4203 3165
rect 3089 3094 3095 3153
rect 4197 3094 4203 3153
rect 3089 3088 4203 3094
rect 4275 4196 4287 4274
rect 4493 4274 5775 4280
rect 4493 4196 4505 4274
rect 4275 4139 4281 4196
rect 4499 4139 4505 4196
rect 4275 4039 4505 4139
rect 4275 3253 4281 4039
rect 4499 3253 4505 4039
rect 4275 3153 4505 3253
rect 4275 3094 4281 3153
rect 4499 3094 4505 3153
rect 4275 3016 4287 3094
rect 3005 3010 4287 3016
rect 4493 3016 4505 3094
rect 4577 4196 5691 4202
rect 4577 4139 4583 4196
rect 5685 4139 5691 4196
rect 4577 4127 5691 4139
rect 4577 4039 4653 4127
rect 4577 3253 4583 4039
rect 4647 3253 4653 4039
rect 4577 3165 4653 3253
rect 4725 4039 5543 4055
rect 4725 3253 4731 4039
rect 4819 3735 4829 3951
rect 5439 3735 5449 3951
rect 4819 3341 4829 3557
rect 5439 3341 5449 3557
rect 5537 3253 5543 4039
rect 4725 3237 5543 3253
rect 5615 4039 5691 4127
rect 5615 3253 5621 4039
rect 5685 3253 5691 4039
rect 5615 3165 5691 3253
rect 4577 3153 5691 3165
rect 4577 3094 4583 3153
rect 5685 3094 5691 3153
rect 4577 3088 5691 3094
rect 5763 4196 5775 4274
rect 5981 4274 7263 4280
rect 5981 4196 5993 4274
rect 5763 4139 5769 4196
rect 5987 4139 5993 4196
rect 5763 4039 5993 4139
rect 5763 3253 5769 4039
rect 5987 3253 5993 4039
rect 5763 3153 5993 3253
rect 5763 3094 5769 3153
rect 5987 3094 5993 3153
rect 5763 3016 5775 3094
rect 4493 3010 5775 3016
rect 5981 3016 5993 3094
rect 6065 4196 7179 4202
rect 6065 4139 6071 4196
rect 6065 4133 6219 4139
rect 6572 4133 6672 4196
rect 7025 4133 7109 4139
rect 6065 4127 7115 4133
rect 6065 4039 6141 4127
rect 6065 3253 6071 4039
rect 6135 3253 6141 4039
rect 6065 3165 6141 3253
rect 6213 4049 7031 4055
rect 6213 3243 6219 4049
rect 6572 3243 6672 4049
rect 7025 3243 7031 4049
rect 6213 3237 7031 3243
rect 7103 4049 7115 4127
rect 7103 3243 7109 4049
rect 7103 3165 7115 3243
rect 6065 3159 7115 3165
rect 6065 3153 6219 3159
rect 6065 3094 6071 3153
rect 6572 3094 6672 3159
rect 7025 3153 7109 3159
rect 7173 3094 7179 4196
rect 6065 3088 7179 3094
rect 7251 4196 7263 4274
rect 7251 3094 7257 4196
rect 7251 3016 7263 3094
rect 5981 3010 7263 3016
rect 35 3004 119 3010
rect 35 2792 119 2798
rect 620 2792 720 3010
rect 1221 3004 1305 3010
rect 1523 3004 1607 3010
rect 2709 3004 2793 3010
rect 3011 3004 3095 3010
rect 4197 3004 4281 3010
rect 4499 3004 4583 3010
rect 5685 3004 5769 3010
rect 5987 3004 6071 3010
rect 1221 2792 1305 2798
rect 1523 2792 1607 2798
rect 2709 2792 2793 2798
rect 3011 2792 3095 2798
rect 4197 2792 4281 2798
rect 4499 2792 4583 2798
rect 5685 2792 5769 2798
rect 5987 2792 6071 2798
rect 6572 2792 6672 3010
rect 7173 3004 7257 3010
rect 7173 2792 7257 2798
rect 29 2786 1311 2792
rect 29 2708 41 2786
rect 35 1606 41 2708
rect 29 1528 41 1606
rect 113 2708 1227 2714
rect 113 1606 119 2708
rect 183 2645 267 2651
rect 620 2645 720 2708
rect 1221 2651 1227 2708
rect 1073 2645 1227 2651
rect 177 2639 1227 2645
rect 177 2561 189 2639
rect 183 1755 189 2561
rect 177 1677 189 1755
rect 261 2561 1079 2567
rect 261 1755 267 2561
rect 620 1755 720 2561
rect 1073 1755 1079 2561
rect 261 1749 1079 1755
rect 1151 2551 1227 2639
rect 1151 1765 1157 2551
rect 1221 1765 1227 2551
rect 1151 1677 1227 1765
rect 177 1671 1227 1677
rect 183 1665 267 1671
rect 620 1606 720 1671
rect 1073 1665 1227 1671
rect 1221 1606 1227 1665
rect 113 1600 1227 1606
rect 1299 2708 1311 2786
rect 1517 2786 2799 2792
rect 1517 2708 1529 2786
rect 1299 2651 1305 2708
rect 1523 2651 1529 2708
rect 1299 2551 1529 2651
rect 1299 1765 1305 2551
rect 1523 1765 1529 2551
rect 1299 1665 1529 1765
rect 1299 1606 1305 1665
rect 1523 1606 1529 1665
rect 1299 1528 1311 1606
rect 29 1522 1311 1528
rect 1517 1528 1529 1606
rect 1601 2708 2715 2714
rect 1601 2651 1607 2708
rect 2709 2651 2715 2708
rect 1601 2639 2715 2651
rect 1601 2551 1677 2639
rect 1601 1765 1607 2551
rect 1671 1765 1677 2551
rect 1601 1677 1677 1765
rect 1749 2551 2567 2567
rect 1749 1765 1755 2551
rect 1843 1853 1853 2463
rect 2463 1853 2473 2463
rect 2561 1765 2567 2551
rect 1749 1749 2567 1765
rect 2639 2551 2715 2639
rect 2639 1765 2645 2551
rect 2709 1765 2715 2551
rect 2639 1677 2715 1765
rect 1601 1665 2715 1677
rect 1601 1606 1607 1665
rect 2709 1606 2715 1665
rect 1601 1600 2715 1606
rect 2787 2708 2799 2786
rect 3005 2786 4287 2792
rect 3005 2708 3017 2786
rect 2787 2651 2793 2708
rect 3011 2651 3017 2708
rect 2787 2551 3017 2651
rect 2787 1765 2793 2551
rect 3011 1765 3017 2551
rect 2787 1665 3017 1765
rect 2787 1606 2793 1665
rect 3011 1606 3017 1665
rect 2787 1528 2799 1606
rect 1517 1522 2799 1528
rect 3005 1528 3017 1606
rect 3089 2708 4203 2714
rect 3089 2651 3095 2708
rect 4197 2651 4203 2708
rect 3089 2639 4203 2651
rect 3089 2551 3165 2639
rect 3089 1765 3095 2551
rect 3159 1765 3165 2551
rect 3089 1677 3165 1765
rect 3237 2551 4055 2567
rect 3237 1765 3243 2551
rect 3331 1853 3341 2463
rect 3951 1853 3961 2463
rect 4049 1765 4055 2551
rect 3237 1749 4055 1765
rect 4127 2551 4203 2639
rect 4127 1765 4133 2551
rect 4197 1765 4203 2551
rect 4127 1677 4203 1765
rect 3089 1665 4203 1677
rect 3089 1606 3095 1665
rect 4197 1606 4203 1665
rect 3089 1600 4203 1606
rect 4275 2708 4287 2786
rect 4493 2786 5775 2792
rect 4493 2708 4505 2786
rect 4275 2651 4281 2708
rect 4499 2651 4505 2708
rect 4275 2551 4505 2651
rect 4275 1765 4281 2551
rect 4499 1765 4505 2551
rect 4275 1665 4505 1765
rect 4275 1606 4281 1665
rect 4499 1606 4505 1665
rect 4275 1528 4287 1606
rect 3005 1522 4287 1528
rect 4493 1528 4505 1606
rect 4577 2708 5691 2714
rect 4577 2651 4583 2708
rect 5685 2651 5691 2708
rect 4577 2639 5691 2651
rect 4577 2551 4653 2639
rect 4577 1765 4583 2551
rect 4647 1765 4653 2551
rect 4577 1677 4653 1765
rect 4725 2551 5543 2567
rect 4725 1765 4731 2551
rect 4819 1853 4829 2463
rect 5439 1853 5449 2463
rect 5537 1765 5543 2551
rect 4725 1749 5543 1765
rect 5615 2551 5691 2639
rect 5615 1765 5621 2551
rect 5685 1765 5691 2551
rect 5615 1677 5691 1765
rect 4577 1665 5691 1677
rect 4577 1606 4583 1665
rect 5685 1606 5691 1665
rect 4577 1600 5691 1606
rect 5763 2708 5775 2786
rect 5981 2786 7263 2792
rect 5981 2708 5993 2786
rect 5763 2651 5769 2708
rect 5987 2651 5993 2708
rect 5763 2551 5993 2651
rect 5763 1765 5769 2551
rect 5987 1765 5993 2551
rect 5763 1665 5993 1765
rect 5763 1606 5769 1665
rect 5987 1606 5993 1665
rect 5763 1528 5775 1606
rect 4493 1522 5775 1528
rect 5981 1528 5993 1606
rect 6065 2708 7179 2714
rect 6065 2651 6071 2708
rect 6065 2645 6219 2651
rect 6572 2645 6672 2708
rect 7025 2645 7109 2651
rect 6065 2639 7115 2645
rect 6065 2551 6141 2639
rect 6065 1765 6071 2551
rect 6135 1765 6141 2551
rect 6065 1677 6141 1765
rect 6213 2561 7031 2567
rect 6213 1755 6219 2561
rect 6572 1755 6672 2561
rect 7025 1755 7031 2561
rect 6213 1749 7031 1755
rect 7103 2561 7115 2639
rect 7103 1755 7109 2561
rect 7103 1677 7115 1755
rect 6065 1671 7115 1677
rect 6065 1665 6219 1671
rect 6065 1606 6071 1665
rect 6572 1606 6672 1671
rect 7025 1665 7109 1671
rect 7173 1606 7179 2708
rect 6065 1600 7179 1606
rect 7251 2708 7263 2786
rect 7251 1606 7257 2708
rect 7251 1528 7263 1606
rect 5981 1522 7263 1528
rect 35 1516 119 1522
rect 35 1304 119 1310
rect 620 1304 720 1522
rect 1221 1516 1305 1522
rect 1523 1516 1607 1522
rect 2709 1516 2793 1522
rect 3011 1516 3095 1522
rect 4197 1516 4281 1522
rect 4499 1516 4583 1522
rect 5685 1516 5769 1522
rect 5987 1516 6071 1522
rect 1221 1304 1305 1310
rect 1523 1304 1607 1310
rect 2709 1304 2793 1310
rect 3011 1304 3095 1310
rect 4197 1304 4281 1310
rect 4499 1304 4583 1310
rect 5685 1304 5769 1310
rect 5987 1304 6071 1310
rect 6572 1304 6672 1522
rect 7173 1516 7257 1522
rect 7173 1304 7257 1310
rect 29 1298 1311 1304
rect 29 1220 41 1298
rect 35 118 41 1220
rect 29 40 41 118
rect 113 1220 1227 1226
rect 113 118 119 1220
rect 183 1157 267 1163
rect 620 1157 720 1220
rect 1221 1163 1227 1220
rect 1073 1157 1227 1163
rect 177 1151 1227 1157
rect 177 1073 189 1151
rect 183 267 189 1073
rect 177 189 189 267
rect 261 1073 1079 1079
rect 261 267 267 1073
rect 620 721 720 1073
rect 1073 721 1079 1073
rect 620 621 1079 721
rect 1073 267 1079 621
rect 261 261 1079 267
rect 1151 1063 1227 1151
rect 1151 721 1157 1063
rect 1221 721 1227 1063
rect 1151 621 1227 721
rect 1151 277 1157 621
rect 1221 277 1227 621
rect 1151 189 1227 277
rect 177 183 1227 189
rect 183 177 267 183
rect 1073 177 1227 183
rect 1221 118 1227 177
rect 113 112 1227 118
rect 1299 1220 1311 1298
rect 1517 1298 2799 1304
rect 1517 1220 1529 1298
rect 1299 1163 1305 1220
rect 1523 1163 1529 1220
rect 1299 1063 1529 1163
rect 1299 721 1305 1063
rect 1523 721 1529 1063
rect 1299 621 1529 721
rect 1299 277 1305 621
rect 1523 277 1529 621
rect 1299 177 1529 277
rect 1299 118 1305 177
rect 1523 118 1529 177
rect 1299 40 1311 118
rect 29 34 1311 40
rect 1517 40 1529 118
rect 1601 1220 2715 1226
rect 1601 1163 1607 1220
rect 2709 1163 2715 1220
rect 1601 1151 2715 1163
rect 1601 1063 1677 1151
rect 1601 721 1607 1063
rect 1671 721 1677 1063
rect 1601 621 1677 721
rect 1601 277 1607 621
rect 1671 277 1677 621
rect 1601 189 1677 277
rect 1749 1063 2567 1079
rect 1749 721 1755 1063
rect 2561 721 2567 1063
rect 1749 621 2567 721
rect 1749 277 1755 621
rect 2561 277 2567 621
rect 1749 261 2567 277
rect 2639 1063 2715 1151
rect 2639 721 2645 1063
rect 2709 721 2715 1063
rect 2639 621 2715 721
rect 2639 277 2645 621
rect 2709 277 2715 621
rect 2639 189 2715 277
rect 1601 177 2715 189
rect 1601 118 1607 177
rect 2709 118 2715 177
rect 1601 112 2715 118
rect 2787 1220 2799 1298
rect 3005 1298 4287 1304
rect 3005 1220 3017 1298
rect 2787 1163 2793 1220
rect 3011 1163 3017 1220
rect 2787 1063 3017 1163
rect 2787 721 2793 1063
rect 3011 721 3017 1063
rect 2787 621 3017 721
rect 2787 277 2793 621
rect 3011 277 3017 621
rect 2787 177 3017 277
rect 2787 118 2793 177
rect 3011 118 3017 177
rect 2787 40 2799 118
rect 1517 34 2799 40
rect 3005 40 3017 118
rect 3089 1220 4203 1226
rect 3089 1163 3095 1220
rect 4197 1163 4203 1220
rect 3089 1151 4203 1163
rect 3089 1063 3165 1151
rect 3089 721 3095 1063
rect 3159 721 3165 1063
rect 3089 621 3165 721
rect 3089 277 3095 621
rect 3159 277 3165 621
rect 3089 189 3165 277
rect 3237 1063 4055 1079
rect 3237 721 3243 1063
rect 4049 721 4055 1063
rect 3237 621 4055 721
rect 3237 277 3243 621
rect 4049 277 4055 621
rect 3237 261 4055 277
rect 4127 1063 4203 1151
rect 4127 721 4133 1063
rect 4197 721 4203 1063
rect 4127 621 4203 721
rect 4127 277 4133 621
rect 4197 277 4203 621
rect 4127 189 4203 277
rect 3089 177 4203 189
rect 3089 118 3095 177
rect 4197 118 4203 177
rect 3089 112 4203 118
rect 4275 1220 4287 1298
rect 4493 1298 5775 1304
rect 4493 1220 4505 1298
rect 4275 1163 4281 1220
rect 4499 1163 4505 1220
rect 4275 1063 4505 1163
rect 4275 721 4281 1063
rect 4499 721 4505 1063
rect 4275 621 4505 721
rect 4275 277 4281 621
rect 4499 277 4505 621
rect 4275 177 4505 277
rect 4275 118 4281 177
rect 4499 118 4505 177
rect 4275 40 4287 118
rect 3005 34 4287 40
rect 4493 40 4505 118
rect 4577 1220 5691 1226
rect 4577 1163 4583 1220
rect 5685 1163 5691 1220
rect 4577 1151 5691 1163
rect 4577 1063 4653 1151
rect 4577 721 4583 1063
rect 4647 721 4653 1063
rect 4577 621 4653 721
rect 4577 277 4583 621
rect 4647 277 4653 621
rect 4577 189 4653 277
rect 4725 1063 5543 1079
rect 4725 721 4731 1063
rect 5537 721 5543 1063
rect 4725 621 5543 721
rect 4725 277 4731 621
rect 5537 277 5543 621
rect 4725 261 5543 277
rect 5615 1063 5691 1151
rect 5615 721 5621 1063
rect 5685 721 5691 1063
rect 5615 621 5691 721
rect 5615 277 5621 621
rect 5685 277 5691 621
rect 5615 189 5691 277
rect 4577 177 5691 189
rect 4577 118 4583 177
rect 5685 118 5691 177
rect 4577 112 5691 118
rect 5763 1220 5775 1298
rect 5981 1298 7263 1304
rect 5981 1220 5993 1298
rect 5763 1163 5769 1220
rect 5987 1163 5993 1220
rect 5763 1063 5993 1163
rect 5763 721 5769 1063
rect 5987 721 5993 1063
rect 5763 621 5993 721
rect 5763 277 5769 621
rect 5987 277 5993 621
rect 5763 177 5993 277
rect 5763 118 5769 177
rect 5987 118 5993 177
rect 5763 40 5775 118
rect 4493 34 5775 40
rect 5981 40 5993 118
rect 6065 1220 7179 1226
rect 6065 1163 6071 1220
rect 6065 1157 6219 1163
rect 6572 1157 6672 1220
rect 7025 1157 7109 1163
rect 6065 1151 7115 1157
rect 6065 1063 6141 1151
rect 6065 721 6071 1063
rect 6135 721 6141 1063
rect 6065 621 6141 721
rect 6065 277 6071 621
rect 6135 277 6141 621
rect 6065 189 6141 277
rect 6213 1073 7031 1079
rect 6213 721 6219 1073
rect 6572 721 6672 1073
rect 6213 621 6672 721
rect 6213 267 6219 621
rect 7025 267 7031 1073
rect 6213 261 7031 267
rect 7103 1073 7115 1151
rect 7103 267 7109 1073
rect 7103 189 7115 267
rect 6065 183 7115 189
rect 6065 177 6219 183
rect 7025 177 7109 183
rect 6065 118 6071 177
rect 7173 118 7179 1220
rect 6065 112 7179 118
rect 7251 1220 7263 1298
rect 7251 118 7257 1220
rect 7251 40 7263 118
rect 5981 34 7263 40
rect 35 28 119 34
rect 1221 28 1305 34
rect 1523 28 1607 34
rect 2709 28 2793 34
rect 3011 28 3095 34
rect 4197 28 4281 34
rect 4499 28 4583 34
rect 5685 28 5769 34
rect 5987 28 6071 34
rect 7173 28 7257 34
<< via1 >>
rect 1853 4829 2463 5439
rect 3341 4829 3951 5439
rect 4829 4829 5439 5439
rect 1853 3341 2463 3951
rect 3341 3341 3951 3951
rect 4829 3735 5439 3951
rect 4829 3341 5439 3557
rect 1853 1853 2463 2463
rect 3341 1853 3951 2463
rect 4829 1853 5439 2463
<< metal2 >>
rect 1853 5439 2463 5449
rect 3341 5439 3951 5449
rect 2463 4829 3341 4919
rect 4829 5439 5439 5449
rect 3951 4829 4829 4919
rect 1853 4819 5439 4829
rect 2363 3961 2463 4819
rect 4829 3961 4929 4819
rect 1853 3951 2463 3961
rect 1853 3331 2463 3341
rect 3341 3951 3951 3961
rect 4829 3951 5439 3961
rect 4829 3725 5439 3735
rect 3951 3596 7749 3696
rect 3341 3331 3951 3341
rect 4829 3557 5439 3567
rect 4829 3331 5439 3341
rect 2363 2473 2463 3331
rect 4829 2473 4929 3331
rect 1853 2463 5439 2473
rect 2463 2373 3341 2463
rect 1853 1843 2463 1853
rect 3951 2373 4829 2463
rect 3341 1843 3951 1853
rect 4829 1843 5439 1853
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
array 0 4 1488 0 4 1488
timestamp 1760968059
transform 1 0 0 0 1 0
box 0 0 1340 1340
<< labels >>
flabel metal2 7703 3646 7703 3646 0 FreeSans 800 0 0 0 A
port 0 nsew
flabel metal2 4876 4394 4876 4394 0 FreeSans 800 0 0 0 B
port 1 nsew
flabel metal1 6613 4393 6613 4394 0 FreeSans 800 0 0 0 AVSS
port 2 nsew
<< end >>
