magic
tech sky130A
magscale 1 2
timestamp 1716133296
<< pwell >>
rect -4283 -310 4283 310
<< nmos >>
rect -4087 -100 -2087 100
rect -2029 -100 -29 100
rect 29 -100 2029 100
rect 2087 -100 4087 100
<< ndiff >>
rect -4145 88 -4087 100
rect -4145 -88 -4133 88
rect -4099 -88 -4087 88
rect -4145 -100 -4087 -88
rect -2087 88 -2029 100
rect -2087 -88 -2075 88
rect -2041 -88 -2029 88
rect -2087 -100 -2029 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 2029 88 2087 100
rect 2029 -88 2041 88
rect 2075 -88 2087 88
rect 2029 -100 2087 -88
rect 4087 88 4145 100
rect 4087 -88 4099 88
rect 4133 -88 4145 88
rect 4087 -100 4145 -88
<< ndiffc >>
rect -4133 -88 -4099 88
rect -2075 -88 -2041 88
rect -17 -88 17 88
rect 2041 -88 2075 88
rect 4099 -88 4133 88
<< psubdiff >>
rect -4247 240 -4151 274
rect 4151 240 4247 274
rect -4247 178 -4213 240
rect 4213 178 4247 240
rect -4247 -240 -4213 -178
rect 4213 -240 4247 -178
rect -4247 -274 -4151 -240
rect 4151 -274 4247 -240
<< psubdiffcont >>
rect -4151 240 4151 274
rect -4247 -178 -4213 178
rect 4213 -178 4247 178
rect -4151 -274 4151 -240
<< poly >>
rect -4087 172 -2087 188
rect -4087 138 -4071 172
rect -2103 138 -2087 172
rect -4087 100 -2087 138
rect -2029 172 -29 188
rect -2029 138 -2013 172
rect -45 138 -29 172
rect -2029 100 -29 138
rect 29 172 2029 188
rect 29 138 45 172
rect 2013 138 2029 172
rect 29 100 2029 138
rect 2087 172 4087 188
rect 2087 138 2103 172
rect 4071 138 4087 172
rect 2087 100 4087 138
rect -4087 -138 -2087 -100
rect -4087 -172 -4071 -138
rect -2103 -172 -2087 -138
rect -4087 -188 -2087 -172
rect -2029 -138 -29 -100
rect -2029 -172 -2013 -138
rect -45 -172 -29 -138
rect -2029 -188 -29 -172
rect 29 -138 2029 -100
rect 29 -172 45 -138
rect 2013 -172 2029 -138
rect 29 -188 2029 -172
rect 2087 -138 4087 -100
rect 2087 -172 2103 -138
rect 4071 -172 4087 -138
rect 2087 -188 4087 -172
<< polycont >>
rect -4071 138 -2103 172
rect -2013 138 -45 172
rect 45 138 2013 172
rect 2103 138 4071 172
rect -4071 -172 -2103 -138
rect -2013 -172 -45 -138
rect 45 -172 2013 -138
rect 2103 -172 4071 -138
<< locali >>
rect -4247 240 -4151 274
rect 4151 240 4247 274
rect -4247 178 -4213 240
rect 4213 178 4247 240
rect -4087 138 -4071 172
rect -2103 138 -2087 172
rect -2029 138 -2013 172
rect -45 138 -29 172
rect 29 138 45 172
rect 2013 138 2029 172
rect 2087 138 2103 172
rect 4071 138 4087 172
rect -4133 88 -4099 104
rect -4133 -104 -4099 -88
rect -2075 88 -2041 104
rect -2075 -104 -2041 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 2041 88 2075 104
rect 2041 -104 2075 -88
rect 4099 88 4133 104
rect 4099 -104 4133 -88
rect -4087 -172 -4071 -138
rect -2103 -172 -2087 -138
rect -2029 -172 -2013 -138
rect -45 -172 -29 -138
rect 29 -172 45 -138
rect 2013 -172 2029 -138
rect 2087 -172 2103 -138
rect 4071 -172 4087 -138
rect -4247 -240 -4213 -178
rect 4213 -240 4247 -178
rect -4247 -274 -4151 -240
rect 4151 -274 4247 -240
<< viali >>
rect -4071 138 -2103 172
rect -2013 138 -45 172
rect 45 138 2013 172
rect 2103 138 4071 172
rect -4133 -88 -4099 88
rect -2075 -88 -2041 88
rect -17 -88 17 88
rect 2041 -88 2075 88
rect 4099 -88 4133 88
rect -4071 -172 -2103 -138
rect -2013 -172 -45 -138
rect 45 -172 2013 -138
rect 2103 -172 4071 -138
<< metal1 >>
rect -4083 172 -2091 178
rect -4083 138 -4071 172
rect -2103 138 -2091 172
rect -4083 132 -2091 138
rect -2025 172 -33 178
rect -2025 138 -2013 172
rect -45 138 -33 172
rect -2025 132 -33 138
rect 33 172 2025 178
rect 33 138 45 172
rect 2013 138 2025 172
rect 33 132 2025 138
rect 2091 172 4083 178
rect 2091 138 2103 172
rect 4071 138 4083 172
rect 2091 132 4083 138
rect -4139 88 -4093 100
rect -4139 -88 -4133 88
rect -4099 -88 -4093 88
rect -4139 -100 -4093 -88
rect -2081 88 -2035 100
rect -2081 -88 -2075 88
rect -2041 -88 -2035 88
rect -2081 -100 -2035 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 2035 88 2081 100
rect 2035 -88 2041 88
rect 2075 -88 2081 88
rect 2035 -100 2081 -88
rect 4093 88 4139 100
rect 4093 -88 4099 88
rect 4133 -88 4139 88
rect 4093 -100 4139 -88
rect -4083 -138 -2091 -132
rect -4083 -172 -4071 -138
rect -2103 -172 -2091 -138
rect -4083 -178 -2091 -172
rect -2025 -138 -33 -132
rect -2025 -172 -2013 -138
rect -45 -172 -33 -138
rect -2025 -178 -33 -172
rect 33 -138 2025 -132
rect 33 -172 45 -138
rect 2013 -172 2025 -138
rect 33 -178 2025 -172
rect 2091 -138 4083 -132
rect 2091 -172 2103 -138
rect 4071 -172 4083 -138
rect 2091 -178 4083 -172
<< properties >>
string FIXED_BBOX -4230 -257 4230 257
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 10 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
