magic
tech sky130A
magscale 1 2
timestamp 1762707440
<< error_p >>
rect -4181 18 4181 236
<< nwell >>
rect -4181 18 4181 418
rect -4181 -418 4181 -18
<< pmos >>
rect -4087 118 -2087 318
rect -2029 118 -29 318
rect 29 118 2029 318
rect 2087 118 4087 318
rect -4087 -318 -2087 -118
rect -2029 -318 -29 -118
rect 29 -318 2029 -118
rect 2087 -318 4087 -118
<< pdiff >>
rect -4145 306 -4087 318
rect -4145 130 -4133 306
rect -4099 130 -4087 306
rect -4145 118 -4087 130
rect -2087 306 -2029 318
rect -2087 130 -2075 306
rect -2041 130 -2029 306
rect -2087 118 -2029 130
rect -29 306 29 318
rect -29 130 -17 306
rect 17 130 29 306
rect -29 118 29 130
rect 2029 306 2087 318
rect 2029 130 2041 306
rect 2075 130 2087 306
rect 2029 118 2087 130
rect 4087 306 4145 318
rect 4087 130 4099 306
rect 4133 130 4145 306
rect 4087 118 4145 130
rect -4145 -130 -4087 -118
rect -4145 -306 -4133 -130
rect -4099 -306 -4087 -130
rect -4145 -318 -4087 -306
rect -2087 -130 -2029 -118
rect -2087 -306 -2075 -130
rect -2041 -306 -2029 -130
rect -2087 -318 -2029 -306
rect -29 -130 29 -118
rect -29 -306 -17 -130
rect 17 -306 29 -130
rect -29 -318 29 -306
rect 2029 -130 2087 -118
rect 2029 -306 2041 -130
rect 2075 -306 2087 -130
rect 2029 -318 2087 -306
rect 4087 -130 4145 -118
rect 4087 -306 4099 -130
rect 4133 -306 4145 -130
rect 4087 -318 4145 -306
<< pdiffc >>
rect -4133 130 -4099 306
rect -2075 130 -2041 306
rect -17 130 17 306
rect 2041 130 2075 306
rect 4099 130 4133 306
rect -4133 -306 -4099 -130
rect -2075 -306 -2041 -130
rect -17 -306 17 -130
rect 2041 -306 2075 -130
rect 4099 -306 4133 -130
<< poly >>
rect -4087 399 -2087 415
rect -4087 365 -4071 399
rect -2103 365 -2087 399
rect -4087 318 -2087 365
rect -2029 399 -29 415
rect -2029 365 -2013 399
rect -45 365 -29 399
rect -2029 318 -29 365
rect 29 399 2029 415
rect 29 365 45 399
rect 2013 365 2029 399
rect 29 318 2029 365
rect 2087 399 4087 415
rect 2087 365 2103 399
rect 4071 365 4087 399
rect 2087 318 4087 365
rect -4087 71 -2087 118
rect -4087 37 -4071 71
rect -2103 37 -2087 71
rect -4087 21 -2087 37
rect -2029 71 -29 118
rect -2029 37 -2013 71
rect -45 37 -29 71
rect -2029 21 -29 37
rect 29 71 2029 118
rect 29 37 45 71
rect 2013 37 2029 71
rect 29 21 2029 37
rect 2087 71 4087 118
rect 2087 37 2103 71
rect 4071 37 4087 71
rect 2087 21 4087 37
rect -4087 -37 -2087 -21
rect -4087 -71 -4071 -37
rect -2103 -71 -2087 -37
rect -4087 -118 -2087 -71
rect -2029 -37 -29 -21
rect -2029 -71 -2013 -37
rect -45 -71 -29 -37
rect -2029 -118 -29 -71
rect 29 -37 2029 -21
rect 29 -71 45 -37
rect 2013 -71 2029 -37
rect 29 -118 2029 -71
rect 2087 -37 4087 -21
rect 2087 -71 2103 -37
rect 4071 -71 4087 -37
rect 2087 -118 4087 -71
rect -4087 -365 -2087 -318
rect -4087 -399 -4071 -365
rect -2103 -399 -2087 -365
rect -4087 -415 -2087 -399
rect -2029 -365 -29 -318
rect -2029 -399 -2013 -365
rect -45 -399 -29 -365
rect -2029 -415 -29 -399
rect 29 -365 2029 -318
rect 29 -399 45 -365
rect 2013 -399 2029 -365
rect 29 -415 2029 -399
rect 2087 -365 4087 -318
rect 2087 -399 2103 -365
rect 4071 -399 4087 -365
rect 2087 -415 4087 -399
<< polycont >>
rect -4071 365 -2103 399
rect -2013 365 -45 399
rect 45 365 2013 399
rect 2103 365 4071 399
rect -4071 37 -2103 71
rect -2013 37 -45 71
rect 45 37 2013 71
rect 2103 37 4071 71
rect -4071 -71 -2103 -37
rect -2013 -71 -45 -37
rect 45 -71 2013 -37
rect 2103 -71 4071 -37
rect -4071 -399 -2103 -365
rect -2013 -399 -45 -365
rect 45 -399 2013 -365
rect 2103 -399 4071 -365
<< locali >>
rect -4087 365 -4071 399
rect -2103 365 -2087 399
rect -2029 365 -2013 399
rect -45 365 -29 399
rect 29 365 45 399
rect 2013 365 2029 399
rect 2087 365 2103 399
rect 4071 365 4087 399
rect -4133 306 -4099 322
rect -4133 114 -4099 130
rect -2075 306 -2041 322
rect -2075 114 -2041 130
rect -17 306 17 322
rect -17 114 17 130
rect 2041 306 2075 322
rect 2041 114 2075 130
rect 4099 306 4133 322
rect 4099 114 4133 130
rect -4087 37 -4071 71
rect -2103 37 -2087 71
rect -2029 37 -2013 71
rect -45 37 -29 71
rect 29 37 45 71
rect 2013 37 2029 71
rect 2087 37 2103 71
rect 4071 37 4087 71
rect -4087 -71 -4071 -37
rect -2103 -71 -2087 -37
rect -2029 -71 -2013 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 2013 -71 2029 -37
rect 2087 -71 2103 -37
rect 4071 -71 4087 -37
rect -4133 -130 -4099 -114
rect -4133 -322 -4099 -306
rect -2075 -130 -2041 -114
rect -2075 -322 -2041 -306
rect -17 -130 17 -114
rect -17 -322 17 -306
rect 2041 -130 2075 -114
rect 2041 -322 2075 -306
rect 4099 -130 4133 -114
rect 4099 -322 4133 -306
rect -4087 -399 -4071 -365
rect -2103 -399 -2087 -365
rect -2029 -399 -2013 -365
rect -45 -399 -29 -365
rect 29 -399 45 -365
rect 2013 -399 2029 -365
rect 2087 -399 2103 -365
rect 4071 -399 4087 -365
<< viali >>
rect -4071 365 -2103 399
rect -2013 365 -45 399
rect 45 365 2013 399
rect 2103 365 4071 399
rect -4133 130 -4099 306
rect -2075 130 -2041 306
rect -17 130 17 306
rect 2041 130 2075 306
rect 4099 130 4133 306
rect -4071 37 -2103 71
rect -2013 37 -45 71
rect 45 37 2013 71
rect 2103 37 4071 71
rect -4071 -71 -2103 -37
rect -2013 -71 -45 -37
rect 45 -71 2013 -37
rect 2103 -71 4071 -37
rect -4133 -306 -4099 -130
rect -2075 -306 -2041 -130
rect -17 -306 17 -130
rect 2041 -306 2075 -130
rect 4099 -306 4133 -130
rect -4071 -399 -2103 -365
rect -2013 -399 -45 -365
rect 45 -399 2013 -365
rect 2103 -399 4071 -365
<< metal1 >>
rect -4083 399 -2091 405
rect -4083 365 -4071 399
rect -2103 365 -2091 399
rect -4083 359 -2091 365
rect -2025 399 -33 405
rect -2025 365 -2013 399
rect -45 365 -33 399
rect -2025 359 -33 365
rect 33 399 2025 405
rect 33 365 45 399
rect 2013 365 2025 399
rect 33 359 2025 365
rect 2091 399 4083 405
rect 2091 365 2103 399
rect 4071 365 4083 399
rect 2091 359 4083 365
rect -4139 306 -4093 318
rect -4139 130 -4133 306
rect -4099 130 -4093 306
rect -4139 118 -4093 130
rect -2081 306 -2035 318
rect -2081 130 -2075 306
rect -2041 130 -2035 306
rect -2081 118 -2035 130
rect -23 306 23 318
rect -23 130 -17 306
rect 17 130 23 306
rect -23 118 23 130
rect 2035 306 2081 318
rect 2035 130 2041 306
rect 2075 130 2081 306
rect 2035 118 2081 130
rect 4093 306 4139 318
rect 4093 130 4099 306
rect 4133 130 4139 306
rect 4093 118 4139 130
rect -4083 71 -2091 77
rect -4083 37 -4071 71
rect -2103 37 -2091 71
rect -4083 31 -2091 37
rect -2025 71 -33 77
rect -2025 37 -2013 71
rect -45 37 -33 71
rect -2025 31 -33 37
rect 33 71 2025 77
rect 33 37 45 71
rect 2013 37 2025 71
rect 33 31 2025 37
rect 2091 71 4083 77
rect 2091 37 2103 71
rect 4071 37 4083 71
rect 2091 31 4083 37
rect -4083 -37 -2091 -31
rect -4083 -71 -4071 -37
rect -2103 -71 -2091 -37
rect -4083 -77 -2091 -71
rect -2025 -37 -33 -31
rect -2025 -71 -2013 -37
rect -45 -71 -33 -37
rect -2025 -77 -33 -71
rect 33 -37 2025 -31
rect 33 -71 45 -37
rect 2013 -71 2025 -37
rect 33 -77 2025 -71
rect 2091 -37 4083 -31
rect 2091 -71 2103 -37
rect 4071 -71 4083 -37
rect 2091 -77 4083 -71
rect -4139 -130 -4093 -118
rect -4139 -306 -4133 -130
rect -4099 -306 -4093 -130
rect -4139 -318 -4093 -306
rect -2081 -130 -2035 -118
rect -2081 -306 -2075 -130
rect -2041 -306 -2035 -130
rect -2081 -318 -2035 -306
rect -23 -130 23 -118
rect -23 -306 -17 -130
rect 17 -306 23 -130
rect -23 -318 23 -306
rect 2035 -130 2081 -118
rect 2035 -306 2041 -130
rect 2075 -306 2081 -130
rect 2035 -318 2081 -306
rect 4093 -130 4139 -118
rect 4093 -306 4099 -130
rect 4133 -306 4139 -130
rect 4093 -318 4139 -306
rect -4083 -365 -2091 -359
rect -4083 -399 -4071 -365
rect -2103 -399 -2091 -365
rect -4083 -405 -2091 -399
rect -2025 -365 -33 -359
rect -2025 -399 -2013 -365
rect -45 -399 -33 -365
rect -2025 -405 -33 -399
rect 33 -365 2025 -359
rect 33 -399 45 -365
rect 2013 -399 2025 -365
rect 33 -405 2025 -399
rect 2091 -365 4083 -359
rect 2091 -399 2103 -365
rect 4071 -399 4083 -365
rect 2091 -405 4083 -399
<< labels >>
rlabel pdiffc -4116 -218 -4116 -218 0 D0_0
port 1 nsew
rlabel polycont -3087 -54 -3087 -54 0 G0_0
port 2 nsew
rlabel pdiffc -4116 218 -4116 218 0 D0_1
port 3 nsew
rlabel polycont -3087 382 -3087 382 0 G0_1
port 4 nsew
rlabel pdiffc -2058 -218 -2058 -218 0 S1_0
port 5 nsew
rlabel polycont -1029 -54 -1029 -54 0 G1_0
port 6 nsew
rlabel pdiffc -2058 218 -2058 218 0 S1_1
port 7 nsew
rlabel polycont -1029 382 -1029 382 0 G1_1
port 8 nsew
rlabel pdiffc 0 -218 0 -218 0 D2_0
port 9 nsew
rlabel polycont 1029 -54 1029 -54 0 G2_0
port 10 nsew
rlabel pdiffc 0 218 0 218 0 D2_1
port 11 nsew
rlabel polycont 1029 382 1029 382 0 G2_1
port 12 nsew
rlabel pdiffc 2058 -218 2058 -218 0 S3_0
port 13 nsew
rlabel polycont 3087 -54 3087 -54 0 G3_0
port 14 nsew
rlabel pdiffc 2058 218 2058 218 0 S3_1
port 15 nsew
rlabel polycont 3087 382 3087 382 0 G3_1
port 16 nsew
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 10 m 2 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 conn_gates 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 doports 1
<< end >>
