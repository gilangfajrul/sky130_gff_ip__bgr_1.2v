magic
tech sky130A
magscale 1 2
timestamp 1716453347
<< metal3 >>
rect -7904 7292 -4132 7320
rect -7904 3868 -4216 7292
rect -4152 3868 -4132 7292
rect -7904 3840 -4132 3868
rect -3892 7292 -120 7320
rect -3892 3868 -204 7292
rect -140 3868 -120 7292
rect -3892 3840 -120 3868
rect 120 7292 3892 7320
rect 120 3868 3808 7292
rect 3872 3868 3892 7292
rect 120 3840 3892 3868
rect 4132 7292 7904 7320
rect 4132 3868 7820 7292
rect 7884 3868 7904 7292
rect 4132 3840 7904 3868
rect -7904 3572 -4132 3600
rect -7904 148 -4216 3572
rect -4152 148 -4132 3572
rect -7904 120 -4132 148
rect -3892 3572 -120 3600
rect -3892 148 -204 3572
rect -140 148 -120 3572
rect -3892 120 -120 148
rect 120 3572 3892 3600
rect 120 148 3808 3572
rect 3872 148 3892 3572
rect 120 120 3892 148
rect 4132 3572 7904 3600
rect 4132 148 7820 3572
rect 7884 148 7904 3572
rect 4132 120 7904 148
rect -7904 -148 -4132 -120
rect -7904 -3572 -4216 -148
rect -4152 -3572 -4132 -148
rect -7904 -3600 -4132 -3572
rect -3892 -148 -120 -120
rect -3892 -3572 -204 -148
rect -140 -3572 -120 -148
rect -3892 -3600 -120 -3572
rect 120 -148 3892 -120
rect 120 -3572 3808 -148
rect 3872 -3572 3892 -148
rect 120 -3600 3892 -3572
rect 4132 -148 7904 -120
rect 4132 -3572 7820 -148
rect 7884 -3572 7904 -148
rect 4132 -3600 7904 -3572
rect -7904 -3868 -4132 -3840
rect -7904 -7292 -4216 -3868
rect -4152 -7292 -4132 -3868
rect -7904 -7320 -4132 -7292
rect -3892 -3868 -120 -3840
rect -3892 -7292 -204 -3868
rect -140 -7292 -120 -3868
rect -3892 -7320 -120 -7292
rect 120 -3868 3892 -3840
rect 120 -7292 3808 -3868
rect 3872 -7292 3892 -3868
rect 120 -7320 3892 -7292
rect 4132 -3868 7904 -3840
rect 4132 -7292 7820 -3868
rect 7884 -7292 7904 -3868
rect 4132 -7320 7904 -7292
<< via3 >>
rect -4216 3868 -4152 7292
rect -204 3868 -140 7292
rect 3808 3868 3872 7292
rect 7820 3868 7884 7292
rect -4216 148 -4152 3572
rect -204 148 -140 3572
rect 3808 148 3872 3572
rect 7820 148 7884 3572
rect -4216 -3572 -4152 -148
rect -204 -3572 -140 -148
rect 3808 -3572 3872 -148
rect 7820 -3572 7884 -148
rect -4216 -7292 -4152 -3868
rect -204 -7292 -140 -3868
rect 3808 -7292 3872 -3868
rect 7820 -7292 7884 -3868
<< mimcap >>
rect -7864 7240 -4464 7280
rect -7864 3920 -7824 7240
rect -4504 3920 -4464 7240
rect -7864 3880 -4464 3920
rect -3852 7240 -452 7280
rect -3852 3920 -3812 7240
rect -492 3920 -452 7240
rect -3852 3880 -452 3920
rect 160 7240 3560 7280
rect 160 3920 200 7240
rect 3520 3920 3560 7240
rect 160 3880 3560 3920
rect 4172 7240 7572 7280
rect 4172 3920 4212 7240
rect 7532 3920 7572 7240
rect 4172 3880 7572 3920
rect -7864 3520 -4464 3560
rect -7864 200 -7824 3520
rect -4504 200 -4464 3520
rect -7864 160 -4464 200
rect -3852 3520 -452 3560
rect -3852 200 -3812 3520
rect -492 200 -452 3520
rect -3852 160 -452 200
rect 160 3520 3560 3560
rect 160 200 200 3520
rect 3520 200 3560 3520
rect 160 160 3560 200
rect 4172 3520 7572 3560
rect 4172 200 4212 3520
rect 7532 200 7572 3520
rect 4172 160 7572 200
rect -7864 -200 -4464 -160
rect -7864 -3520 -7824 -200
rect -4504 -3520 -4464 -200
rect -7864 -3560 -4464 -3520
rect -3852 -200 -452 -160
rect -3852 -3520 -3812 -200
rect -492 -3520 -452 -200
rect -3852 -3560 -452 -3520
rect 160 -200 3560 -160
rect 160 -3520 200 -200
rect 3520 -3520 3560 -200
rect 160 -3560 3560 -3520
rect 4172 -200 7572 -160
rect 4172 -3520 4212 -200
rect 7532 -3520 7572 -200
rect 4172 -3560 7572 -3520
rect -7864 -3920 -4464 -3880
rect -7864 -7240 -7824 -3920
rect -4504 -7240 -4464 -3920
rect -7864 -7280 -4464 -7240
rect -3852 -3920 -452 -3880
rect -3852 -7240 -3812 -3920
rect -492 -7240 -452 -3920
rect -3852 -7280 -452 -7240
rect 160 -3920 3560 -3880
rect 160 -7240 200 -3920
rect 3520 -7240 3560 -3920
rect 160 -7280 3560 -7240
rect 4172 -3920 7572 -3880
rect 4172 -7240 4212 -3920
rect 7532 -7240 7572 -3920
rect 4172 -7280 7572 -7240
<< mimcapcontact >>
rect -7824 3920 -4504 7240
rect -3812 3920 -492 7240
rect 200 3920 3520 7240
rect 4212 3920 7532 7240
rect -7824 200 -4504 3520
rect -3812 200 -492 3520
rect 200 200 3520 3520
rect 4212 200 7532 3520
rect -7824 -3520 -4504 -200
rect -3812 -3520 -492 -200
rect 200 -3520 3520 -200
rect 4212 -3520 7532 -200
rect -7824 -7240 -4504 -3920
rect -3812 -7240 -492 -3920
rect 200 -7240 3520 -3920
rect 4212 -7240 7532 -3920
<< metal4 >>
rect -4232 7292 -4136 7308
rect -7825 7240 -4503 7241
rect -7825 3920 -7824 7240
rect -4504 3920 -4503 7240
rect -7825 3919 -4503 3920
rect -4232 3868 -4216 7292
rect -4152 3868 -4136 7292
rect -220 7292 -124 7308
rect -3813 7240 -491 7241
rect -3813 3920 -3812 7240
rect -492 3920 -491 7240
rect -3813 3919 -491 3920
rect -4232 3852 -4136 3868
rect -220 3868 -204 7292
rect -140 3868 -124 7292
rect 3792 7292 3888 7308
rect 199 7240 3521 7241
rect 199 3920 200 7240
rect 3520 3920 3521 7240
rect 199 3919 3521 3920
rect -220 3852 -124 3868
rect 3792 3868 3808 7292
rect 3872 3868 3888 7292
rect 7804 7292 7900 7308
rect 4211 7240 7533 7241
rect 4211 3920 4212 7240
rect 7532 3920 7533 7240
rect 4211 3919 7533 3920
rect 3792 3852 3888 3868
rect 7804 3868 7820 7292
rect 7884 3868 7900 7292
rect 7804 3852 7900 3868
rect -4232 3572 -4136 3588
rect -7825 3520 -4503 3521
rect -7825 200 -7824 3520
rect -4504 200 -4503 3520
rect -7825 199 -4503 200
rect -4232 148 -4216 3572
rect -4152 148 -4136 3572
rect -220 3572 -124 3588
rect -3813 3520 -491 3521
rect -3813 200 -3812 3520
rect -492 200 -491 3520
rect -3813 199 -491 200
rect -4232 132 -4136 148
rect -220 148 -204 3572
rect -140 148 -124 3572
rect 3792 3572 3888 3588
rect 199 3520 3521 3521
rect 199 200 200 3520
rect 3520 200 3521 3520
rect 199 199 3521 200
rect -220 132 -124 148
rect 3792 148 3808 3572
rect 3872 148 3888 3572
rect 7804 3572 7900 3588
rect 4211 3520 7533 3521
rect 4211 200 4212 3520
rect 7532 200 7533 3520
rect 4211 199 7533 200
rect 3792 132 3888 148
rect 7804 148 7820 3572
rect 7884 148 7900 3572
rect 7804 132 7900 148
rect -4232 -148 -4136 -132
rect -7825 -200 -4503 -199
rect -7825 -3520 -7824 -200
rect -4504 -3520 -4503 -200
rect -7825 -3521 -4503 -3520
rect -4232 -3572 -4216 -148
rect -4152 -3572 -4136 -148
rect -220 -148 -124 -132
rect -3813 -200 -491 -199
rect -3813 -3520 -3812 -200
rect -492 -3520 -491 -200
rect -3813 -3521 -491 -3520
rect -4232 -3588 -4136 -3572
rect -220 -3572 -204 -148
rect -140 -3572 -124 -148
rect 3792 -148 3888 -132
rect 199 -200 3521 -199
rect 199 -3520 200 -200
rect 3520 -3520 3521 -200
rect 199 -3521 3521 -3520
rect -220 -3588 -124 -3572
rect 3792 -3572 3808 -148
rect 3872 -3572 3888 -148
rect 7804 -148 7900 -132
rect 4211 -200 7533 -199
rect 4211 -3520 4212 -200
rect 7532 -3520 7533 -200
rect 4211 -3521 7533 -3520
rect 3792 -3588 3888 -3572
rect 7804 -3572 7820 -148
rect 7884 -3572 7900 -148
rect 7804 -3588 7900 -3572
rect -4232 -3868 -4136 -3852
rect -7825 -3920 -4503 -3919
rect -7825 -7240 -7824 -3920
rect -4504 -7240 -4503 -3920
rect -7825 -7241 -4503 -7240
rect -4232 -7292 -4216 -3868
rect -4152 -7292 -4136 -3868
rect -220 -3868 -124 -3852
rect -3813 -3920 -491 -3919
rect -3813 -7240 -3812 -3920
rect -492 -7240 -491 -3920
rect -3813 -7241 -491 -7240
rect -4232 -7308 -4136 -7292
rect -220 -7292 -204 -3868
rect -140 -7292 -124 -3868
rect 3792 -3868 3888 -3852
rect 199 -3920 3521 -3919
rect 199 -7240 200 -3920
rect 3520 -7240 3521 -3920
rect 199 -7241 3521 -7240
rect -220 -7308 -124 -7292
rect 3792 -7292 3808 -3868
rect 3872 -7292 3888 -3868
rect 7804 -3868 7900 -3852
rect 4211 -3920 7533 -3919
rect 4211 -7240 4212 -3920
rect 7532 -7240 7533 -3920
rect 4211 -7241 7533 -7240
rect 3792 -7308 3888 -7292
rect 7804 -7292 7820 -3868
rect 7884 -7292 7900 -3868
rect 7804 -7308 7900 -7292
<< properties >>
string FIXED_BBOX 4132 3840 7612 7320
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 17 l 17 val 590.92 carea 2.00 cperi 0.19 nx 4 ny 4 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 0 tconnect 0 ccov 100
<< end >>
