magic
tech sky130A
magscale 1 2
timestamp 1717000582
<< nwell >>
rect -2123 -309 2123 309
<< pmos >>
rect -2029 47 -29 247
rect 29 47 2029 247
rect -2029 -247 -29 -47
rect 29 -247 2029 -47
<< pdiff >>
rect -2087 235 -2029 247
rect -2087 59 -2075 235
rect -2041 59 -2029 235
rect -2087 47 -2029 59
rect -29 235 29 247
rect -29 59 -17 235
rect 17 59 29 235
rect -29 47 29 59
rect 2029 235 2087 247
rect 2029 59 2041 235
rect 2075 59 2087 235
rect 2029 47 2087 59
rect -2087 -59 -2029 -47
rect -2087 -235 -2075 -59
rect -2041 -235 -2029 -59
rect -2087 -247 -2029 -235
rect -29 -59 29 -47
rect -29 -235 -17 -59
rect 17 -235 29 -59
rect -29 -247 29 -235
rect 2029 -59 2087 -47
rect 2029 -235 2041 -59
rect 2075 -235 2087 -59
rect 2029 -247 2087 -235
<< pdiffc >>
rect -2075 59 -2041 235
rect -17 59 17 235
rect 2041 59 2075 235
rect -2075 -235 -2041 -59
rect -17 -235 17 -59
rect 2041 -235 2075 -59
<< poly >>
rect -2029 247 -29 273
rect 29 247 2029 273
rect -2029 21 -29 47
rect 29 21 2029 47
rect -2029 -47 -29 -21
rect 29 -47 2029 -21
rect -2029 -273 -29 -247
rect 29 -273 2029 -247
<< locali >>
rect -2075 235 -2041 251
rect -2075 43 -2041 59
rect -17 235 17 251
rect -17 43 17 59
rect 2041 235 2075 251
rect 2041 43 2075 59
rect -2075 -59 -2041 -43
rect -2075 -251 -2041 -235
rect -17 -59 17 -43
rect -17 -251 17 -235
rect 2041 -59 2075 -43
rect 2041 -251 2075 -235
<< viali >>
rect -2075 59 -2041 235
rect -17 59 17 235
rect 2041 59 2075 235
rect -2075 -235 -2041 -59
rect -17 -235 17 -59
rect 2041 -235 2075 -59
<< metal1 >>
rect -2081 235 -2035 247
rect -2081 59 -2075 235
rect -2041 59 -2035 235
rect -2081 47 -2035 59
rect -23 235 23 247
rect -23 59 -17 235
rect 17 59 23 235
rect -23 47 23 59
rect 2035 235 2081 247
rect 2035 59 2041 235
rect 2075 59 2081 235
rect 2035 47 2081 59
rect -2081 -59 -2035 -47
rect -2081 -235 -2075 -59
rect -2041 -235 -2035 -59
rect -2081 -247 -2035 -235
rect -23 -59 23 -47
rect -23 -235 -17 -59
rect 17 -235 23 -59
rect -23 -247 23 -235
rect 2035 -59 2081 -47
rect 2035 -235 2041 -59
rect 2075 -235 2081 -59
rect 2035 -247 2081 -235
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 10 m 2 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
