magic
tech sky130A
magscale 1 2
timestamp 1718095057
<< dnwell >>
rect 50494 9426 83924 10858
rect 50494 6051 78611 9426
rect 79871 9424 83924 9426
rect 79871 9423 81845 9424
rect 83323 9399 83924 9424
rect 50494 2852 78610 6051
rect 50494 1592 78608 2852
rect 79871 1721 82059 8163
rect 50494 459 78616 1592
rect 83324 464 83924 9399
rect 82420 461 83924 464
rect 82152 459 83924 461
rect 50494 -2911 83924 459
rect 50494 -2912 76268 -2911
rect 50494 -12406 68036 -2912
rect 69296 -11144 76268 -4172
rect 77528 -11144 83924 -2911
rect 77529 -12404 83924 -11144
rect 69296 -12406 83924 -12404
rect 50494 -13006 83924 -12406
<< nwell >>
rect 50414 10652 84004 10938
rect 50414 -12800 50700 10652
rect 67967 495 77368 4655
rect 83718 -12800 84004 10652
rect 50414 -13086 84004 -12800
<< pwell >>
rect 52104 4755 78348 9848
rect 79911 7574 80929 8123
rect 79911 6504 80504 7574
rect 52104 370 67949 4755
rect 79911 2894 82020 6504
rect 52104 -2759 77403 370
<< nsubdiff >>
rect 50451 10881 83967 10901
rect 50451 10847 50531 10881
rect 83887 10847 83967 10881
rect 50451 10827 83967 10847
rect 50451 10821 50525 10827
rect 50451 -12969 50471 10821
rect 50505 -12969 50525 10821
rect 50451 -12975 50525 -12969
rect 83893 10821 83967 10827
rect 83893 -12969 83913 10821
rect 83947 -12969 83967 10821
rect 83893 -12975 83967 -12969
rect 50451 -12995 83967 -12975
rect 50451 -13029 50531 -12995
rect 83887 -13029 83967 -12995
rect 50451 -13049 83967 -13029
<< nsubdiffcont >>
rect 50531 10847 83887 10881
rect 50471 -12969 50505 10821
rect 83913 -12969 83947 10821
rect 50531 -13029 83887 -12995
<< locali >>
rect 50471 10847 50531 10881
rect 83887 10847 83947 10881
rect 50471 10821 50505 10847
rect 50471 -12995 50505 -12969
rect 83913 10821 83947 10847
rect 83913 -12995 83947 -12969
rect 50471 -13029 50531 -12995
rect 83887 -13029 83947 -12995
<< metal1 >>
rect 79438 9189 79448 9212
rect 77959 9124 79448 9189
rect 79438 9068 79448 9124
rect 79598 9068 79608 9212
rect 77841 8510 78886 8627
rect 51879 7923 51951 7928
rect 51879 7922 52697 7923
rect 51951 7851 52697 7922
rect 51879 7844 51951 7850
rect 51720 7686 52697 7756
rect 51720 4052 51849 7686
rect 70157 7658 70167 7662
rect 69973 7657 70167 7658
rect 69537 7613 70167 7657
rect 69537 7566 70041 7613
rect 70157 7610 70167 7613
rect 70219 7610 70229 7662
rect 69537 7530 69587 7566
rect 73873 7331 73923 7520
rect 73873 7281 78592 7331
rect 78542 7083 78592 7281
rect 78541 7077 78593 7083
rect 78541 7019 78593 7025
rect 51978 6856 52702 6926
rect 51978 5252 52105 6856
rect 52198 6758 52264 6764
rect 52264 6692 52424 6758
rect 52198 6686 52264 6692
rect 51978 4933 51988 5252
rect 52095 4933 52105 5252
rect 78769 6097 78886 8510
rect 80603 7991 80949 8037
rect 80362 7771 80372 7947
rect 80424 7771 80434 7947
rect 80903 7594 80949 7991
rect 80012 7548 80949 7594
rect 80012 7231 80058 7548
rect 80092 7025 80102 7077
rect 80278 7025 80288 7077
rect 78769 5980 79719 6097
rect 79886 5980 79896 6096
rect 77507 5087 78354 5157
rect 78284 4322 78354 5087
rect 77635 4252 78354 4322
rect 51720 3994 68290 4052
rect 68244 3961 68290 3994
rect 68238 3295 68300 3961
rect 76468 3295 76530 3965
rect 73524 2365 73534 2417
rect 74518 2365 74528 2417
rect 75582 2364 75592 2416
rect 76576 2364 76586 2416
rect 67789 1952 68149 2011
rect 67789 -1473 67865 1952
rect 77635 1513 77705 4252
rect 77083 1455 77705 1513
rect 68234 1094 68280 1270
rect 72960 1143 72970 1319
rect 73022 1143 73032 1319
rect 77083 1131 77141 1455
rect 67894 1030 68280 1094
rect 67894 -45 67969 1030
rect 77079 462 77145 861
rect 68715 396 77145 462
rect 68715 136 68781 396
rect 68705 70 68715 136
rect 68781 70 68791 136
rect 72251 100 72261 192
rect 72493 160 72503 192
rect 72493 100 72595 160
rect 67894 -99 68202 -45
rect 68150 -175 68202 -99
rect 68703 -107 68713 -55
rect 69697 -107 69707 -55
rect 70761 -107 70771 -55
rect 71755 -107 71765 -55
rect 68141 -216 68193 -175
rect 72535 -219 72595 100
rect 77079 85 77145 396
rect 76662 19 77145 85
rect 76662 -118 76728 19
rect 72535 -279 72734 -219
rect 75755 -270 75960 -220
rect 75898 -908 75960 -270
rect 76251 -373 76261 -197
rect 76313 -373 76323 -197
rect 75898 -970 77027 -908
rect 68198 -1048 68204 -988
rect 68264 -1048 68270 -988
rect 68204 -1130 68264 -1048
rect 68204 -1208 68288 -1130
rect 68204 -1296 68264 -1208
rect 67783 -1479 67865 -1473
rect 67783 -1538 67789 -1479
rect 67783 -1545 67865 -1538
rect 76958 -2960 77027 -970
rect 76913 -3074 76923 -2960
rect 77062 -3074 77072 -2960
rect 78769 -3890 78886 5980
rect 80070 5753 80080 5805
rect 80856 5753 80866 5805
rect 81064 5753 81074 5805
rect 81850 5753 81860 5805
rect 80070 4861 80080 4913
rect 80856 4861 80866 4913
rect 81064 4861 81074 4913
rect 81850 4861 81860 4913
rect 80070 3969 80080 4021
rect 80856 3969 80866 4021
rect 81064 3969 81074 4021
rect 81850 3969 81860 4021
rect 80070 3077 80080 3129
rect 80856 3077 80866 3129
rect 81064 3077 81074 3129
rect 81850 3077 81860 3129
rect 74349 -4007 74355 -3890
rect 74472 -4007 78886 -3890
rect 73999 -6414 74009 -6114
rect 74309 -6414 74319 -6114
<< via1 >>
rect 79448 9068 79598 9212
rect 51879 7850 51951 7922
rect 70167 7610 70219 7662
rect 78541 7025 78593 7077
rect 52198 6692 52264 6758
rect 51988 4933 52095 5252
rect 80372 7771 80424 7947
rect 80102 7025 80278 7077
rect 79719 5980 79886 6096
rect 73534 2365 74518 2417
rect 75592 2364 76576 2416
rect 72970 1143 73022 1319
rect 68715 70 68781 136
rect 72261 100 72493 192
rect 68713 -107 69697 -55
rect 70771 -107 71755 -55
rect 76261 -373 76313 -197
rect 68204 -1048 68264 -988
rect 67789 -1538 67865 -1479
rect 76923 -3074 77062 -2960
rect 80080 5753 80856 5805
rect 81074 5753 81850 5805
rect 80080 4861 80856 4913
rect 81074 4861 81850 4913
rect 80080 3969 80856 4021
rect 81074 3969 81850 4021
rect 80080 3077 80856 3129
rect 81074 3077 81850 3129
rect 74355 -4007 74472 -3890
rect 74009 -6414 74309 -6114
<< metal2 >>
rect 79448 9212 79598 9222
rect 79448 9058 79598 9068
rect 79344 8524 79434 8533
rect 77958 8434 79344 8524
rect 79344 8425 79434 8434
rect 80372 7947 80424 7957
rect 51873 7850 51879 7922
rect 51951 7850 51957 7922
rect 70163 7666 70223 7676
rect 78300 7666 78356 7673
rect 80372 7666 80424 7771
rect 78298 7664 80424 7666
rect 78298 7608 78300 7664
rect 78356 7608 80424 7664
rect 78298 7606 80424 7608
rect 70163 7596 70223 7606
rect 78300 7599 78356 7606
rect 69436 7417 69492 7427
rect 69436 7351 69492 7361
rect 60950 7195 60960 7251
rect 61016 7195 61026 7251
rect 80102 7080 80278 7087
rect 78535 7077 80278 7080
rect 78535 7025 78541 7077
rect 78593 7025 80102 7077
rect 78535 7022 80278 7025
rect 80102 7015 80278 7022
rect 52203 6758 52259 6762
rect 52192 6692 52198 6758
rect 52264 6692 52270 6758
rect 52203 6688 52259 6692
rect 79719 6096 79886 6106
rect 80080 6065 80856 6075
rect 80080 5999 80856 6009
rect 79719 5970 79886 5980
rect 79760 5815 79820 5816
rect 79760 5807 81850 5815
rect 79820 5805 81850 5807
rect 79820 5753 80080 5805
rect 80856 5753 81074 5805
rect 79820 5751 81850 5753
rect 79760 5743 81850 5751
rect 79760 5742 79820 5743
rect 51973 5252 52110 5262
rect 51973 4933 51988 5252
rect 52095 4933 52110 5252
rect 80939 5127 80991 5743
rect 51973 3923 52110 4933
rect 79735 4932 79825 4941
rect 79825 4913 81850 4923
rect 79825 4861 80080 4913
rect 80856 4861 81074 4913
rect 79825 4851 81850 4861
rect 79735 4833 79825 4842
rect 60861 4428 67821 4437
rect 60861 4372 60870 4428
rect 60926 4372 67821 4428
rect 60861 4363 67821 4372
rect 51973 3786 67711 3923
rect 51980 3785 67711 3786
rect 67587 140 67711 3785
rect 67747 334 67821 4363
rect 80939 4229 80991 4851
rect 79798 4031 79864 4037
rect 79798 4028 81850 4031
rect 72355 3953 72411 3963
rect 79864 4021 81850 4028
rect 79864 3969 80080 4021
rect 80856 3969 81074 4021
rect 79864 3962 81850 3969
rect 79798 3959 81850 3962
rect 79798 3953 79864 3959
rect 72355 3767 72411 3777
rect 80939 3335 80991 3959
rect 67905 3118 68115 3196
rect 79790 3139 79856 3146
rect 79790 3136 81850 3139
rect 67905 519 67983 3118
rect 79856 3129 81850 3136
rect 79856 3077 80080 3129
rect 80856 3077 81074 3129
rect 79856 3070 81850 3077
rect 79790 3067 81850 3070
rect 79790 3060 79856 3067
rect 73534 2426 74518 2427
rect 75024 2426 75086 2778
rect 73534 2417 76576 2426
rect 74518 2416 76576 2417
rect 74518 2365 75592 2416
rect 73534 2355 74518 2365
rect 75592 2354 76576 2364
rect 72345 1331 72401 1341
rect 72345 1145 72401 1155
rect 72970 1319 73022 1329
rect 67905 441 72339 519
rect 72970 503 73022 1143
rect 72970 451 76313 503
rect 67747 260 70845 334
rect 68715 140 68781 146
rect 67587 136 68785 140
rect 67587 74 68715 136
rect 67587 -3136 67711 74
rect 68713 70 68715 74
rect 68781 70 68785 136
rect 68713 -45 68785 70
rect 68713 -55 69697 -45
rect 68713 -117 69697 -107
rect 70771 -49 70845 260
rect 72261 202 72339 441
rect 72261 192 72493 202
rect 72261 90 72493 100
rect 70771 -55 71755 -49
rect 70771 -117 71755 -107
rect 76261 -197 76313 451
rect 76261 -423 76313 -373
rect 67771 -750 68063 -749
rect 67762 -817 68063 -750
rect 67762 -1218 67848 -817
rect 68204 -988 68264 -982
rect 72679 -986 72740 -604
rect 68197 -1046 68204 -990
rect 68264 -1046 68271 -990
rect 68204 -1054 68264 -1048
rect 72428 -1047 72740 -986
rect 67762 -1318 67771 -1218
rect 67839 -1318 67848 -1218
rect 72428 -1341 72489 -1047
rect 67771 -1390 67839 -1380
rect 67783 -1479 67865 -1473
rect 67783 -1538 67789 -1479
rect 67865 -1538 68046 -1479
rect 67783 -1545 67865 -1538
rect 76545 -2008 76601 -1998
rect 76545 -2194 76601 -2184
rect 76923 -2960 77062 -2950
rect 76923 -3084 77062 -3074
rect 67587 -3260 72836 -3136
rect 72712 -3905 72836 -3260
rect 74355 -3890 74472 -3884
rect 74110 -4007 74355 -3890
rect 74110 -6104 74214 -4007
rect 74355 -4013 74472 -4007
rect 74009 -6114 74309 -6104
rect 74009 -6424 74309 -6414
<< via2 >>
rect 79448 9068 79598 9212
rect 79344 8434 79434 8524
rect 51884 7855 51946 7917
rect 70163 7662 70223 7666
rect 70163 7610 70167 7662
rect 70167 7610 70219 7662
rect 70219 7610 70223 7662
rect 70163 7606 70223 7610
rect 78300 7608 78356 7664
rect 69436 7361 69492 7417
rect 60960 7195 61016 7251
rect 52203 6697 52259 6753
rect 79719 5980 79886 6096
rect 80080 6009 80856 6065
rect 79760 5751 79820 5807
rect 79735 4842 79825 4932
rect 60870 4372 60926 4428
rect 79798 3962 79864 4028
rect 72355 3777 72411 3953
rect 79790 3070 79856 3136
rect 72345 1155 72401 1331
rect 72261 100 72493 192
rect 68206 -1046 68262 -990
rect 67771 -1380 67839 -1218
rect 76545 -2184 76601 -2008
rect 76923 -3074 77062 -2960
<< metal3 >>
rect 79438 9212 79608 9217
rect 79438 9068 79448 9212
rect 79598 9068 79608 9212
rect 79438 9063 79608 9068
rect 77942 8945 79278 9021
rect 78472 8434 78537 8435
rect 78462 8370 78472 8434
rect 78536 8370 78546 8434
rect 51879 7917 51951 7922
rect 51879 7866 51884 7917
rect 51865 7855 51884 7866
rect 51946 7866 51951 7917
rect 51946 7855 51966 7866
rect 51865 4307 51966 7855
rect 70153 7666 70233 7671
rect 78295 7666 78361 7669
rect 70153 7606 70163 7666
rect 70223 7664 78361 7666
rect 70223 7608 78300 7664
rect 78356 7608 78361 7664
rect 70223 7606 78361 7608
rect 70153 7601 70233 7606
rect 78295 7603 78361 7606
rect 69426 7417 69502 7422
rect 69426 7361 69436 7417
rect 69492 7361 69502 7417
rect 69426 7344 69502 7361
rect 78472 7344 78537 8370
rect 52198 7273 61021 7339
rect 52198 6753 52264 7273
rect 52198 6697 52203 6753
rect 52259 6697 52264 6753
rect 52198 6692 52264 6697
rect 60865 7251 61021 7273
rect 69426 7268 79123 7344
rect 60865 7195 60960 7251
rect 61016 7195 61021 7251
rect 60865 7185 61021 7195
rect 60865 6410 60931 7185
rect 60618 6344 60931 6410
rect 60618 4739 60684 6344
rect 60618 4673 60931 4739
rect 60865 4428 60931 4673
rect 60865 4372 60870 4428
rect 60926 4372 60931 4428
rect 60865 4367 60931 4372
rect 61380 4629 72433 4730
rect 61380 4307 61481 4629
rect 51865 4206 61481 4307
rect 72332 3953 72433 4629
rect 72332 3777 72355 3953
rect 72411 3777 72433 3953
rect 72332 3772 72433 3777
rect 76644 2638 76704 3224
rect 79047 3141 79123 7268
rect 79202 4033 79278 8945
rect 79339 8524 79439 8529
rect 79339 8434 79344 8524
rect 79434 8434 79439 8524
rect 79339 8429 79439 8434
rect 79346 4925 79422 8429
rect 79500 5818 79577 9063
rect 79709 6097 79896 6101
rect 79709 6096 80856 6097
rect 79709 5980 79719 6096
rect 79886 6070 80856 6096
rect 79886 6065 80866 6070
rect 79886 6009 80080 6065
rect 80856 6009 80866 6065
rect 79886 6004 80866 6009
rect 79886 5980 80856 6004
rect 79709 5975 79896 5980
rect 79500 5807 79825 5818
rect 79500 5751 79760 5807
rect 79820 5751 79825 5807
rect 79500 5741 79825 5751
rect 79730 4932 79830 4937
rect 79730 4925 79735 4932
rect 79346 4849 79735 4925
rect 79730 4842 79735 4849
rect 79825 4842 79830 4932
rect 79730 4837 79830 4842
rect 79202 4028 79869 4033
rect 79202 3962 79798 4028
rect 79864 3962 79869 4028
rect 79202 3957 79869 3962
rect 79047 3136 79866 3141
rect 79047 3070 79790 3136
rect 79856 3070 79866 3136
rect 79047 3065 79866 3070
rect 76644 2578 77447 2638
rect 72335 1331 72411 1336
rect 72335 1155 72345 1331
rect 72401 1155 72411 1331
rect 72335 1150 72411 1155
rect 72343 1090 72403 1150
rect 72343 1030 72564 1090
rect 68227 504 68287 798
rect 67815 444 68287 504
rect 67815 -988 67875 444
rect 72504 197 72564 1030
rect 72251 192 72564 197
rect 72251 100 72261 192
rect 72493 112 72564 192
rect 72493 100 72503 112
rect 72251 95 72503 100
rect 72262 -242 72322 95
rect 68201 -988 68267 -985
rect 67815 -990 68267 -988
rect 67815 -1046 68206 -990
rect 68262 -1046 68267 -990
rect 67815 -1048 68267 -1046
rect 68201 -1051 68267 -1048
rect 67761 -1218 67849 -1213
rect 67761 -1380 67771 -1218
rect 67839 -1380 67849 -1218
rect 67761 -1385 67849 -1380
rect 67762 -1854 67848 -1385
rect 67762 -1940 68263 -1854
rect 76535 -2008 76611 -2003
rect 76531 -2184 76541 -2008
rect 76605 -2184 76615 -2008
rect 76535 -2189 76611 -2184
rect 76538 -2262 76608 -2189
rect 77387 -2262 77447 2578
rect 76538 -2322 77447 -2262
rect 76913 -2960 77072 -2955
rect 76913 -3074 76923 -2960
rect 77062 -3074 77072 -2960
rect 76913 -3079 77072 -3074
<< via3 >>
rect 78472 8370 78536 8434
rect 76541 -2184 76545 -2008
rect 76545 -2184 76601 -2008
rect 76601 -2184 76605 -2008
rect 76923 -3074 77062 -2960
<< metal4 >>
rect 78471 8434 78537 8435
rect 77662 8370 78472 8434
rect 78536 8370 78537 8434
rect 77662 8369 78537 8370
rect 67793 -2816 67889 -1956
rect 76538 -2008 76608 -2007
rect 76538 -2184 76541 -2008
rect 76605 -2184 76608 -2008
rect 76538 -2816 76608 -2184
rect 67793 -2912 76608 -2816
rect 76922 -2960 77063 -2959
rect 76922 -2973 76923 -2960
rect 68214 -3054 76923 -2973
rect 68214 -3910 68293 -3054
rect 76922 -3074 76923 -3054
rect 77062 -3074 77063 -2960
rect 76922 -3075 77063 -3074
use bjt  bjt_0
timestamp 1717930986
transform 0 -1 76228 1 0 -11104
box 0 0 7324 6892
use cap_op  cap_op_0
timestamp 1718012278
transform 1 0 63910 0 1 -22
box -12037 -11160 4383 3480
use differential_pair  differential_pair_0
timestamp 1717432846
transform -1 0 71951 0 1 -764
box -567 -89 4001 858
use nmos_startup  nmos_startup_0
timestamp 1717696245
transform -1 0 76816 0 -1 -171
box -204 -148 746 686
use nmos_tail_current  nmos_tail_current_0
timestamp 1717870580
transform 1 0 68264 0 1 -2618
box -315 -141 8593 1579
use pmos_current_bgr  pmos_current_bgr_0
timestamp 1717985588
transform 1 0 68204 0 1 4099
box -227 -1493 8585 556
use pmos_current_bgr_2  pmos_current_bgr_2_0
timestamp 1717930986
transform 1 0 68192 0 1 1945
box -225 -1450 4471 516
use pmos_ena  pmos_ena_0
timestamp 1717771017
transform 1 0 80695 0 1 7108
box -191 -536 1237 466
use pmos_iptat  pmos_iptat_0
timestamp 1717930986
transform 1 0 72931 0 1 1632
box -191 -104 4438 898
use pmos_startup  pmos_startup_0
timestamp 1717930986
transform 1 0 72931 0 1 1031
box -191 -509 4437 439
use res_trim  res_trim_0
timestamp 1717917475
transform 0 -1 78047 1 0 8315
box -31 -51 1533 15873
use resist_const  resist_const_0
timestamp 1717597558
transform 1 0 49856 0 1 10331
box 2248 -3973 28492 -2077
use resistor_op_tt  resistor_op_tt_0
timestamp 1717870769
transform 0 1 70379 -1 0 -71
box -441 2216 791 5516
use resistorstart  resistorstart_0
timestamp 1717756107
transform -1 0 78052 0 -1 6266
box -53 -53 21855 1511
use trim  trim_0
timestamp 1717913952
transform 0 -1 80894 1 0 5750
box -182 -1121 756 979
use trim  trim_1
timestamp 1717913952
transform 0 -1 80894 1 0 4858
box -182 -1121 756 979
use trim  trim_2
timestamp 1717913952
transform 0 -1 80894 1 0 3966
box -182 -1121 756 979
use trim  trim_3
timestamp 1717913952
transform 0 -1 80894 1 0 3074
box -182 -1121 756 979
use vena  vena_0
timestamp 1717912414
transform 0 -1 80378 1 0 6764
box -182 -68 756 444
use vena  vena_1
timestamp 1717912414
transform 1 0 80111 0 1 7671
box -182 -68 756 444
<< labels >>
flabel pwell 76554 -1493 76554 -1493 0 FreeSans 800 0 0 0 D1
flabel pwell 76573 -1824 76573 -1824 0 FreeSans 800 0 0 0 D4
flabel pwell 76565 -1981 76565 -1981 0 FreeSans 800 0 0 0 D3
flabel pwell 72396 -1245 72396 -1245 0 FreeSans 800 0 0 0 S2
flabel pwell 68179 -375 68179 -375 0 FreeSans 800 0 0 0 D4
flabel pwell 70234 -783 70234 -783 0 FreeSans 800 0 0 0 S
flabel nwell 72377 3736 72377 3736 0 FreeSans 800 0 0 0 D1
flabel nwell 75009 3623 75009 3623 0 FreeSans 800 0 0 0 G
flabel nwell 76491 3691 76491 3691 0 FreeSans 800 0 0 0 D2
flabel nwell 72363 1364 72363 1364 0 FreeSans 800 0 0 0 D8
flabel nwell 72366 1591 72366 1591 0 FreeSans 800 0 0 0 D9
flabel nwell 72381 2019 72381 2019 0 FreeSans 800 0 0 0 D3
flabel nwell 72200 1973 72200 1973 0 FreeSans 800 0 0 0 D4
flabel pwell 70389 -363 70389 -363 0 FreeSans 800 0 0 0 Plus
flabel pwell 69881 -358 69881 -358 0 FreeSans 800 0 0 0 Minus
flabel metal1 52053 7716 52053 7716 0 FreeSans 800 0 0 0 C
flabel metal1 52271 6727 52271 6727 0 FreeSans 800 0 0 0 B
flabel metal3 60990 7191 60990 7191 0 FreeSans 800 270 0 0 E
flabel metal1 51996 6889 51996 6889 0 FreeSans 800 0 0 0 D
flabel via2 69478 7383 69478 7383 0 FreeSans 800 0 0 0 F
flabel pwell 68837 7468 68837 7469 0 FreeSans 800 0 0 0 VBGSC
flabel pwell 73932 7388 73932 7388 0 FreeSans 800 0 0 0 VBGTC
<< end >>
