magic
tech sky130A
magscale 1 2
timestamp 1717428712
<< metal1 >>
rect 3770 530 3860 560
rect -360 390 -330 480
rect 1440 430 1450 460
rect 1190 400 1450 430
rect -370 290 -360 390
rect -260 290 -250 390
rect 1440 370 1450 400
rect 1540 370 1550 460
rect 1440 220 1450 240
rect 1180 190 1450 220
rect 1440 150 1450 190
rect 1540 150 1550 240
rect 1700 140 1730 480
rect 1900 370 1910 460
rect 2000 430 2010 460
rect 2000 400 2250 430
rect 2000 370 2010 400
rect 1900 150 1910 240
rect 2000 220 2010 240
rect 3680 230 3690 330
rect 3790 230 3800 330
rect 2000 190 2250 220
rect 2000 150 2010 190
rect 3760 140 3790 230
rect -360 -100 -330 -10
rect 3830 -100 3860 530
rect -360 -130 3860 -100
<< via1 >>
rect -360 290 -260 390
rect 1450 370 1540 460
rect 1450 150 1540 240
rect 1910 370 2000 460
rect 1910 150 2000 240
rect 3690 230 3790 330
<< metal2 >>
rect -300 680 3730 720
rect -300 400 -260 680
rect -360 390 -260 400
rect 1450 460 1540 470
rect 1910 460 2000 470
rect 1540 390 1740 430
rect 1450 360 1540 370
rect -360 280 -260 290
rect 1450 240 1540 250
rect 1700 210 1740 390
rect 1910 360 2000 370
rect 3690 340 3730 680
rect 3690 330 3790 340
rect 1910 240 2000 250
rect 1700 170 1910 210
rect 1450 140 1540 150
rect 3690 220 3790 230
rect 1910 140 2000 150
<< via2 >>
rect 1450 150 1540 240
rect 1910 370 2000 460
<< metal3 >>
rect 1900 460 2010 465
rect 1900 450 1910 460
rect 1680 380 1910 450
rect 1440 240 1550 245
rect 1440 150 1450 240
rect 1540 230 1550 240
rect 1680 230 1750 380
rect 1900 370 1910 380
rect 2000 370 2010 460
rect 1900 365 2010 370
rect 1540 160 1750 230
rect 1540 150 1550 160
rect 1440 145 1550 150
use sky130_fd_pr__nfet_01v8_N7TR4F  sky130_fd_pr__nfet_01v8_N7TR4F_0
timestamp 1717428712
transform 1 0 1717 0 -1 517
box -2087 -137 2087 137
use sky130_fd_pr__nfet_01v8_N7TR4F  sky130_fd_pr__nfet_01v8_N7TR4F_1
timestamp 1717428712
transform 1 0 1717 0 1 97
box -2087 -137 2087 137
<< end >>
