magic
tech sky130A
magscale 1 2
timestamp 1716303658
<< nmos >>
rect -15 -80 15 80
<< ndiff >>
rect -73 68 -15 80
rect -73 -68 -61 68
rect -27 -68 -15 68
rect -73 -80 -15 -68
rect 15 68 73 80
rect 15 -68 27 68
rect 61 -68 73 68
rect 15 -80 73 -68
<< ndiffc >>
rect -61 -68 -27 68
rect 27 -68 61 68
<< poly >>
rect -15 80 15 106
rect -15 -106 15 -80
<< locali >>
rect -61 68 -27 84
rect -61 -84 -27 -68
rect 27 68 61 84
rect 27 -84 61 -68
<< viali >>
rect -61 -68 -27 68
rect 27 -68 61 68
<< metal1 >>
rect -67 68 -21 80
rect -67 -68 -61 68
rect -27 -68 -21 68
rect -67 -80 -21 -68
rect 21 68 67 80
rect 21 -68 27 68
rect 61 -68 67 68
rect 21 -80 67 -68
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.8 l 0.150 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
