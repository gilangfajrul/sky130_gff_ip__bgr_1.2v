magic
tech sky130A
magscale 1 2
timestamp 1718517160
<< pwell >>
rect -31 2797 1533 16353
rect -31 2792 618 2797
rect 706 2792 1533 2797
rect -31 -51 1533 2792
<< metal1 >>
rect 311 16214 1440 16264
rect 311 16169 361 16214
rect 643 16169 693 16214
rect 1390 16181 1440 16214
rect 134 16117 144 16169
rect 196 16117 206 16169
rect 466 16117 476 16169
rect 528 16117 538 16169
rect 798 16117 808 16169
rect 860 16117 870 16169
rect 1141 16131 1440 16181
rect 964 15944 974 15996
rect 1026 15944 1036 15996
rect 964 13785 974 13837
rect 1026 13785 1036 13837
rect 134 13613 144 13665
rect 196 13613 206 13665
rect 466 13613 476 13665
rect 528 13613 538 13665
rect 798 13613 808 13665
rect 860 13613 870 13665
rect 1390 13651 1440 16131
rect 311 13568 361 13613
rect 643 13568 693 13613
rect 1143 13601 1440 13651
rect 62 13518 1191 13568
rect 62 13485 112 13518
rect 62 13435 360 13485
rect 477 13473 527 13518
rect 809 13473 859 13518
rect 1141 13473 1191 13518
rect 1390 13485 1440 13601
rect 62 10955 112 13435
rect 632 13421 642 13473
rect 694 13421 704 13473
rect 964 13421 974 13473
rect 1026 13421 1036 13473
rect 1307 13435 1440 13485
rect 62 10905 361 10955
rect 632 10917 642 10969
rect 694 10917 704 10969
rect 964 10917 974 10969
rect 1026 10917 1036 10969
rect 1390 10955 1440 13435
rect 62 10789 112 10905
rect 477 10872 527 10917
rect 809 10872 859 10917
rect 1141 10872 1191 10917
rect 1307 10905 1440 10955
rect 1390 10872 1440 10905
rect 311 10822 1440 10872
rect 62 10739 195 10789
rect 311 10777 361 10822
rect 643 10777 693 10822
rect 975 10777 1025 10822
rect 1390 10789 1440 10822
rect 62 8259 112 10739
rect 466 10725 476 10777
rect 528 10725 538 10777
rect 798 10725 808 10777
rect 860 10725 870 10777
rect 1141 10739 1440 10789
rect 1390 10343 1440 10739
rect 1379 8655 1389 10343
rect 1441 8655 1451 10343
rect 62 8209 195 8259
rect 466 8221 476 8273
rect 528 8221 538 8273
rect 798 8221 808 8273
rect 860 8221 870 8273
rect 1390 8259 1440 8655
rect 62 8176 112 8209
rect 311 8176 361 8221
rect 643 8176 693 8221
rect 975 8176 1025 8221
rect 1141 8209 1440 8259
rect 62 8126 1191 8176
rect 62 8093 112 8126
rect 62 8043 361 8093
rect 477 8081 527 8126
rect 809 8081 859 8126
rect 1141 8081 1191 8126
rect 1390 8093 1440 8209
rect 62 5563 112 8043
rect 632 8029 642 8081
rect 694 8029 704 8081
rect 964 8029 974 8081
rect 1026 8029 1036 8081
rect 1307 8043 1440 8093
rect 1390 7647 1440 8043
rect 1379 5959 1389 7647
rect 1441 5959 1451 7647
rect 62 5513 360 5563
rect 632 5525 642 5577
rect 694 5525 704 5577
rect 964 5525 974 5577
rect 1026 5525 1036 5577
rect 1390 5563 1440 5959
rect 62 5397 112 5513
rect 477 5480 527 5525
rect 809 5480 859 5525
rect 1141 5480 1191 5525
rect 1307 5513 1440 5563
rect 1390 5480 1440 5513
rect 311 5430 1440 5480
rect 62 5347 195 5397
rect 311 5385 361 5430
rect 643 5385 693 5430
rect 975 5385 1025 5430
rect 1390 5397 1440 5430
rect 62 2867 112 5347
rect 466 5333 476 5385
rect 528 5333 538 5385
rect 798 5333 808 5385
rect 860 5333 870 5385
rect 1141 5347 1440 5397
rect 62 2817 188 2867
rect 466 2829 476 2881
rect 528 2829 538 2881
rect 798 2829 808 2881
rect 860 2829 870 2881
rect 1390 2867 1440 5347
rect 62 2784 112 2817
rect 311 2784 361 2829
rect 643 2784 693 2829
rect 975 2784 1025 2829
rect 1141 2817 1440 2867
rect 62 2734 1191 2784
rect 145 2691 195 2734
rect 228 171 278 2734
rect 311 2693 361 2734
rect 809 2689 859 2734
rect 1141 2689 1191 2734
rect 1390 2701 1440 2817
rect 632 2637 642 2689
rect 694 2637 704 2689
rect 964 2637 974 2689
rect 1026 2637 1036 2689
rect 1307 2651 1440 2701
rect 466 2464 476 2516
rect 528 2464 538 2516
rect 466 305 476 357
rect 528 305 538 357
rect 145 121 346 171
rect 632 133 642 185
rect 694 133 704 185
rect 964 133 974 185
rect 1026 133 1036 185
rect 1390 171 1440 2651
rect 809 88 859 133
rect 1141 88 1191 133
rect 1307 121 1440 171
rect 1390 88 1440 121
rect 809 38 1440 88
<< via1 >>
rect 144 16117 196 16169
rect 476 16117 528 16169
rect 808 16117 860 16169
rect 974 15944 1026 15996
rect 974 13785 1026 13837
rect 144 13613 196 13665
rect 476 13613 528 13665
rect 808 13613 860 13665
rect 642 13421 694 13473
rect 974 13421 1026 13473
rect 642 10917 694 10969
rect 974 10917 1026 10969
rect 476 10725 528 10777
rect 808 10725 860 10777
rect 1389 8655 1441 10343
rect 476 8221 528 8273
rect 808 8221 860 8273
rect 642 8029 694 8081
rect 974 8029 1026 8081
rect 1389 5959 1441 7647
rect 642 5525 694 5577
rect 974 5525 1026 5577
rect 476 5333 528 5385
rect 808 5333 860 5385
rect 476 2829 528 2881
rect 808 2829 860 2881
rect 642 2637 694 2689
rect 974 2637 1026 2689
rect 476 2464 528 2516
rect 476 305 528 357
rect 642 133 694 185
rect 974 133 1026 185
<< metal2 >>
rect 61 16209 528 16261
rect 61 16179 113 16209
rect 61 16169 196 16179
rect 61 16117 144 16169
rect 61 16107 196 16117
rect 476 16169 528 16209
rect 476 16107 528 16117
rect 806 16171 862 16181
rect 61 13675 113 16107
rect 806 16105 862 16115
rect 972 15998 1028 16008
rect 972 15932 1028 15942
rect 972 13839 1028 13849
rect 972 13773 1028 13783
rect 61 13665 196 13675
rect 61 13613 144 13665
rect 61 13603 196 13613
rect 476 13665 528 13675
rect 61 10873 113 13603
rect 476 13569 528 13613
rect 806 13667 862 13677
rect 806 13601 862 13611
rect 476 13517 1441 13569
rect 642 13473 694 13517
rect 642 13411 694 13421
rect 972 13475 1028 13485
rect 972 13409 1028 13419
rect 642 10969 694 10979
rect 642 10873 694 10917
rect 972 10971 1028 10981
rect 972 10905 1028 10915
rect 61 10821 860 10873
rect 61 10353 113 10821
rect 476 10777 528 10821
rect 476 10715 528 10725
rect 808 10777 860 10821
rect 808 10715 860 10725
rect 54 10343 120 10353
rect 54 8645 120 8655
rect 1389 10343 1441 13517
rect 61 7657 113 8645
rect 476 8273 528 8283
rect 476 8177 528 8221
rect 808 8273 860 8283
rect 808 8177 860 8221
rect 1389 8177 1441 8655
rect 476 8125 1441 8177
rect 642 8081 694 8125
rect 642 8019 694 8029
rect 974 8081 1026 8125
rect 974 8019 1026 8029
rect 54 7647 120 7657
rect 54 5949 120 5959
rect 1389 7647 1441 8125
rect 61 5481 113 5949
rect 642 5577 694 5587
rect 642 5481 694 5525
rect 974 5577 1026 5587
rect 974 5481 1026 5525
rect 61 5429 1026 5481
rect 61 89 113 5429
rect 474 5387 530 5397
rect 474 5321 530 5331
rect 808 5385 860 5429
rect 808 5323 860 5333
rect 474 2883 530 2893
rect 474 2817 530 2827
rect 808 2881 860 2891
rect 808 2785 860 2829
rect 1389 2785 1441 5959
rect 808 2733 1441 2785
rect 640 2691 696 2701
rect 640 2625 696 2635
rect 974 2689 1026 2733
rect 974 2627 1026 2637
rect 474 2518 530 2528
rect 474 2452 530 2462
rect 474 359 530 369
rect 474 293 530 303
rect 640 187 696 197
rect 640 121 696 131
rect 974 185 1026 195
rect 974 89 1026 133
rect 61 37 1026 89
<< via2 >>
rect 806 16169 862 16171
rect 806 16117 808 16169
rect 808 16117 860 16169
rect 860 16117 862 16169
rect 806 16115 862 16117
rect 972 15996 1028 15998
rect 972 15944 974 15996
rect 974 15944 1026 15996
rect 1026 15944 1028 15996
rect 972 15942 1028 15944
rect 972 13837 1028 13839
rect 972 13785 974 13837
rect 974 13785 1026 13837
rect 1026 13785 1028 13837
rect 972 13783 1028 13785
rect 806 13665 862 13667
rect 806 13613 808 13665
rect 808 13613 860 13665
rect 860 13613 862 13665
rect 806 13611 862 13613
rect 972 13473 1028 13475
rect 972 13421 974 13473
rect 974 13421 1026 13473
rect 1026 13421 1028 13473
rect 972 13419 1028 13421
rect 972 10969 1028 10971
rect 972 10917 974 10969
rect 974 10917 1026 10969
rect 1026 10917 1028 10969
rect 972 10915 1028 10917
rect 54 8655 120 10343
rect 54 5959 120 7647
rect 474 5385 530 5387
rect 474 5333 476 5385
rect 476 5333 528 5385
rect 528 5333 530 5385
rect 474 5331 530 5333
rect 474 2881 530 2883
rect 474 2829 476 2881
rect 476 2829 528 2881
rect 528 2829 530 2881
rect 474 2827 530 2829
rect 640 2689 696 2691
rect 640 2637 642 2689
rect 642 2637 694 2689
rect 694 2637 696 2689
rect 640 2635 696 2637
rect 474 2516 530 2518
rect 474 2464 476 2516
rect 476 2464 528 2516
rect 528 2464 530 2516
rect 474 2462 530 2464
rect 474 357 530 359
rect 474 305 476 357
rect 476 305 528 357
rect 528 305 530 357
rect 474 303 530 305
rect 640 185 696 187
rect 640 133 642 185
rect 642 133 694 185
rect 694 133 696 185
rect 640 131 696 133
<< metal3 >>
rect 796 16197 1448 16273
rect 796 16171 872 16197
rect 796 16115 806 16171
rect 862 16115 872 16171
rect 796 16110 872 16115
rect 962 16002 1038 16047
rect 958 15938 968 16002
rect 1032 15938 1042 16002
rect 962 15893 1038 15938
rect 962 13843 1038 13888
rect 958 13779 968 13843
rect 1032 13779 1042 13843
rect 962 13734 1038 13779
rect 796 13667 950 13672
rect 796 13611 806 13667
rect 862 13611 950 13667
rect 796 13576 950 13611
rect 54 13510 1038 13576
rect 54 10348 120 13510
rect 884 13475 1038 13510
rect 884 13419 972 13475
rect 1028 13419 1038 13475
rect 884 13414 1038 13419
rect 962 10971 1038 10976
rect 962 10915 972 10971
rect 1028 10915 1038 10971
rect 962 10885 1038 10915
rect 1382 10885 1448 16197
rect 962 10809 1448 10885
rect 44 10343 130 10348
rect 1382 10343 1448 10809
rect 44 8655 54 10343
rect 120 8655 130 10343
rect 1372 8655 1382 10343
rect 1448 8655 1458 10343
rect 44 8650 130 8655
rect 54 7652 120 8650
rect 44 7647 130 7652
rect 1382 7647 1448 8655
rect 44 5959 54 7647
rect 120 5959 130 7647
rect 1372 5959 1382 7647
rect 1448 5959 1458 7647
rect 44 5954 130 5959
rect 54 2792 120 5954
rect 1382 5493 1448 5959
rect 464 5417 1448 5493
rect 464 5387 540 5417
rect 464 5331 474 5387
rect 530 5331 540 5387
rect 464 5326 540 5331
rect 464 2883 618 2888
rect 464 2827 474 2883
rect 530 2827 618 2883
rect 464 2792 618 2827
rect 54 2726 706 2792
rect 552 2691 706 2726
rect 552 2635 640 2691
rect 696 2635 706 2691
rect 552 2630 706 2635
rect 464 2522 540 2567
rect 460 2458 470 2522
rect 534 2458 544 2522
rect 464 2413 540 2458
rect 464 363 540 407
rect 460 299 470 363
rect 534 299 544 363
rect 464 254 540 299
rect 630 187 706 192
rect 630 131 640 187
rect 696 131 706 187
rect 630 105 706 131
rect 1382 105 1448 5417
rect 630 29 1448 105
<< via3 >>
rect 968 15998 1032 16002
rect 968 15942 972 15998
rect 972 15942 1028 15998
rect 1028 15942 1032 15998
rect 968 15938 1032 15942
rect 968 13839 1032 13843
rect 968 13783 972 13839
rect 972 13783 1028 13839
rect 1028 13783 1032 13839
rect 968 13779 1032 13783
rect 1382 8655 1448 10343
rect 1382 5959 1448 7647
rect 470 2518 534 2522
rect 470 2462 474 2518
rect 474 2462 530 2518
rect 530 2462 534 2518
rect 470 2458 534 2462
rect 470 359 534 363
rect 470 303 474 359
rect 474 303 530 359
rect 530 303 534 359
rect 470 299 534 303
<< metal4 >>
rect 54 16002 1033 16003
rect 54 15938 968 16002
rect 1032 15938 1033 16002
rect 54 15937 1033 15938
rect 54 364 120 15937
rect 967 13843 1448 13844
rect 967 13779 968 13843
rect 1032 13779 1448 13843
rect 967 13778 1448 13779
rect 1382 10344 1448 13778
rect 1381 10343 1449 10344
rect 1381 8655 1382 10343
rect 1448 8655 1449 10343
rect 1381 8654 1449 8655
rect 1382 7648 1448 8654
rect 1381 7647 1449 7648
rect 1381 5959 1382 7647
rect 1448 5959 1449 7647
rect 1381 5958 1449 5959
rect 1382 2523 1448 5958
rect 469 2522 1448 2523
rect 469 2458 470 2522
rect 534 2458 1448 2522
rect 469 2457 1448 2458
rect 54 363 535 364
rect 54 299 470 363
rect 534 299 535 363
rect 54 298 535 299
use sky130_fd_pr__res_high_po_0p35_5N3J8V  sky130_fd_pr__res_high_po_0p35_5N3J8V_0
timestamp 1718386057
transform 1 0 751 0 1 8151
box -782 -8202 782 8202
<< labels >>
flabel pwell 12 -35 12 -35 0 FreeSans 1600 0 0 0 AVSS
port 4 nsew
flabel metal1 224 8148 224 8148 0 FreeSans 1600 0 0 0 B
port 0 nsew
flabel metal4 80 7714 80 7714 0 FreeSans 1600 0 0 0 A
port 1 nsew
flabel metal4 1420 8186 1420 8186 0 FreeSans 1600 0 0 0 1
port 5 nsew
flabel metal3 118 8310 118 8310 0 FreeSans 1600 0 0 0 2
port 6 nsew
flabel metal2 1418 8514 1418 8514 0 FreeSans 1600 0 0 0 3
port 7 nsew
<< end >>
