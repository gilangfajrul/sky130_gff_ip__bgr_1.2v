magic
tech sky130A
magscale 1 2
timestamp 1717755416
<< pwell >>
rect -782 -10954 782 10954
<< psubdiff >>
rect -746 10884 -650 10918
rect 650 10884 746 10918
rect -746 10822 -712 10884
rect 712 10822 746 10884
rect -746 -10884 -712 -10822
rect 712 -10884 746 -10822
rect -746 -10918 -650 -10884
rect 650 -10918 746 -10884
<< psubdiffcont >>
rect -650 10884 650 10918
rect -746 -10822 -712 10822
rect 712 -10822 746 10822
rect -650 -10918 650 -10884
<< xpolycontact >>
rect -616 10356 -546 10788
rect -616 6556 -546 6988
rect -450 10356 -380 10788
rect -450 6556 -380 6988
rect -284 10356 -214 10788
rect -284 6556 -214 6988
rect -118 10356 -48 10788
rect -118 6556 -48 6988
rect 48 10356 118 10788
rect 48 6556 118 6988
rect 214 10356 284 10788
rect 214 6556 284 6988
rect 380 10356 450 10788
rect 380 6556 450 6988
rect 546 10356 616 10788
rect 546 6556 616 6988
rect -616 6020 -546 6452
rect -616 2220 -546 2652
rect -450 6020 -380 6452
rect -450 2220 -380 2652
rect -284 6020 -214 6452
rect -284 2220 -214 2652
rect -118 6020 -48 6452
rect -118 2220 -48 2652
rect 48 6020 118 6452
rect 48 2220 118 2652
rect 214 6020 284 6452
rect 214 2220 284 2652
rect 380 6020 450 6452
rect 380 2220 450 2652
rect 546 6020 616 6452
rect 546 2220 616 2652
rect -616 1684 -546 2116
rect -616 -2116 -546 -1684
rect -450 1684 -380 2116
rect -450 -2116 -380 -1684
rect -284 1684 -214 2116
rect -284 -2116 -214 -1684
rect -118 1684 -48 2116
rect -118 -2116 -48 -1684
rect 48 1684 118 2116
rect 48 -2116 118 -1684
rect 214 1684 284 2116
rect 214 -2116 284 -1684
rect 380 1684 450 2116
rect 380 -2116 450 -1684
rect 546 1684 616 2116
rect 546 -2116 616 -1684
rect -616 -2652 -546 -2220
rect -616 -6452 -546 -6020
rect -450 -2652 -380 -2220
rect -450 -6452 -380 -6020
rect -284 -2652 -214 -2220
rect -284 -6452 -214 -6020
rect -118 -2652 -48 -2220
rect -118 -6452 -48 -6020
rect 48 -2652 118 -2220
rect 48 -6452 118 -6020
rect 214 -2652 284 -2220
rect 214 -6452 284 -6020
rect 380 -2652 450 -2220
rect 380 -6452 450 -6020
rect 546 -2652 616 -2220
rect 546 -6452 616 -6020
rect -616 -6988 -546 -6556
rect -616 -10788 -546 -10356
rect -450 -6988 -380 -6556
rect -450 -10788 -380 -10356
rect -284 -6988 -214 -6556
rect -284 -10788 -214 -10356
rect -118 -6988 -48 -6556
rect -118 -10788 -48 -10356
rect 48 -6988 118 -6556
rect 48 -10788 118 -10356
rect 214 -6988 284 -6556
rect 214 -10788 284 -10356
rect 380 -6988 450 -6556
rect 380 -10788 450 -10356
rect 546 -6988 616 -6556
rect 546 -10788 616 -10356
<< ppolyres >>
rect -616 6988 -546 10356
rect -450 6988 -380 10356
rect -284 6988 -214 10356
rect -118 6988 -48 10356
rect 48 6988 118 10356
rect 214 6988 284 10356
rect 380 6988 450 10356
rect 546 6988 616 10356
rect -616 2652 -546 6020
rect -450 2652 -380 6020
rect -284 2652 -214 6020
rect -118 2652 -48 6020
rect 48 2652 118 6020
rect 214 2652 284 6020
rect 380 2652 450 6020
rect 546 2652 616 6020
rect -616 -1684 -546 1684
rect -450 -1684 -380 1684
rect -284 -1684 -214 1684
rect -118 -1684 -48 1684
rect 48 -1684 118 1684
rect 214 -1684 284 1684
rect 380 -1684 450 1684
rect 546 -1684 616 1684
rect -616 -6020 -546 -2652
rect -450 -6020 -380 -2652
rect -284 -6020 -214 -2652
rect -118 -6020 -48 -2652
rect 48 -6020 118 -2652
rect 214 -6020 284 -2652
rect 380 -6020 450 -2652
rect 546 -6020 616 -2652
rect -616 -10356 -546 -6988
rect -450 -10356 -380 -6988
rect -284 -10356 -214 -6988
rect -118 -10356 -48 -6988
rect 48 -10356 118 -6988
rect 214 -10356 284 -6988
rect 380 -10356 450 -6988
rect 546 -10356 616 -6988
<< locali >>
rect -746 10884 -650 10918
rect 650 10884 746 10918
rect -746 10822 -712 10884
rect 712 10822 746 10884
rect -746 -10884 -712 -10822
rect 712 -10884 746 -10822
rect -746 -10918 -650 -10884
rect 650 -10918 746 -10884
<< viali >>
rect -600 10373 -562 10770
rect -434 10373 -396 10770
rect -268 10373 -230 10770
rect -102 10373 -64 10770
rect 64 10373 102 10770
rect 230 10373 268 10770
rect 396 10373 434 10770
rect 562 10373 600 10770
rect -600 6574 -562 6971
rect -434 6574 -396 6971
rect -268 6574 -230 6971
rect -102 6574 -64 6971
rect 64 6574 102 6971
rect 230 6574 268 6971
rect 396 6574 434 6971
rect 562 6574 600 6971
rect -600 6037 -562 6434
rect -434 6037 -396 6434
rect -268 6037 -230 6434
rect -102 6037 -64 6434
rect 64 6037 102 6434
rect 230 6037 268 6434
rect 396 6037 434 6434
rect 562 6037 600 6434
rect -600 2238 -562 2635
rect -434 2238 -396 2635
rect -268 2238 -230 2635
rect -102 2238 -64 2635
rect 64 2238 102 2635
rect 230 2238 268 2635
rect 396 2238 434 2635
rect 562 2238 600 2635
rect -600 1701 -562 2098
rect -434 1701 -396 2098
rect -268 1701 -230 2098
rect -102 1701 -64 2098
rect 64 1701 102 2098
rect 230 1701 268 2098
rect 396 1701 434 2098
rect 562 1701 600 2098
rect -600 -2098 -562 -1701
rect -434 -2098 -396 -1701
rect -268 -2098 -230 -1701
rect -102 -2098 -64 -1701
rect 64 -2098 102 -1701
rect 230 -2098 268 -1701
rect 396 -2098 434 -1701
rect 562 -2098 600 -1701
rect -600 -2635 -562 -2238
rect -434 -2635 -396 -2238
rect -268 -2635 -230 -2238
rect -102 -2635 -64 -2238
rect 64 -2635 102 -2238
rect 230 -2635 268 -2238
rect 396 -2635 434 -2238
rect 562 -2635 600 -2238
rect -600 -6434 -562 -6037
rect -434 -6434 -396 -6037
rect -268 -6434 -230 -6037
rect -102 -6434 -64 -6037
rect 64 -6434 102 -6037
rect 230 -6434 268 -6037
rect 396 -6434 434 -6037
rect 562 -6434 600 -6037
rect -600 -6971 -562 -6574
rect -434 -6971 -396 -6574
rect -268 -6971 -230 -6574
rect -102 -6971 -64 -6574
rect 64 -6971 102 -6574
rect 230 -6971 268 -6574
rect 396 -6971 434 -6574
rect 562 -6971 600 -6574
rect -600 -10770 -562 -10373
rect -434 -10770 -396 -10373
rect -268 -10770 -230 -10373
rect -102 -10770 -64 -10373
rect 64 -10770 102 -10373
rect 230 -10770 268 -10373
rect 396 -10770 434 -10373
rect 562 -10770 600 -10373
<< metal1 >>
rect -606 10770 -556 10782
rect -606 10373 -600 10770
rect -562 10373 -556 10770
rect -606 10361 -556 10373
rect -440 10770 -390 10782
rect -440 10373 -434 10770
rect -396 10373 -390 10770
rect -440 10361 -390 10373
rect -274 10770 -224 10782
rect -274 10373 -268 10770
rect -230 10373 -224 10770
rect -274 10361 -224 10373
rect -108 10770 -58 10782
rect -108 10373 -102 10770
rect -64 10373 -58 10770
rect -108 10361 -58 10373
rect 58 10770 108 10782
rect 58 10373 64 10770
rect 102 10373 108 10770
rect 58 10361 108 10373
rect 224 10770 274 10782
rect 224 10373 230 10770
rect 268 10373 274 10770
rect 224 10361 274 10373
rect 390 10770 440 10782
rect 390 10373 396 10770
rect 434 10373 440 10770
rect 390 10361 440 10373
rect 556 10770 606 10782
rect 556 10373 562 10770
rect 600 10373 606 10770
rect 556 10361 606 10373
rect -606 6971 -556 6983
rect -606 6574 -600 6971
rect -562 6574 -556 6971
rect -606 6562 -556 6574
rect -440 6971 -390 6983
rect -440 6574 -434 6971
rect -396 6574 -390 6971
rect -440 6562 -390 6574
rect -274 6971 -224 6983
rect -274 6574 -268 6971
rect -230 6574 -224 6971
rect -274 6562 -224 6574
rect -108 6971 -58 6983
rect -108 6574 -102 6971
rect -64 6574 -58 6971
rect -108 6562 -58 6574
rect 58 6971 108 6983
rect 58 6574 64 6971
rect 102 6574 108 6971
rect 58 6562 108 6574
rect 224 6971 274 6983
rect 224 6574 230 6971
rect 268 6574 274 6971
rect 224 6562 274 6574
rect 390 6971 440 6983
rect 390 6574 396 6971
rect 434 6574 440 6971
rect 390 6562 440 6574
rect 556 6971 606 6983
rect 556 6574 562 6971
rect 600 6574 606 6971
rect 556 6562 606 6574
rect -606 6434 -556 6446
rect -606 6037 -600 6434
rect -562 6037 -556 6434
rect -606 6025 -556 6037
rect -440 6434 -390 6446
rect -440 6037 -434 6434
rect -396 6037 -390 6434
rect -440 6025 -390 6037
rect -274 6434 -224 6446
rect -274 6037 -268 6434
rect -230 6037 -224 6434
rect -274 6025 -224 6037
rect -108 6434 -58 6446
rect -108 6037 -102 6434
rect -64 6037 -58 6434
rect -108 6025 -58 6037
rect 58 6434 108 6446
rect 58 6037 64 6434
rect 102 6037 108 6434
rect 58 6025 108 6037
rect 224 6434 274 6446
rect 224 6037 230 6434
rect 268 6037 274 6434
rect 224 6025 274 6037
rect 390 6434 440 6446
rect 390 6037 396 6434
rect 434 6037 440 6434
rect 390 6025 440 6037
rect 556 6434 606 6446
rect 556 6037 562 6434
rect 600 6037 606 6434
rect 556 6025 606 6037
rect -606 2635 -556 2647
rect -606 2238 -600 2635
rect -562 2238 -556 2635
rect -606 2226 -556 2238
rect -440 2635 -390 2647
rect -440 2238 -434 2635
rect -396 2238 -390 2635
rect -440 2226 -390 2238
rect -274 2635 -224 2647
rect -274 2238 -268 2635
rect -230 2238 -224 2635
rect -274 2226 -224 2238
rect -108 2635 -58 2647
rect -108 2238 -102 2635
rect -64 2238 -58 2635
rect -108 2226 -58 2238
rect 58 2635 108 2647
rect 58 2238 64 2635
rect 102 2238 108 2635
rect 58 2226 108 2238
rect 224 2635 274 2647
rect 224 2238 230 2635
rect 268 2238 274 2635
rect 224 2226 274 2238
rect 390 2635 440 2647
rect 390 2238 396 2635
rect 434 2238 440 2635
rect 390 2226 440 2238
rect 556 2635 606 2647
rect 556 2238 562 2635
rect 600 2238 606 2635
rect 556 2226 606 2238
rect -606 2098 -556 2110
rect -606 1701 -600 2098
rect -562 1701 -556 2098
rect -606 1689 -556 1701
rect -440 2098 -390 2110
rect -440 1701 -434 2098
rect -396 1701 -390 2098
rect -440 1689 -390 1701
rect -274 2098 -224 2110
rect -274 1701 -268 2098
rect -230 1701 -224 2098
rect -274 1689 -224 1701
rect -108 2098 -58 2110
rect -108 1701 -102 2098
rect -64 1701 -58 2098
rect -108 1689 -58 1701
rect 58 2098 108 2110
rect 58 1701 64 2098
rect 102 1701 108 2098
rect 58 1689 108 1701
rect 224 2098 274 2110
rect 224 1701 230 2098
rect 268 1701 274 2098
rect 224 1689 274 1701
rect 390 2098 440 2110
rect 390 1701 396 2098
rect 434 1701 440 2098
rect 390 1689 440 1701
rect 556 2098 606 2110
rect 556 1701 562 2098
rect 600 1701 606 2098
rect 556 1689 606 1701
rect -606 -1701 -556 -1689
rect -606 -2098 -600 -1701
rect -562 -2098 -556 -1701
rect -606 -2110 -556 -2098
rect -440 -1701 -390 -1689
rect -440 -2098 -434 -1701
rect -396 -2098 -390 -1701
rect -440 -2110 -390 -2098
rect -274 -1701 -224 -1689
rect -274 -2098 -268 -1701
rect -230 -2098 -224 -1701
rect -274 -2110 -224 -2098
rect -108 -1701 -58 -1689
rect -108 -2098 -102 -1701
rect -64 -2098 -58 -1701
rect -108 -2110 -58 -2098
rect 58 -1701 108 -1689
rect 58 -2098 64 -1701
rect 102 -2098 108 -1701
rect 58 -2110 108 -2098
rect 224 -1701 274 -1689
rect 224 -2098 230 -1701
rect 268 -2098 274 -1701
rect 224 -2110 274 -2098
rect 390 -1701 440 -1689
rect 390 -2098 396 -1701
rect 434 -2098 440 -1701
rect 390 -2110 440 -2098
rect 556 -1701 606 -1689
rect 556 -2098 562 -1701
rect 600 -2098 606 -1701
rect 556 -2110 606 -2098
rect -606 -2238 -556 -2226
rect -606 -2635 -600 -2238
rect -562 -2635 -556 -2238
rect -606 -2647 -556 -2635
rect -440 -2238 -390 -2226
rect -440 -2635 -434 -2238
rect -396 -2635 -390 -2238
rect -440 -2647 -390 -2635
rect -274 -2238 -224 -2226
rect -274 -2635 -268 -2238
rect -230 -2635 -224 -2238
rect -274 -2647 -224 -2635
rect -108 -2238 -58 -2226
rect -108 -2635 -102 -2238
rect -64 -2635 -58 -2238
rect -108 -2647 -58 -2635
rect 58 -2238 108 -2226
rect 58 -2635 64 -2238
rect 102 -2635 108 -2238
rect 58 -2647 108 -2635
rect 224 -2238 274 -2226
rect 224 -2635 230 -2238
rect 268 -2635 274 -2238
rect 224 -2647 274 -2635
rect 390 -2238 440 -2226
rect 390 -2635 396 -2238
rect 434 -2635 440 -2238
rect 390 -2647 440 -2635
rect 556 -2238 606 -2226
rect 556 -2635 562 -2238
rect 600 -2635 606 -2238
rect 556 -2647 606 -2635
rect -606 -6037 -556 -6025
rect -606 -6434 -600 -6037
rect -562 -6434 -556 -6037
rect -606 -6446 -556 -6434
rect -440 -6037 -390 -6025
rect -440 -6434 -434 -6037
rect -396 -6434 -390 -6037
rect -440 -6446 -390 -6434
rect -274 -6037 -224 -6025
rect -274 -6434 -268 -6037
rect -230 -6434 -224 -6037
rect -274 -6446 -224 -6434
rect -108 -6037 -58 -6025
rect -108 -6434 -102 -6037
rect -64 -6434 -58 -6037
rect -108 -6446 -58 -6434
rect 58 -6037 108 -6025
rect 58 -6434 64 -6037
rect 102 -6434 108 -6037
rect 58 -6446 108 -6434
rect 224 -6037 274 -6025
rect 224 -6434 230 -6037
rect 268 -6434 274 -6037
rect 224 -6446 274 -6434
rect 390 -6037 440 -6025
rect 390 -6434 396 -6037
rect 434 -6434 440 -6037
rect 390 -6446 440 -6434
rect 556 -6037 606 -6025
rect 556 -6434 562 -6037
rect 600 -6434 606 -6037
rect 556 -6446 606 -6434
rect -606 -6574 -556 -6562
rect -606 -6971 -600 -6574
rect -562 -6971 -556 -6574
rect -606 -6983 -556 -6971
rect -440 -6574 -390 -6562
rect -440 -6971 -434 -6574
rect -396 -6971 -390 -6574
rect -440 -6983 -390 -6971
rect -274 -6574 -224 -6562
rect -274 -6971 -268 -6574
rect -230 -6971 -224 -6574
rect -274 -6983 -224 -6971
rect -108 -6574 -58 -6562
rect -108 -6971 -102 -6574
rect -64 -6971 -58 -6574
rect -108 -6983 -58 -6971
rect 58 -6574 108 -6562
rect 58 -6971 64 -6574
rect 102 -6971 108 -6574
rect 58 -6983 108 -6971
rect 224 -6574 274 -6562
rect 224 -6971 230 -6574
rect 268 -6971 274 -6574
rect 224 -6983 274 -6971
rect 390 -6574 440 -6562
rect 390 -6971 396 -6574
rect 434 -6971 440 -6574
rect 390 -6983 440 -6971
rect 556 -6574 606 -6562
rect 556 -6971 562 -6574
rect 600 -6971 606 -6574
rect 556 -6983 606 -6971
rect -606 -10373 -556 -10361
rect -606 -10770 -600 -10373
rect -562 -10770 -556 -10373
rect -606 -10782 -556 -10770
rect -440 -10373 -390 -10361
rect -440 -10770 -434 -10373
rect -396 -10770 -390 -10373
rect -440 -10782 -390 -10770
rect -274 -10373 -224 -10361
rect -274 -10770 -268 -10373
rect -230 -10770 -224 -10373
rect -274 -10782 -224 -10770
rect -108 -10373 -58 -10361
rect -108 -10770 -102 -10373
rect -64 -10770 -58 -10373
rect -108 -10782 -58 -10770
rect 58 -10373 108 -10361
rect 58 -10770 64 -10373
rect 102 -10770 108 -10373
rect 58 -10782 108 -10770
rect 224 -10373 274 -10361
rect 224 -10770 230 -10373
rect 268 -10770 274 -10373
rect 224 -10782 274 -10770
rect 390 -10373 440 -10361
rect 390 -10770 396 -10373
rect 434 -10770 440 -10373
rect 390 -10782 440 -10770
rect 556 -10373 606 -10361
rect 556 -10770 562 -10373
rect 600 -10770 606 -10373
rect 556 -10782 606 -10770
<< properties >>
string FIXED_BBOX -729 -10901 729 10901
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.350 l 17 m 5 nx 8 wmin 0.350 lmin 0.50 rho 319.8 val 16.646k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
