magic
tech sky130A
magscale 1 2
timestamp 1716632848
<< metal1 >>
rect 350 13175 400 13220
rect 682 13175 732 13220
rect 350 13125 732 13175
rect 516 10559 566 10604
rect 599 10559 649 13125
rect 848 10559 898 10633
rect 1180 10559 1230 10604
rect 516 10509 1230 10559
rect 350 7943 400 7988
rect 682 7943 732 7980
rect 765 7943 815 10509
rect 1014 7943 1064 7976
rect 350 7893 1230 7943
rect 516 7848 566 7893
rect 599 5327 649 7893
rect 848 7848 898 7893
rect 1180 7848 1230 7893
rect 350 5277 1064 5327
rect 350 5232 400 5277
rect 682 5232 732 5277
rect 931 2711 981 5277
rect 1014 5232 1064 5277
rect 848 2661 1230 2711
rect 848 2616 898 2661
rect 1180 2616 1230 2661
use sky130_fd_pr__res_high_po_0p35_KQ9YB9  sky130_fd_pr__res_high_po_0p35_KQ9YB9_0
timestamp 1716599135
transform -1 0 790 0 -1 7918
box -843 -7971 843 7971
<< end >>
