magic
tech sky130A
magscale 1 2
timestamp 1717768872
<< nwell >>
rect -323 -264 323 298
<< pmos >>
rect -229 -164 -29 236
rect 29 -164 229 236
<< pdiff >>
rect -287 224 -229 236
rect -287 -152 -275 224
rect -241 -152 -229 224
rect -287 -164 -229 -152
rect -29 224 29 236
rect -29 -152 -17 224
rect 17 -152 29 224
rect -29 -164 29 -152
rect 229 224 287 236
rect 229 -152 241 224
rect 275 -152 287 224
rect 229 -164 287 -152
<< pdiffc >>
rect -275 -152 -241 224
rect -17 -152 17 224
rect 241 -152 275 224
<< poly >>
rect -229 236 -29 262
rect 29 236 229 262
rect -229 -211 -29 -164
rect -229 -228 -171 -211
rect -187 -245 -171 -228
rect -87 -228 -29 -211
rect 29 -211 229 -164
rect 29 -228 87 -211
rect -87 -245 -71 -228
rect -187 -261 -71 -245
rect 71 -245 87 -228
rect 171 -228 229 -211
rect 171 -245 187 -228
rect 71 -261 187 -245
<< polycont >>
rect -171 -245 -87 -211
rect 87 -245 171 -211
<< locali >>
rect -275 224 -241 240
rect -275 -168 -241 -152
rect -17 224 17 240
rect -17 -168 17 -152
rect 241 224 275 240
rect 241 -168 275 -152
rect -187 -245 -171 -211
rect -87 -245 -71 -211
rect 71 -245 87 -211
rect 171 -245 187 -211
<< viali >>
rect -275 -152 -241 224
rect -17 -152 17 224
rect 241 -152 275 224
rect -171 -245 -87 -211
rect 87 -245 171 -211
<< metal1 >>
rect -281 224 -235 236
rect -281 -152 -275 224
rect -241 -152 -235 224
rect -281 -164 -235 -152
rect -23 224 23 236
rect -23 -152 -17 224
rect 17 -152 23 224
rect -23 -164 23 -152
rect 235 224 281 236
rect 235 -152 241 224
rect 275 -152 281 224
rect 235 -164 281 -152
rect -183 -211 -75 -205
rect -183 -245 -171 -211
rect -87 -245 -75 -211
rect -183 -251 -75 -245
rect 75 -211 183 -205
rect 75 -245 87 -211
rect 171 -245 183 -211
rect 75 -251 183 -245
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2 l 1 m 1 nf 2 diffcov 100 polycov 50 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
