magic
tech sky130A
magscale 1 2
timestamp 1716190229
<< nwell >>
rect 680 15 5394 648
<< nsubdiff >>
rect 716 523 776 557
rect 5298 523 5358 557
rect 716 497 750 523
rect 5324 497 5358 523
rect 716 85 750 111
rect 5324 85 5358 111
rect 716 51 776 85
rect 5298 51 5358 85
<< nsubdiffcont >>
rect 776 523 5298 557
rect 716 111 750 497
rect 5324 111 5358 497
rect 776 51 5298 85
<< poly >>
rect 798 422 892 470
rect 862 411 892 422
rect 1137 417 1763 458
rect 2195 417 2821 458
rect 3253 417 3879 458
rect 4311 417 4937 458
rect 5182 422 5276 470
rect 2191 408 2829 417
rect 3249 408 3887 417
rect 4307 408 4945 417
rect 5182 391 5212 422
<< locali >>
rect 716 523 776 557
rect 5298 523 5358 557
rect 716 497 750 523
rect 5324 497 5358 523
rect 5224 391 5258 395
rect 716 85 750 111
rect 5324 85 5358 111
rect 716 51 776 85
rect 5298 51 5358 85
<< viali >>
rect 716 383 750 457
rect 811 429 879 463
rect 1150 417 1750 451
rect 2208 417 2808 451
rect 3266 417 3866 451
rect 4324 417 4924 451
rect 5195 429 5263 463
rect 5324 383 5358 457
rect 2981 51 3093 85
<< metal1 >>
rect 1138 470 4936 510
rect 710 463 891 469
rect 710 457 811 463
rect 710 383 716 457
rect 750 429 811 457
rect 879 429 891 463
rect 750 423 891 429
rect 1138 451 1762 470
rect 750 383 756 423
rect 810 391 856 423
rect 1138 417 1150 451
rect 1750 417 1762 451
rect 1138 411 1762 417
rect 2196 451 2820 470
rect 2196 417 2208 451
rect 2808 417 2820 451
rect 2196 411 2820 417
rect 3254 451 3878 470
rect 3254 417 3266 451
rect 3866 417 3878 451
rect 3254 411 3878 417
rect 4312 451 4936 470
rect 4312 417 4324 451
rect 4924 417 4936 451
rect 5183 463 5364 469
rect 5183 429 5195 463
rect 5263 457 5364 463
rect 5263 429 5324 457
rect 5183 423 5324 429
rect 4312 411 4936 417
rect 5218 391 5264 423
rect 710 371 756 383
rect 5318 383 5324 423
rect 5358 383 5364 457
rect 885 237 895 379
rect 947 237 957 379
rect 885 203 957 237
rect 3001 203 3011 379
rect 3063 203 3073 379
rect 5117 237 5127 379
rect 5179 237 5189 379
rect 5318 371 5364 383
rect 5117 203 5189 237
rect 1956 157 2002 195
rect 4072 157 4118 191
rect 1955 125 4118 157
rect 3011 91 3063 125
rect 2969 85 3105 91
rect 2969 51 2981 85
rect 3093 51 3105 85
rect 2969 45 3105 51
<< via1 >>
rect 895 237 947 379
rect 3011 203 3063 379
rect 5127 237 5179 379
<< metal2 >>
rect 895 379 947 389
rect 895 159 947 237
rect 3011 379 3063 389
rect 3011 159 3063 203
rect 5127 379 5179 389
rect 5127 159 5179 237
rect 895 111 5179 159
use sky130_fd_pr__pfet_01v8_2XU96L  sky130_fd_pr__pfet_01v8_2XU96L_0
timestamp 1716189928
transform 1 0 5197 0 1 291
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XU96L  sky130_fd_pr__pfet_01v8_2XU96L_1
timestamp 1716189928
transform 1 0 877 0 1 291
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_9QGYG3  sky130_fd_pr__pfet_01v8_9QGYG3_0
timestamp 1716188352
transform 1 0 3037 0 1 291
box -2181 -162 2181 162
<< end >>
