magic
tech sky130A
magscale 1 2
timestamp 1720112176
<< nwell >>
rect -250 -1450 4496 516
<< nsubdiff >>
rect -214 446 -129 480
rect 4375 446 4460 480
rect -214 420 -180 446
rect 4426 420 4460 446
rect -214 -1380 -180 -1354
rect 4426 -1380 4460 -1354
rect -214 -1414 -129 -1380
rect 4375 -1414 4460 -1380
<< nsubdiffcont >>
rect -129 446 4375 480
rect -214 -1354 -180 420
rect 4426 -1354 4460 420
rect -129 -1414 4375 -1380
<< poly >>
rect -56 381 36 397
rect -56 347 -40 381
rect -6 347 36 381
rect -56 331 36 347
rect 6 300 36 331
rect 4210 381 4302 397
rect 4210 347 4252 381
rect 4286 347 4302 381
rect 4210 331 4302 347
rect 4210 326 4240 331
rect -56 -51 36 -35
rect -56 -85 -40 -51
rect -6 -85 36 -51
rect -56 -101 36 -85
rect 6 -106 36 -101
rect 4210 -51 4302 -35
rect 4210 -85 4252 -51
rect 4286 -85 4302 -51
rect 4210 -101 4302 -85
rect 4210 -132 4240 -101
rect 6 -833 36 -821
rect -56 -849 36 -833
rect -56 -883 -40 -849
rect -6 -883 36 -849
rect -56 -898 36 -883
rect 4210 -833 4240 -802
rect 4210 -849 4302 -833
rect 4210 -883 4252 -849
rect 4286 -883 4302 -849
rect -56 -899 10 -898
rect 4210 -899 4302 -883
rect 6 -1265 36 -1234
rect -56 -1281 36 -1265
rect -56 -1315 -40 -1281
rect -6 -1315 36 -1281
rect -56 -1331 36 -1315
rect 4210 -1265 4240 -1234
rect 4210 -1281 4302 -1265
rect 4210 -1315 4252 -1281
rect 4286 -1315 4302 -1281
rect 4210 -1331 4302 -1315
<< polycont >>
rect -40 347 -6 381
rect 4252 347 4286 381
rect -40 -85 -6 -51
rect 4252 -85 4286 -51
rect -40 -883 -6 -849
rect 4252 -883 4286 -849
rect -40 -1315 -6 -1281
rect 4252 -1315 4286 -1281
<< locali >>
rect -40 381 -6 397
rect -40 300 -6 347
rect 4252 381 4286 397
rect 4252 298 4286 347
rect -40 -51 -6 -35
rect -40 -137 -6 -85
rect 4252 -51 4286 -35
rect 4252 -132 4286 -85
rect -40 -849 -6 -792
rect -40 -899 -6 -883
rect 4252 -849 4286 -802
rect 4252 -899 4286 -883
rect -40 -1281 -6 -1234
rect -40 -1331 -6 -1315
rect 4252 -1281 4286 -1234
rect 4252 -1331 4286 -1315
<< viali >>
rect -214 446 -129 480
rect -129 446 4375 480
rect 4375 446 4460 480
rect -214 420 -180 446
rect -214 -1354 -180 420
rect 4426 420 4460 446
rect -40 347 -6 381
rect 4252 347 4286 381
rect -40 -85 -6 -51
rect 4252 -85 4286 -51
rect -40 -883 -6 -849
rect 4252 -883 4286 -849
rect -40 -1315 -6 -1281
rect 4252 -1315 4286 -1281
rect -214 -1380 -180 -1354
rect 4426 -1354 4460 420
rect 4426 -1380 4460 -1354
rect -214 -1414 -129 -1380
rect -129 -1414 4375 -1380
rect 4375 -1414 4460 -1380
<< metal1 >>
rect -220 486 -174 492
rect 2100 486 2146 492
rect 4420 486 4466 492
rect -226 480 4472 486
rect -226 440 -214 480
rect -220 -1374 -214 440
rect -226 -1414 -214 -1374
rect -180 440 4426 446
rect -180 -1374 -174 440
rect -46 381 0 393
rect -46 347 -40 381
rect -6 347 0 381
rect -46 300 0 347
rect 2100 288 2146 440
rect 4246 381 4292 393
rect 4246 347 4252 381
rect 4286 347 4292 381
rect 4246 300 4292 347
rect 4194 295 4292 300
rect 4194 288 4272 295
rect -46 59 0 116
rect 2087 112 2097 288
rect 2149 112 2159 288
rect 4145 112 4155 288
rect 4207 112 4272 288
rect 42 59 88 108
rect 4194 100 4272 112
rect -133 13 4379 59
rect -133 -346 -87 13
rect -46 -51 0 -39
rect -46 -85 -40 -51
rect -6 -85 0 -51
rect -46 -132 0 -85
rect 4246 -51 4292 -39
rect 4246 -85 4252 -51
rect 4286 -85 4292 -51
rect 4246 -132 4292 -85
rect -46 -144 61 -132
rect -46 -145 39 -144
rect -21 -320 39 -145
rect 91 -320 101 -144
rect 2087 -320 2097 -144
rect 2149 -320 2159 -144
rect -21 -332 61 -320
rect 4175 -322 4274 -132
rect 4158 -332 4274 -322
rect -142 -352 -78 -346
rect -142 -404 -136 -352
rect -84 -404 -78 -352
rect -142 -410 -78 -404
rect 590 -444 1598 -411
rect 2648 -444 3656 -412
rect 4158 -444 4204 -332
rect 4333 -346 4379 13
rect 4324 -352 4388 -346
rect 4324 -404 4330 -352
rect 4382 -404 4388 -352
rect 4324 -410 4388 -404
rect 42 -490 4204 -444
rect -142 -530 -78 -524
rect -142 -582 -136 -530
rect -84 -582 -78 -530
rect -142 -588 -78 -582
rect -133 -947 -87 -588
rect 42 -602 88 -490
rect 590 -518 1598 -490
rect 2648 -519 3656 -490
rect 4324 -530 4388 -524
rect 4324 -582 4330 -530
rect 4382 -582 4388 -530
rect 4324 -588 4388 -582
rect -44 -611 88 -602
rect -44 -791 62 -611
rect 4180 -614 4279 -602
rect 2087 -790 2097 -614
rect 2149 -790 2159 -614
rect 4145 -790 4155 -614
rect 4207 -790 4279 -614
rect -46 -802 62 -791
rect 4180 -802 4279 -790
rect -46 -849 0 -802
rect -46 -883 -40 -849
rect -6 -883 0 -849
rect -46 -895 0 -883
rect 4246 -849 4292 -802
rect 4246 -883 4252 -849
rect 4286 -883 4292 -849
rect 4246 -895 4292 -883
rect 4333 -947 4379 -588
rect -133 -993 740 -947
rect 1575 -993 2671 -947
rect 3624 -993 4379 -947
rect -19 -1046 59 -1034
rect 4158 -1041 4204 -993
rect -19 -1222 39 -1046
rect 91 -1222 101 -1046
rect 2087 -1222 2097 -1046
rect 2149 -1222 2159 -1046
rect 4246 -1047 4292 -993
rect -19 -1234 59 -1222
rect -46 -1281 0 -1234
rect -46 -1315 -40 -1281
rect -6 -1315 0 -1281
rect -46 -1327 0 -1315
rect 2100 -1374 2146 -1222
rect 4246 -1281 4292 -1234
rect 4246 -1315 4252 -1281
rect 4286 -1315 4292 -1281
rect 4246 -1327 4292 -1315
rect 4420 -1374 4426 440
rect -180 -1380 4426 -1374
rect 4460 440 4472 480
rect 4460 -1374 4466 440
rect 4460 -1414 4472 -1374
rect -226 -1420 4472 -1414
rect -220 -1426 -174 -1420
rect 2100 -1426 2146 -1420
rect 4420 -1426 4466 -1420
<< via1 >>
rect 2097 112 2149 288
rect 4155 112 4207 288
rect 39 -320 91 -144
rect 2097 -320 2149 -144
rect -136 -404 -84 -352
rect 4330 -404 4382 -352
rect -136 -582 -84 -530
rect 4330 -582 4382 -530
rect 2097 -790 2149 -614
rect 4155 -790 4207 -614
rect 39 -1222 91 -1046
rect 2097 -1222 2149 -1046
<< metal2 >>
rect 2097 288 2149 298
rect 2095 112 2097 152
rect 2095 -134 2149 112
rect 4153 288 4209 298
rect 4153 102 4209 112
rect 39 -144 91 -134
rect -142 -352 -78 -346
rect -142 -404 -136 -352
rect -84 -404 -78 -352
rect -142 -410 -78 -404
rect -133 -524 -87 -410
rect 39 -441 91 -320
rect 2095 -144 2151 -134
rect 2095 -330 2151 -320
rect 4324 -352 4388 -346
rect 4324 -404 4330 -352
rect 4382 -404 4388 -352
rect 4324 -410 4388 -404
rect 39 -493 4207 -441
rect -142 -530 -78 -524
rect -142 -582 -136 -530
rect -84 -582 -78 -530
rect -142 -588 -78 -582
rect 2095 -614 2151 -604
rect 2095 -800 2151 -790
rect 4155 -614 4207 -493
rect 4333 -524 4379 -410
rect 4324 -530 4388 -524
rect 4324 -582 4330 -530
rect 4382 -582 4388 -530
rect 4324 -588 4388 -582
rect 4155 -800 4207 -790
rect 37 -1046 93 -1036
rect 37 -1232 93 -1222
rect 2097 -1046 2151 -800
rect 2149 -1064 2151 -1046
rect 2097 -1232 2149 -1222
<< via2 >>
rect 4153 112 4155 288
rect 4155 112 4207 288
rect 4207 112 4209 288
rect 2095 -320 2097 -144
rect 2097 -320 2149 -144
rect 2149 -320 2151 -144
rect 2095 -790 2097 -614
rect 2097 -790 2149 -614
rect 2149 -790 2151 -614
rect 37 -1222 39 -1046
rect 39 -1222 91 -1046
rect 91 -1222 93 -1046
<< metal3 >>
rect 4143 288 4219 293
rect 4143 112 4153 288
rect 4209 112 4219 288
rect 4143 107 4219 112
rect 4151 26 4211 107
rect 4151 -34 4386 26
rect 2085 -144 2161 -139
rect 2081 -320 2091 -144
rect 2155 -320 2165 -144
rect 2085 -325 2161 -320
rect 4326 -437 4386 -34
rect -140 -497 4386 -437
rect -140 -900 -80 -497
rect 2085 -614 2161 -609
rect 2081 -790 2091 -614
rect 2155 -790 2165 -614
rect 2085 -795 2161 -790
rect -140 -960 95 -900
rect 35 -1041 95 -960
rect 27 -1046 103 -1041
rect 27 -1222 37 -1046
rect 93 -1222 103 -1046
rect 27 -1227 103 -1222
<< via3 >>
rect 2091 -320 2095 -144
rect 2095 -320 2151 -144
rect 2151 -320 2155 -144
rect 2091 -790 2095 -614
rect 2095 -790 2151 -614
rect 2151 -790 2155 -614
<< metal4 >>
rect 2090 -144 2156 -143
rect 2090 -320 2091 -144
rect 2155 -320 2156 -144
rect 2090 -321 2156 -320
rect 2091 -613 2155 -321
rect 2090 -614 2156 -613
rect 2090 -790 2091 -614
rect 2155 -790 2156 -614
rect 2090 -791 2156 -790
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_0
timestamp 1717765832
transform 1 0 21 0 1 -702
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_1
timestamp 1717765832
transform 1 0 4225 0 1 -1134
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_2
timestamp 1717765832
transform 1 0 4225 0 1 -702
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_3
timestamp 1717765832
transform 1 0 4225 0 1 -232
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_4
timestamp 1717765832
transform 1 0 4225 0 1 200
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_5
timestamp 1717765832
transform 1 0 21 0 1 200
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_6
timestamp 1717765832
transform 1 0 21 0 1 -232
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_7
timestamp 1717765832
transform 1 0 21 0 1 -1134
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_8RMJP2  sky130_fd_pr__pfet_01v8_8RMJP2_0
timestamp 1717765832
transform 1 0 2123 0 1 -1098
box -2123 -198 2123 164
use sky130_fd_pr__pfet_01v8_8RMJP2  sky130_fd_pr__pfet_01v8_8RMJP2_1
timestamp 1717765832
transform 1 0 2123 0 1 -666
box -2123 -198 2123 164
use sky130_fd_pr__pfet_01v8_CVRJBD  sky130_fd_pr__pfet_01v8_CVRJBD_0
timestamp 1717765832
transform 1 0 2123 0 1 -268
box -2123 -164 2123 198
use sky130_fd_pr__pfet_01v8_CVRJBD  sky130_fd_pr__pfet_01v8_CVRJBD_1
timestamp 1717765832
transform 1 0 2123 0 1 164
box -2123 -164 2123 198
<< labels >>
flabel metal1 2119 423 2119 423 1 FreeSans 160 0 0 0 vdde
port 0 n
flabel metal3 4176 73 4176 73 1 FreeSans 160 0 0 0 D3
port 1 n
flabel metal1 4190 -425 4190 -425 1 FreeSans 160 0 0 0 D9
port 4 n
flabel metal2 4182 -560 4182 -560 1 FreeSans 160 0 0 0 D8
port 5 n
flabel metal1 -209 -1418 -209 -1418 0 FreeSans 1600 0 0 0 VDDE
port 7 nsew
flabel metal1 4058 25 4058 25 1 FreeSans 160 0 0 0 D4
port 3 n
<< end >>
