magic
tech sky130A
magscale 1 2
timestamp 1718866891
<< xpolycontact >>
rect -450 1052 -380 1484
rect -450 52 -380 484
rect -284 1052 -214 1484
rect -284 52 -214 484
rect -118 1052 -48 1484
rect -118 52 -48 484
rect 48 1052 118 1484
rect 48 52 118 484
rect 214 1052 284 1484
rect 214 52 284 484
rect 380 1052 450 1484
rect 380 52 450 484
rect -450 -484 -380 -52
rect -450 -1484 -380 -1052
rect -284 -484 -214 -52
rect -284 -1484 -214 -1052
rect -118 -484 -48 -52
rect -118 -1484 -48 -1052
rect 48 -484 118 -52
rect 48 -1484 118 -1052
rect 214 -484 284 -52
rect 214 -1484 284 -1052
rect 380 -484 450 -52
rect 380 -1484 450 -1052
<< ppolyres >>
rect -450 484 -380 1052
rect -284 484 -214 1052
rect -118 484 -48 1052
rect 48 484 118 1052
rect 214 484 284 1052
rect 380 484 450 1052
rect -450 -1052 -380 -484
rect -284 -1052 -214 -484
rect -118 -1052 -48 -484
rect 48 -1052 118 -484
rect 214 -1052 284 -484
rect 380 -1052 450 -484
<< viali >>
rect -434 1069 -396 1466
rect -268 1069 -230 1466
rect -102 1069 -64 1466
rect 64 1069 102 1466
rect 230 1069 268 1466
rect 396 1069 434 1466
rect -434 70 -396 467
rect -268 70 -230 467
rect -102 70 -64 467
rect 64 70 102 467
rect 230 70 268 467
rect 396 70 434 467
rect -434 -467 -396 -70
rect -268 -467 -230 -70
rect -102 -467 -64 -70
rect 64 -467 102 -70
rect 230 -467 268 -70
rect 396 -467 434 -70
rect -434 -1466 -396 -1069
rect -268 -1466 -230 -1069
rect -102 -1466 -64 -1069
rect 64 -1466 102 -1069
rect 230 -1466 268 -1069
rect 396 -1466 434 -1069
<< metal1 >>
rect -440 1466 -390 1478
rect -440 1069 -434 1466
rect -396 1069 -390 1466
rect -440 1057 -390 1069
rect -274 1466 -224 1478
rect -274 1069 -268 1466
rect -230 1069 -224 1466
rect -274 1057 -224 1069
rect -108 1466 -58 1478
rect -108 1069 -102 1466
rect -64 1069 -58 1466
rect -108 1057 -58 1069
rect 58 1466 108 1478
rect 58 1069 64 1466
rect 102 1069 108 1466
rect 58 1057 108 1069
rect 224 1466 274 1478
rect 224 1069 230 1466
rect 268 1069 274 1466
rect 224 1057 274 1069
rect 390 1466 440 1478
rect 390 1069 396 1466
rect 434 1069 440 1466
rect 390 1057 440 1069
rect -440 467 -390 479
rect -440 70 -434 467
rect -396 70 -390 467
rect -440 58 -390 70
rect -274 467 -224 479
rect -274 70 -268 467
rect -230 70 -224 467
rect -274 58 -224 70
rect -108 467 -58 479
rect -108 70 -102 467
rect -64 70 -58 467
rect -108 58 -58 70
rect 58 467 108 479
rect 58 70 64 467
rect 102 70 108 467
rect 58 58 108 70
rect 224 467 274 479
rect 224 70 230 467
rect 268 70 274 467
rect 224 58 274 70
rect 390 467 440 479
rect 390 70 396 467
rect 434 70 440 467
rect 390 58 440 70
rect -440 -70 -390 -58
rect -440 -467 -434 -70
rect -396 -467 -390 -70
rect -440 -479 -390 -467
rect -274 -70 -224 -58
rect -274 -467 -268 -70
rect -230 -467 -224 -70
rect -274 -479 -224 -467
rect -108 -70 -58 -58
rect -108 -467 -102 -70
rect -64 -467 -58 -70
rect -108 -479 -58 -467
rect 58 -70 108 -58
rect 58 -467 64 -70
rect 102 -467 108 -70
rect 58 -479 108 -467
rect 224 -70 274 -58
rect 224 -467 230 -70
rect 268 -467 274 -70
rect 224 -479 274 -467
rect 390 -70 440 -58
rect 390 -467 396 -70
rect 434 -467 440 -70
rect 390 -479 440 -467
rect -440 -1069 -390 -1057
rect -440 -1466 -434 -1069
rect -396 -1466 -390 -1069
rect -440 -1478 -390 -1466
rect -274 -1069 -224 -1057
rect -274 -1466 -268 -1069
rect -230 -1466 -224 -1069
rect -274 -1478 -224 -1466
rect -108 -1069 -58 -1057
rect -108 -1466 -102 -1069
rect -64 -1466 -58 -1069
rect -108 -1478 -58 -1466
rect 58 -1069 108 -1057
rect 58 -1466 64 -1069
rect 102 -1466 108 -1069
rect 58 -1478 108 -1466
rect 224 -1069 274 -1057
rect 224 -1466 230 -1069
rect 268 -1466 274 -1069
rect 224 -1478 274 -1466
rect 390 -1069 440 -1057
rect 390 -1466 396 -1069
rect 434 -1466 440 -1069
rect 390 -1478 440 -1466
<< properties >>
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.350 l 3 m 2 nx 6 wmin 0.350 lmin 0.50 rho 319.8 val 3.854k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
